/*E5M2
inf:        S.11111.00
NaN:        S.11111.{01, 10, 11}
zero:       S.00000.00
normal_max: S.11110.11 = ±57,344
normal_min: S.00001.00 = ±2^(-14)
subnor_max: S.00000.11 = ±0.75 * 2^(-14)
subnor_min: S.00000.01 = ±2^(-16)
exp_bias:   15
*/

//scalar mul, should be vector tho
module e5m2_MULT #(
    //parameters
) (
    /* implement these later
    input  logic                 clk_i,
    input  logic                 rst_ni,
    output logic                 a_ready_o,
    input  logic                 a_valid_o,
    output logic                 b_ready_o,
    input  logic                 b_valid_o,
    output logic                 b_ready_o,
    input  logic                 b_valid_o,
    input  logic                 mode_i,                  
    */
    input  logic [7:0]           a_i,
    input  logic [7:0]           b_i,
    output logic [7:0]           c_o,
    output logic                 inf,
    output logic                 NaN 
    //store intermediate in E6M4
    //output of MAC should be fp16 or fp32, TODO: verify this, should we convert it back in FP8 again?

);

    //////////////////////////////////parameters//////////////////////////////////////////////
    localparam int MANT_BITS  = 2;
    localparam int EXP_BITS   = 5;
    localparam int EXP_MAX    = (1<<EXP_BITS)-1;   // 31
    localparam int EXP_BIAS   = 15;                // e5 bias
    localparam int SIG_NORM_HI_BIT = MANT_BITS;    // for e5m2, 2 (so '1xx' => [4..7])
 
    //////////////////////////////////variables////////////////////////////////////////////////       
    logic a_sign;                 logic b_sign;              logic c_sign;
    logic [EXP_BITS-1:0]  a_exp;  logic [EXP_BITS-1:0]    b_exp;
    logic [MANT_BITS-1:0] a_man;  logic [MANT_BITS-1:0]   b_man;
    logic [EXP_BITS*2-1:0]    c_exp;  logic [MANT_BITS*2+1:0] c_man;
    //////////////////////////////////Functions////////////////////////////////////////////////
    //get sign, mentissa, exp
    function automatic void unpack(
    input  logic [7:0] in,
    output logic       sign,
    output logic [EXP_BITS-1:0] exp,
    output logic [MANT_BITS-1:0] mant
    );
    sign = in[7];
    exp  = in[6:2];
    mant = in[1:0];
    endfunction
    
    //////////////////////////////////Main logic////////////////////////////////////////////////
    
    /*E5M2
    inf:        S.11111.00
    NaN:        S.11111.{01, 10, 11}
    zero:       S.00000.00
    normal_max: S.11110.11 = ±57,344
    normal_min: S.00001.00 = ±2^(-14)
    subnor_max: S.00000.11 = ±0.75 * 2^(-14)
    subnor_min: S.00000.01 = ±2^(-16)
    exp_bias:   15
    */

    //exponent add
    always_comb begin
        unpack(a_i, a_sign, a_exp, a_man);
        unpack(b_i, b_sign, b_exp, b_man);
        if((a_exp==EXP_MAX&&a_man!=0)||(b_exp==EXP_MAX&&b_man!=0))begin
            //NaN prod anything is NaN
            c_exp = 6'b011111;
            c_man = 4'b0100;
            c_sign = 0;
            NaN = 1;
            inf = 0;
        end else if((a_exp==EXP_MAX&&a_man==0)||(b_exp==EXP_MAX&&b_man==0)) begin
            //when one of them is inf
            if((a_exp==0&&a_man==0)||(b_exp==0&&b_man==0))begin
                //when one inf one zero, set as NaN
                c_exp = 6'b011111;
                c_man = 4'b0100;
                c_sign = 0;
                NaN = 1;
                inf = 0;
            end else begin
                //otherwise also inf
                c_exp = 6'b011111;
                c_man = 0;
                c_sign = 0;
                NaN = 0;
                inf = 1;
            end
        end else if ((a_exp==0&&a_man==0)||(b_exp==0&&b_man==0)) begin
            //zero
            if((a_exp==EXP_MAX&&a_man==0)||(b_exp==EXP_MAX&&b_man==0))begin
                //when one inf one zero, set as NaN
                c_exp = 6'b011111;
                c_man = 4'b0100;
                c_sign = 0;
                NaN = 1;
                inf = 0;
            end else begin
                c_exp = 0;
                c_man = 0;
                c_sign = 0;
                NaN = 0;
                inf = 0;
            end    
        end else begin
            c_sign = a_sign^b_sign;
            NaN = 0;
            inf = c_exp[EXP_BITS];
            if (a_exp==0&&b_exp==0) begin   
                //subnormal*subnormal
                c_exp = a_exp + b_exp-EXP_BIAS+2;
                c_man = {1'b0,a_man}*{1'b0,b_man};
            end else if (a_exp==0&&b_exp!=0) begin
                //subnormal*normal
                c_exp = a_exp + b_exp-EXP_BIAS+1;
                c_man = {1'b0,a_man}*{1'b1,b_man};
            end else if (a_exp!=0&&b_exp==0) begin
                //normal*subnormal
                c_exp = a_exp + b_exp-EXP_BIAS+1;
                c_man = {1'b1,a_man}*{1'b0,b_man};
            end else begin
                //normal*normal
                c_exp = a_exp + b_exp-EXP_BIAS;
                if (inf) begin
                    //TODO: overflow case
                    c_exp = 6'b011111;
                    c_man = 0;
                end else begin
                    c_man = {1'b1,a_man}*{1'b1,b_man};
                    if(c_man[EXP_BITS*2-1]==1)begin
                        c_exp = c_exp+1;
                        c_man = c_man>>1;
                    end
                end
            end
            
        end   
    end
    assign c_o = {c_sign,c_exp[EXP_BITS-1:0],c_man[MANT_BITS*2-1 -:MANT_BITS-1]};
    

    

    //normally, Xa+Xb, Pa+Pb
    //remember when doing mult,加上尾数隐含的一位，比如mantissa：10， 实际大小为1.10
    //case like 1.10* 1.10 = 10.0100, need to put the extra 1 in the exponent
    //
    

endmodule


/*detect special cases
    function automatic bit is_nan   (input logic [EXP_BITS-1:0] e, input logic [MANT_BITS-1:0] m);
    return (e == EXP_MAX) && (m != 0);
    endfunction
    function automatic bit is_inf   (input logic [EXP_BITS-1:0] e, input logic [MANT_BITS-1:0] m);
    return (e == EXP_MAX) && (m == 0);
    endfunction
    function automatic bit is_zero  (input logic [EXP_BITS-1:0] e, input logic [MANT_BITS-1:0] m);
    return (e == 0) && (m == 0);
    endfunction
    function automatic bit is_sub   (input logic [EXP_BITS-1:0] e, input logic [MANT_BITS-1:0] m);
    return (e == 0) && (m != 0);
    endfunction
    function automatic bit is_norm  (input logic [EXP_BITS-1:0] e);
    return (e != 0) && (e != EXP_MAX);
    endfunction*/