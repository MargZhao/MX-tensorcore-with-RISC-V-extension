module tb_pt_MAC_long_better;

timeunit 1ns;
timeprecision 1ps;

logic clk_i;
logic rstn;

always begin #{CLK_HALF}ns; clk_i <= ~clk_i; end

localparam M_out_width = {M_OUT_WIDTH};

logic [7:0] a_mant0,a_mant1,a_mant2,a_mant3;
logic [7:0] b_mant0,b_mant1,b_mant2,b_mant3;
logic [9:0] a_exp0,a_exp1,a_exp2,a_exp3;
logic [9:0] b_exp0,b_exp1,b_exp2,b_exp3;
logic [3:0] a_sign0,a_sign1,a_sign2,a_sign3;
logic [3:0] b_sign0,b_sign1,b_sign2,b_sign3;
logic [1:0] prec_mode;
logic [1:0] FP_mode;/*
logic [22:0] out_mant;
logic [7:0]  out_exp;
logic        out_sign;*/
logic [M_out_width-1:0] MAC_mant_out;
logic [7:0]  MAC_exp_out;
logic        MAC_sign_out;
logic [7:0] shared_exps0;
logic [7:0] shared_exps1;


//DUT
/*
  MX_MAC_EA MX_MAC0 (.clk_i(clk_i), .rstn(rstn), .a_mant0(a_mant0), .a_mant1(a_mant1), .a_mant2(a_mant2), .a_mant3(a_mant3), 
  .b_mant0(b_mant0), .b_mant1(b_mant1), .b_mant2(b_mant2), .b_mant3(b_mant3), .a_exp_in0(a_exp0), .a_exp_in1(a_exp1), .a_exp_in2(a_exp2), .a_exp_in3(a_exp3),
  .b_exp_in0(b_exp0), .b_exp_in1(b_exp1), .b_exp_in2(b_exp2), .b_exp_in3(b_exp3), .a_sign_in0(a_sign0), .a_sign_in1(a_sign1), .a_sign_in2(a_sign2), .a_sign_in3(a_sign3),
  .b_sign_in0(b_sign0), .b_sign_in1(b_sign1), .b_sign_in2(b_sign2), .b_sign_in3(b_sign3), .prec_mode(prec_mode), .FP_mode(FP_mode), .MAC_mant_out(MAC_mant_out), .MAC_exp_out(MAC_exp_out), .MAC_sign_out(MAC_sign_out),
  .shared_exps0(shared_exps0), .shared_exps1(shared_exps1));
*/

  MX_MAC MX_MAC0 (.clk_i(clk_i), .rstn(rstn), .a_mant0(a_mant0), .a_mant1(a_mant1), .a_mant2(a_mant2), .a_mant3(a_mant3), 
  .b_mant0(b_mant0), .b_mant1(b_mant1), .b_mant2(b_mant2), .b_mant3(b_mant3), .a_exp_in0(a_exp0), .a_exp_in1(a_exp1), .a_exp_in2(a_exp2), .a_exp_in3(a_exp3),
  .b_exp_in0(b_exp0), .b_exp_in1(b_exp1), .b_exp_in2(b_exp2), .b_exp_in3(b_exp3), .a_sign_in0(a_sign0), .a_sign_in1(a_sign1), .a_sign_in2(a_sign2), .a_sign_in3(a_sign3),
  .b_sign_in0(b_sign0), .b_sign_in1(b_sign1), .b_sign_in2(b_sign2), .b_sign_in3(b_sign3), .prec_mode(prec_mode), .FP_mode(FP_mode), .MAC_mant_out(MAC_mant_out), .MAC_exp_out(MAC_exp_out), .MAC_sign_out(MAC_sign_out),
  .shared_exps0(shared_exps0), .shared_exps1(shared_exps1));


/*
ST_mul ST_mul0 (.a_mant0(a_mant0), .a_mant1(a_mant1), .a_mant2(a_mant2), .a_mant3(a_mant3), .b_mant0(b_mant0), .b_mant1(b_mant1), .b_mant2(b_mant2), .b_mant3(b_mant3), 
.a_exp_in0(a_exp0), .a_exp_in1(a_exp1), .a_exp_in2(a_exp2), .a_exp_in3(a_exp3), .b_exp_in0(b_exp0), .b_exp_in1(b_exp1), .b_exp_in2(b_exp2), .b_exp_in3(b_exp3), .a_sign_in0(a_sign0), .a_sign_in1(a_sign1), .a_sign_in2(a_sign2), .a_sign_in3(a_sign3), 
.b_sign_in0(b_sign0), .b_sign_in1(b_sign1), .b_sign_in2(b_sign2), .b_sign_in3(b_sign3), .prec_mode(prec_mode), .FP_mode(FP_mode), .out_mant(out_mant), .out_exp(out_exp), .out_sign(out_sign));
*/

// SDF annotation
initial begin
	$sdf_annotate("/{OUTER_FOLDER}/Ours_old/syn/outputs/{DIR_LOC_TEMP}/MX_MAC_mapped.sdf", MX_MAC0);
end

initial begin
prec_mode = {PREC_MODE};
FP_mode = {FP_MODE};
shared_exps0 = 'd127;
shared_exps1 = 'd127;

clk_i = 0;
rstn = 0;

a_mant0 = 8'd95; a_mant1 = 8'd95; a_mant2 = 8'd95; a_mant3 = '0;
b_mant0 = 8'd112; b_mant1 = 8'd112; b_mant2 = 8'd112; b_mant3 = 8'd112;
a_exp0 = 10'd6; a_exp1 = 10'd6; a_exp2 = 10'd6; a_exp3 = 10'd6;
b_exp0 = 10'd520; b_exp1 = 10'd520; b_exp2 = 10'd520; b_exp3 = 10'd520;
a_sign0 = 4'd0; a_sign1 = 4'd0; a_sign2 = 4'd0; a_sign3 = 4'd0;
b_sign0 = 4'd0; b_sign1 = 4'd0; b_sign2 = 4'd0; b_sign3 = 4'd0;


@(posedge clk_i);
#0.1ns;
rstn = 1;

$dumpfile("/{OUTER_FOLDER}/Ours_old/sim-syn/vcd/{DIR_LOC_TEMP}/MX_MAC_{WORKLOAD}.vcd");
$dumpvars(0, tb_pt_MAC_long_better);
$dumpon;

@(posedge clk_i);
shared_exps0 = 8'd152;
shared_exps1 = 8'd135;
rstn = 0;
@(posedge clk_i);
rstn = 1;
a_mant0 = 8'd188; a_mant1 = 8'd228; a_mant2 = 8'd73; a_mant3 = 8'd244;
b_mant0 = 8'd25; b_mant1 = 8'd161; b_mant2 = 8'd100; b_mant3 = 8'd218;
a_exp0 = 10'd638; a_exp1 = 10'd381; a_exp2 = 10'd682; a_exp3 = 10'd750;
b_exp0 = 10'd760; b_exp1 = 10'd732; b_exp2 = 10'd42; b_exp3 = 10'd355;
a_sign0 = 4'd5; a_sign1 = 4'd10; a_sign2 = 4'd10; a_sign3 = 4'd6;
b_sign0 = 4'd14; b_sign1 = 4'd11; b_sign2 = 4'd15; b_sign3 = 4'd16;
@(posedge clk_i);
a_mant0 = 8'd30; a_mant1 = 8'd9; a_mant2 = 8'd201; a_mant3 = 8'd133;
b_mant0 = 8'd35; b_mant1 = 8'd75; b_mant2 = 8'd185; b_mant3 = 8'd91;
a_exp0 = 10'd905; a_exp1 = 10'd589; a_exp2 = 10'd29; a_exp3 = 10'd474;
b_exp0 = 10'd794; b_exp1 = 10'd87; b_exp2 = 10'd550; b_exp3 = 10'd573;
a_sign0 = 4'd8; a_sign1 = 4'd12; a_sign2 = 4'd9; a_sign3 = 4'd12;
b_sign0 = 4'd10; b_sign1 = 4'd6; b_sign2 = 4'd1; b_sign3 = 4'd6;
@(posedge clk_i);
a_mant0 = 8'd177; a_mant1 = 8'd35; a_mant2 = 8'd44; a_mant3 = 8'd211;
b_mant0 = 8'd92; b_mant1 = 8'd65; b_mant2 = 8'd86; b_mant3 = 8'd252;
a_exp0 = 10'd186; a_exp1 = 10'd68; a_exp2 = 10'd403; a_exp3 = 10'd4;
b_exp0 = 10'd260; b_exp1 = 10'd551; b_exp2 = 10'd986; b_exp3 = 10'd53;
a_sign0 = 4'd14; a_sign1 = 4'd12; a_sign2 = 4'd10; a_sign3 = 4'd4;
b_sign0 = 4'd7; b_sign1 = 4'd2; b_sign2 = 4'd1; b_sign3 = 4'd1;
@(posedge clk_i);
a_mant0 = 8'd7; a_mant1 = 8'd109; a_mant2 = 8'd163; a_mant3 = 8'd64;
b_mant0 = 8'd39; b_mant1 = 8'd87; b_mant2 = 8'd212; b_mant3 = 8'd155;
a_exp0 = 10'd746; a_exp1 = 10'd79; a_exp2 = 10'd611; a_exp3 = 10'd130;
b_exp0 = 10'd541; b_exp1 = 10'd190; b_exp2 = 10'd705; b_exp3 = 10'd190;
a_sign0 = 4'd11; a_sign1 = 4'd4; a_sign2 = 4'd13; a_sign3 = 4'd2;
b_sign0 = 4'd2; b_sign1 = 4'd6; b_sign2 = 4'd7; b_sign3 = 4'd0;
@(posedge clk_i);
a_mant0 = 8'd140; a_mant1 = 8'd21; a_mant2 = 8'd163; a_mant3 = 8'd192;
b_mant0 = 8'd250; b_mant1 = 8'd63; b_mant2 = 8'd30; b_mant3 = 8'd225;
a_exp0 = 10'd270; a_exp1 = 10'd917; a_exp2 = 10'd74; a_exp3 = 10'd694;
b_exp0 = 10'd245; b_exp1 = 10'd581; b_exp2 = 10'd216; b_exp3 = 10'd374;
a_sign0 = 4'd6; a_sign1 = 4'd12; a_sign2 = 4'd2; a_sign3 = 4'd2;
b_sign0 = 4'd4; b_sign1 = 4'd15; b_sign2 = 4'd3; b_sign3 = 4'd15;
@(posedge clk_i);
a_mant0 = 8'd16; a_mant1 = 8'd112; a_mant2 = 8'd119; a_mant3 = 8'd128;
b_mant0 = 8'd209; b_mant1 = 8'd73; b_mant2 = 8'd7; b_mant3 = 8'd111;
a_exp0 = 10'd371; a_exp1 = 10'd1019; a_exp2 = 10'd175; a_exp3 = 10'd471;
b_exp0 = 10'd554; b_exp1 = 10'd269; b_exp2 = 10'd252; b_exp3 = 10'd105;
a_sign0 = 4'd15; a_sign1 = 4'd10; a_sign2 = 4'd16; a_sign3 = 4'd7;
b_sign0 = 4'd16; b_sign1 = 4'd3; b_sign2 = 4'd16; b_sign3 = 4'd7;
@(posedge clk_i);
a_mant0 = 8'd76; a_mant1 = 8'd98; a_mant2 = 8'd96; a_mant3 = 8'd155;
b_mant0 = 8'd120; b_mant1 = 8'd95; b_mant2 = 8'd133; b_mant3 = 8'd111;
a_exp0 = 10'd485; a_exp1 = 10'd93; a_exp2 = 10'd975; a_exp3 = 10'd210;
b_exp0 = 10'd573; b_exp1 = 10'd494; b_exp2 = 10'd814; b_exp3 = 10'd722;
a_sign0 = 4'd5; a_sign1 = 4'd0; a_sign2 = 4'd13; a_sign3 = 4'd12;
b_sign0 = 4'd11; b_sign1 = 4'd8; b_sign2 = 4'd16; b_sign3 = 4'd0;
@(posedge clk_i);
shared_exps0 = 8'd130;
shared_exps1 = 8'd111;
a_mant0 = 8'd19; a_mant1 = 8'd228; a_mant2 = 8'd116; a_mant3 = 8'd171;
b_mant0 = 8'd51; b_mant1 = 8'd5; b_mant2 = 8'd128; b_mant3 = 8'd101;
a_exp0 = 10'd545; a_exp1 = 10'd550; a_exp2 = 10'd863; a_exp3 = 10'd302;
b_exp0 = 10'd818; b_exp1 = 10'd986; b_exp2 = 10'd999; b_exp3 = 10'd968;
a_sign0 = 4'd6; a_sign1 = 4'd11; a_sign2 = 4'd6; a_sign3 = 4'd1;
b_sign0 = 4'd6; b_sign1 = 4'd16; b_sign2 = 4'd14; b_sign3 = 4'd5;
@(posedge clk_i);
a_mant0 = 8'd192; a_mant1 = 8'd49; a_mant2 = 8'd231; a_mant3 = 8'd34;
b_mant0 = 8'd0; b_mant1 = 8'd215; b_mant2 = 8'd138; b_mant3 = 8'd129;
a_exp0 = 10'd991; a_exp1 = 10'd131; a_exp2 = 10'd876; a_exp3 = 10'd759;
b_exp0 = 10'd557; b_exp1 = 10'd293; b_exp2 = 10'd642; b_exp3 = 10'd241;
a_sign0 = 4'd4; a_sign1 = 4'd13; a_sign2 = 4'd5; a_sign3 = 4'd13;
b_sign0 = 4'd10; b_sign1 = 4'd4; b_sign2 = 4'd13; b_sign3 = 4'd4;
@(posedge clk_i);
a_mant0 = 8'd109; a_mant1 = 8'd63; a_mant2 = 8'd145; a_mant3 = 8'd116;
b_mant0 = 8'd187; b_mant1 = 8'd32; b_mant2 = 8'd230; b_mant3 = 8'd139;
a_exp0 = 10'd284; a_exp1 = 10'd440; a_exp2 = 10'd235; a_exp3 = 10'd683;
b_exp0 = 10'd82; b_exp1 = 10'd725; b_exp2 = 10'd232; b_exp3 = 10'd558;
a_sign0 = 4'd0; a_sign1 = 4'd5; a_sign2 = 4'd14; a_sign3 = 4'd2;
b_sign0 = 4'd16; b_sign1 = 4'd0; b_sign2 = 4'd14; b_sign3 = 4'd15;
@(posedge clk_i);
a_mant0 = 8'd13; a_mant1 = 8'd89; a_mant2 = 8'd231; a_mant3 = 8'd27;
b_mant0 = 8'd216; b_mant1 = 8'd79; b_mant2 = 8'd1; b_mant3 = 8'd50;
a_exp0 = 10'd513; a_exp1 = 10'd523; a_exp2 = 10'd640; a_exp3 = 10'd634;
b_exp0 = 10'd817; b_exp1 = 10'd416; b_exp2 = 10'd747; b_exp3 = 10'd289;
a_sign0 = 4'd11; a_sign1 = 4'd2; a_sign2 = 4'd11; a_sign3 = 4'd3;
b_sign0 = 4'd13; b_sign1 = 4'd0; b_sign2 = 4'd13; b_sign3 = 4'd6;
@(posedge clk_i);
a_mant0 = 8'd228; a_mant1 = 8'd213; a_mant2 = 8'd177; a_mant3 = 8'd181;
b_mant0 = 8'd128; b_mant1 = 8'd185; b_mant2 = 8'd151; b_mant3 = 8'd117;
a_exp0 = 10'd36; a_exp1 = 10'd846; a_exp2 = 10'd274; a_exp3 = 10'd615;
b_exp0 = 10'd196; b_exp1 = 10'd940; b_exp2 = 10'd882; b_exp3 = 10'd125;
a_sign0 = 4'd4; a_sign1 = 4'd14; a_sign2 = 4'd8; a_sign3 = 4'd3;
b_sign0 = 4'd13; b_sign1 = 4'd12; b_sign2 = 4'd10; b_sign3 = 4'd1;
@(posedge clk_i);
a_mant0 = 8'd159; a_mant1 = 8'd147; a_mant2 = 8'd24; a_mant3 = 8'd212;
b_mant0 = 8'd191; b_mant1 = 8'd46; b_mant2 = 8'd99; b_mant3 = 8'd192;
a_exp0 = 10'd93; a_exp1 = 10'd776; a_exp2 = 10'd206; a_exp3 = 10'd65;
b_exp0 = 10'd319; b_exp1 = 10'd841; b_exp2 = 10'd537; b_exp3 = 10'd706;
a_sign0 = 4'd4; a_sign1 = 4'd3; a_sign2 = 4'd6; a_sign3 = 4'd8;
b_sign0 = 4'd10; b_sign1 = 4'd12; b_sign2 = 4'd10; b_sign3 = 4'd5;
@(posedge clk_i);
a_mant0 = 8'd12; a_mant1 = 8'd93; a_mant2 = 8'd210; a_mant3 = 8'd200;
b_mant0 = 8'd63; b_mant1 = 8'd81; b_mant2 = 8'd37; b_mant3 = 8'd79;
a_exp0 = 10'd755; a_exp1 = 10'd67; a_exp2 = 10'd467; a_exp3 = 10'd148;
b_exp0 = 10'd735; b_exp1 = 10'd888; b_exp2 = 10'd219; b_exp3 = 10'd817;
a_sign0 = 4'd10; a_sign1 = 4'd7; a_sign2 = 4'd0; a_sign3 = 4'd12;
b_sign0 = 4'd2; b_sign1 = 4'd11; b_sign2 = 4'd2; b_sign3 = 4'd3;
@(posedge clk_i);
a_mant0 = 8'd95; a_mant1 = 8'd179; a_mant2 = 8'd242; a_mant3 = 8'd239;
b_mant0 = 8'd60; b_mant1 = 8'd130; b_mant2 = 8'd82; b_mant3 = 8'd117;
a_exp0 = 10'd183; a_exp1 = 10'd326; a_exp2 = 10'd542; a_exp3 = 10'd266;
b_exp0 = 10'd819; b_exp1 = 10'd288; b_exp2 = 10'd747; b_exp3 = 10'd882;
a_sign0 = 4'd6; a_sign1 = 4'd10; a_sign2 = 4'd16; a_sign3 = 4'd9;
b_sign0 = 4'd5; b_sign1 = 4'd1; b_sign2 = 4'd14; b_sign3 = 4'd14;
@(posedge clk_i);
shared_exps0 = 8'd140;
shared_exps1 = 8'd121;
a_mant0 = 8'd237; a_mant1 = 8'd203; a_mant2 = 8'd160; a_mant3 = 8'd19;
b_mant0 = 8'd6; b_mant1 = 8'd51; b_mant2 = 8'd59; b_mant3 = 8'd148;
a_exp0 = 10'd320; a_exp1 = 10'd289; a_exp2 = 10'd798; a_exp3 = 10'd283;
b_exp0 = 10'd258; b_exp1 = 10'd717; b_exp2 = 10'd257; b_exp3 = 10'd612;
a_sign0 = 4'd16; a_sign1 = 4'd16; a_sign2 = 4'd13; a_sign3 = 4'd3;
b_sign0 = 4'd0; b_sign1 = 4'd13; b_sign2 = 4'd3; b_sign3 = 4'd14;
@(posedge clk_i);
a_mant0 = 8'd88; a_mant1 = 8'd172; a_mant2 = 8'd66; a_mant3 = 8'd164;
b_mant0 = 8'd96; b_mant1 = 8'd166; b_mant2 = 8'd106; b_mant3 = 8'd40;
a_exp0 = 10'd543; a_exp1 = 10'd790; a_exp2 = 10'd316; a_exp3 = 10'd375;
b_exp0 = 10'd686; b_exp1 = 10'd626; b_exp2 = 10'd1; b_exp3 = 10'd1009;
a_sign0 = 4'd12; a_sign1 = 4'd10; a_sign2 = 4'd9; a_sign3 = 4'd16;
b_sign0 = 4'd8; b_sign1 = 4'd4; b_sign2 = 4'd11; b_sign3 = 4'd16;
@(posedge clk_i);
a_mant0 = 8'd19; a_mant1 = 8'd31; a_mant2 = 8'd245; a_mant3 = 8'd121;
b_mant0 = 8'd77; b_mant1 = 8'd158; b_mant2 = 8'd210; b_mant3 = 8'd177;
a_exp0 = 10'd185; a_exp1 = 10'd468; a_exp2 = 10'd227; a_exp3 = 10'd0;
b_exp0 = 10'd956; b_exp1 = 10'd1008; b_exp2 = 10'd752; b_exp3 = 10'd933;
a_sign0 = 4'd10; a_sign1 = 4'd16; a_sign2 = 4'd11; a_sign3 = 4'd3;
b_sign0 = 4'd4; b_sign1 = 4'd0; b_sign2 = 4'd8; b_sign3 = 4'd16;
@(posedge clk_i);
a_mant0 = 8'd191; a_mant1 = 8'd23; a_mant2 = 8'd228; a_mant3 = 8'd127;
b_mant0 = 8'd13; b_mant1 = 8'd140; b_mant2 = 8'd43; b_mant3 = 8'd17;
a_exp0 = 10'd563; a_exp1 = 10'd990; a_exp2 = 10'd824; a_exp3 = 10'd632;
b_exp0 = 10'd291; b_exp1 = 10'd797; b_exp2 = 10'd351; b_exp3 = 10'd687;
a_sign0 = 4'd5; a_sign1 = 4'd11; a_sign2 = 4'd12; a_sign3 = 4'd3;
b_sign0 = 4'd9; b_sign1 = 4'd8; b_sign2 = 4'd15; b_sign3 = 4'd3;
@(posedge clk_i);
a_mant0 = 8'd52; a_mant1 = 8'd105; a_mant2 = 8'd254; a_mant3 = 8'd103;
b_mant0 = 8'd214; b_mant1 = 8'd131; b_mant2 = 8'd16; b_mant3 = 8'd135;
a_exp0 = 10'd915; a_exp1 = 10'd551; a_exp2 = 10'd642; a_exp3 = 10'd675;
b_exp0 = 10'd714; b_exp1 = 10'd63; b_exp2 = 10'd465; b_exp3 = 10'd802;
a_sign0 = 4'd0; a_sign1 = 4'd8; a_sign2 = 4'd10; a_sign3 = 4'd3;
b_sign0 = 4'd3; b_sign1 = 4'd10; b_sign2 = 4'd14; b_sign3 = 4'd7;
@(posedge clk_i);
a_mant0 = 8'd181; a_mant1 = 8'd171; a_mant2 = 8'd104; a_mant3 = 8'd168;
b_mant0 = 8'd178; b_mant1 = 8'd217; b_mant2 = 8'd29; b_mant3 = 8'd193;
a_exp0 = 10'd331; a_exp1 = 10'd598; a_exp2 = 10'd208; a_exp3 = 10'd883;
b_exp0 = 10'd107; b_exp1 = 10'd758; b_exp2 = 10'd120; b_exp3 = 10'd395;
a_sign0 = 4'd0; a_sign1 = 4'd15; a_sign2 = 4'd3; a_sign3 = 4'd5;
b_sign0 = 4'd16; b_sign1 = 4'd12; b_sign2 = 4'd3; b_sign3 = 4'd15;
@(posedge clk_i);
a_mant0 = 8'd210; a_mant1 = 8'd74; a_mant2 = 8'd74; a_mant3 = 8'd197;
b_mant0 = 8'd210; b_mant1 = 8'd5; b_mant2 = 8'd81; b_mant3 = 8'd206;
a_exp0 = 10'd118; a_exp1 = 10'd31; a_exp2 = 10'd774; a_exp3 = 10'd355;
b_exp0 = 10'd180; b_exp1 = 10'd96; b_exp2 = 10'd623; b_exp3 = 10'd806;
a_sign0 = 4'd15; a_sign1 = 4'd1; a_sign2 = 4'd1; a_sign3 = 4'd2;
b_sign0 = 4'd11; b_sign1 = 4'd3; b_sign2 = 4'd6; b_sign3 = 4'd2;
@(posedge clk_i);
a_mant0 = 8'd53; a_mant1 = 8'd21; a_mant2 = 8'd112; a_mant3 = 8'd73;
b_mant0 = 8'd198; b_mant1 = 8'd56; b_mant2 = 8'd111; b_mant3 = 8'd1;
a_exp0 = 10'd198; a_exp1 = 10'd527; a_exp2 = 10'd198; a_exp3 = 10'd106;
b_exp0 = 10'd743; b_exp1 = 10'd961; b_exp2 = 10'd996; b_exp3 = 10'd742;
a_sign0 = 4'd3; a_sign1 = 4'd4; a_sign2 = 4'd11; a_sign3 = 4'd6;
b_sign0 = 4'd8; b_sign1 = 4'd3; b_sign2 = 4'd14; b_sign3 = 4'd13;
@(posedge clk_i);
shared_exps0 = 8'd127;
shared_exps1 = 8'd129;
a_mant0 = 8'd17; a_mant1 = 8'd206; a_mant2 = 8'd189; a_mant3 = 8'd157;
b_mant0 = 8'd83; b_mant1 = 8'd251; b_mant2 = 8'd81; b_mant3 = 8'd44;
a_exp0 = 10'd590; a_exp1 = 10'd576; a_exp2 = 10'd468; a_exp3 = 10'd358;
b_exp0 = 10'd675; b_exp1 = 10'd14; b_exp2 = 10'd67; b_exp3 = 10'd489;
a_sign0 = 4'd8; a_sign1 = 4'd13; a_sign2 = 4'd12; a_sign3 = 4'd7;
b_sign0 = 4'd4; b_sign1 = 4'd15; b_sign2 = 4'd15; b_sign3 = 4'd7;
@(posedge clk_i);
a_mant0 = 8'd81; a_mant1 = 8'd74; a_mant2 = 8'd125; a_mant3 = 8'd198;
b_mant0 = 8'd156; b_mant1 = 8'd53; b_mant2 = 8'd90; b_mant3 = 8'd14;
a_exp0 = 10'd353; a_exp1 = 10'd765; a_exp2 = 10'd562; a_exp3 = 10'd996;
b_exp0 = 10'd334; b_exp1 = 10'd647; b_exp2 = 10'd112; b_exp3 = 10'd455;
a_sign0 = 4'd0; a_sign1 = 4'd5; a_sign2 = 4'd7; a_sign3 = 4'd3;
b_sign0 = 4'd4; b_sign1 = 4'd7; b_sign2 = 4'd16; b_sign3 = 4'd14;
@(posedge clk_i);
a_mant0 = 8'd154; a_mant1 = 8'd12; a_mant2 = 8'd120; a_mant3 = 8'd42;
b_mant0 = 8'd24; b_mant1 = 8'd139; b_mant2 = 8'd120; b_mant3 = 8'd152;
a_exp0 = 10'd21; a_exp1 = 10'd836; a_exp2 = 10'd404; a_exp3 = 10'd73;
b_exp0 = 10'd864; b_exp1 = 10'd635; b_exp2 = 10'd512; b_exp3 = 10'd867;
a_sign0 = 4'd13; a_sign1 = 4'd4; a_sign2 = 4'd3; a_sign3 = 4'd6;
b_sign0 = 4'd16; b_sign1 = 4'd4; b_sign2 = 4'd8; b_sign3 = 4'd5;
@(posedge clk_i);
a_mant0 = 8'd165; a_mant1 = 8'd92; a_mant2 = 8'd131; a_mant3 = 8'd104;
b_mant0 = 8'd19; b_mant1 = 8'd173; b_mant2 = 8'd208; b_mant3 = 8'd49;
a_exp0 = 10'd216; a_exp1 = 10'd498; a_exp2 = 10'd85; a_exp3 = 10'd460;
b_exp0 = 10'd138; b_exp1 = 10'd609; b_exp2 = 10'd208; b_exp3 = 10'd360;
a_sign0 = 4'd16; a_sign1 = 4'd14; a_sign2 = 4'd13; a_sign3 = 4'd2;
b_sign0 = 4'd0; b_sign1 = 4'd14; b_sign2 = 4'd14; b_sign3 = 4'd0;
@(posedge clk_i);
a_mant0 = 8'd158; a_mant1 = 8'd83; a_mant2 = 8'd124; a_mant3 = 8'd94;
b_mant0 = 8'd174; b_mant1 = 8'd68; b_mant2 = 8'd200; b_mant3 = 8'd206;
a_exp0 = 10'd436; a_exp1 = 10'd291; a_exp2 = 10'd2; a_exp3 = 10'd85;
b_exp0 = 10'd37; b_exp1 = 10'd907; b_exp2 = 10'd781; b_exp3 = 10'd853;
a_sign0 = 4'd2; a_sign1 = 4'd11; a_sign2 = 4'd14; a_sign3 = 4'd14;
b_sign0 = 4'd8; b_sign1 = 4'd8; b_sign2 = 4'd5; b_sign3 = 4'd7;
@(posedge clk_i);
a_mant0 = 8'd155; a_mant1 = 8'd125; a_mant2 = 8'd28; a_mant3 = 8'd172;
b_mant0 = 8'd121; b_mant1 = 8'd2; b_mant2 = 8'd164; b_mant3 = 8'd213;
a_exp0 = 10'd648; a_exp1 = 10'd681; a_exp2 = 10'd382; a_exp3 = 10'd600;
b_exp0 = 10'd525; b_exp1 = 10'd760; b_exp2 = 10'd569; b_exp3 = 10'd724;
a_sign0 = 4'd2; a_sign1 = 4'd13; a_sign2 = 4'd1; a_sign3 = 4'd0;
b_sign0 = 4'd10; b_sign1 = 4'd3; b_sign2 = 4'd8; b_sign3 = 4'd13;
@(posedge clk_i);
a_mant0 = 8'd41; a_mant1 = 8'd199; a_mant2 = 8'd107; a_mant3 = 8'd60;
b_mant0 = 8'd185; b_mant1 = 8'd63; b_mant2 = 8'd40; b_mant3 = 8'd88;
a_exp0 = 10'd450; a_exp1 = 10'd462; a_exp2 = 10'd353; a_exp3 = 10'd771;
b_exp0 = 10'd702; b_exp1 = 10'd257; b_exp2 = 10'd723; b_exp3 = 10'd646;
a_sign0 = 4'd13; a_sign1 = 4'd8; a_sign2 = 4'd13; a_sign3 = 4'd2;
b_sign0 = 4'd9; b_sign1 = 4'd4; b_sign2 = 4'd13; b_sign3 = 4'd2;
@(posedge clk_i);
a_mant0 = 8'd149; a_mant1 = 8'd102; a_mant2 = 8'd182; a_mant3 = 8'd26;
b_mant0 = 8'd204; b_mant1 = 8'd223; b_mant2 = 8'd106; b_mant3 = 8'd218;
a_exp0 = 10'd729; a_exp1 = 10'd655; a_exp2 = 10'd195; a_exp3 = 10'd418;
b_exp0 = 10'd622; b_exp1 = 10'd102; b_exp2 = 10'd630; b_exp3 = 10'd649;
a_sign0 = 4'd14; a_sign1 = 4'd1; a_sign2 = 4'd12; a_sign3 = 4'd9;
b_sign0 = 4'd11; b_sign1 = 4'd12; b_sign2 = 4'd11; b_sign3 = 4'd6;
@(posedge clk_i);
shared_exps0 = 8'd146;
shared_exps1 = 8'd144;
rstn = 0;
@(posedge clk_i);
rstn = 1;
a_mant0 = 8'd17; a_mant1 = 8'd3; a_mant2 = 8'd245; a_mant3 = 8'd198;
b_mant0 = 8'd184; b_mant1 = 8'd184; b_mant2 = 8'd127; b_mant3 = 8'd106;
a_exp0 = 10'd978; a_exp1 = 10'd104; a_exp2 = 10'd477; a_exp3 = 10'd415;
b_exp0 = 10'd690; b_exp1 = 10'd945; b_exp2 = 10'd110; b_exp3 = 10'd115;
a_sign0 = 4'd7; a_sign1 = 4'd9; a_sign2 = 4'd6; a_sign3 = 4'd5;
b_sign0 = 4'd8; b_sign1 = 4'd1; b_sign2 = 4'd11; b_sign3 = 4'd9;
@(posedge clk_i);
a_mant0 = 8'd157; a_mant1 = 8'd35; a_mant2 = 8'd5; a_mant3 = 8'd104;
b_mant0 = 8'd116; b_mant1 = 8'd60; b_mant2 = 8'd133; b_mant3 = 8'd31;
a_exp0 = 10'd799; a_exp1 = 10'd288; a_exp2 = 10'd313; a_exp3 = 10'd825;
b_exp0 = 10'd689; b_exp1 = 10'd910; b_exp2 = 10'd203; b_exp3 = 10'd1022;
a_sign0 = 4'd10; a_sign1 = 4'd0; a_sign2 = 4'd15; a_sign3 = 4'd1;
b_sign0 = 4'd9; b_sign1 = 4'd6; b_sign2 = 4'd1; b_sign3 = 4'd5;
@(posedge clk_i);
a_mant0 = 8'd138; a_mant1 = 8'd49; a_mant2 = 8'd130; a_mant3 = 8'd228;
b_mant0 = 8'd195; b_mant1 = 8'd189; b_mant2 = 8'd18; b_mant3 = 8'd203;
a_exp0 = 10'd758; a_exp1 = 10'd350; a_exp2 = 10'd427; a_exp3 = 10'd107;
b_exp0 = 10'd212; b_exp1 = 10'd921; b_exp2 = 10'd427; b_exp3 = 10'd189;
a_sign0 = 4'd16; a_sign1 = 4'd9; a_sign2 = 4'd6; a_sign3 = 4'd0;
b_sign0 = 4'd4; b_sign1 = 4'd16; b_sign2 = 4'd11; b_sign3 = 4'd7;
@(posedge clk_i);
a_mant0 = 8'd0; a_mant1 = 8'd218; a_mant2 = 8'd198; a_mant3 = 8'd241;
b_mant0 = 8'd231; b_mant1 = 8'd52; b_mant2 = 8'd54; b_mant3 = 8'd91;
a_exp0 = 10'd634; a_exp1 = 10'd456; a_exp2 = 10'd196; a_exp3 = 10'd15;
b_exp0 = 10'd630; b_exp1 = 10'd204; b_exp2 = 10'd911; b_exp3 = 10'd156;
a_sign0 = 4'd14; a_sign1 = 4'd15; a_sign2 = 4'd14; a_sign3 = 4'd6;
b_sign0 = 4'd15; b_sign1 = 4'd0; b_sign2 = 4'd13; b_sign3 = 4'd9;
@(posedge clk_i);
a_mant0 = 8'd163; a_mant1 = 8'd128; a_mant2 = 8'd58; a_mant3 = 8'd100;
b_mant0 = 8'd109; b_mant1 = 8'd239; b_mant2 = 8'd156; b_mant3 = 8'd211;
a_exp0 = 10'd930; a_exp1 = 10'd835; a_exp2 = 10'd738; a_exp3 = 10'd635;
b_exp0 = 10'd483; b_exp1 = 10'd864; b_exp2 = 10'd283; b_exp3 = 10'd1004;
a_sign0 = 4'd15; a_sign1 = 4'd12; a_sign2 = 4'd5; a_sign3 = 4'd2;
b_sign0 = 4'd8; b_sign1 = 4'd8; b_sign2 = 4'd8; b_sign3 = 4'd4;
@(posedge clk_i);
a_mant0 = 8'd17; a_mant1 = 8'd115; a_mant2 = 8'd72; a_mant3 = 8'd40;
b_mant0 = 8'd152; b_mant1 = 8'd245; b_mant2 = 8'd222; b_mant3 = 8'd137;
a_exp0 = 10'd371; a_exp1 = 10'd826; a_exp2 = 10'd298; a_exp3 = 10'd393;
b_exp0 = 10'd130; b_exp1 = 10'd112; b_exp2 = 10'd560; b_exp3 = 10'd971;
a_sign0 = 4'd1; a_sign1 = 4'd5; a_sign2 = 4'd4; a_sign3 = 4'd15;
b_sign0 = 4'd13; b_sign1 = 4'd7; b_sign2 = 4'd14; b_sign3 = 4'd4;
@(posedge clk_i);
a_mant0 = 8'd85; a_mant1 = 8'd82; a_mant2 = 8'd236; a_mant3 = 8'd140;
b_mant0 = 8'd142; b_mant1 = 8'd192; b_mant2 = 8'd149; b_mant3 = 8'd15;
a_exp0 = 10'd470; a_exp1 = 10'd337; a_exp2 = 10'd530; a_exp3 = 10'd640;
b_exp0 = 10'd437; b_exp1 = 10'd676; b_exp2 = 10'd464; b_exp3 = 10'd796;
a_sign0 = 4'd14; a_sign1 = 4'd10; a_sign2 = 4'd10; a_sign3 = 4'd2;
b_sign0 = 4'd10; b_sign1 = 4'd8; b_sign2 = 4'd12; b_sign3 = 4'd1;
@(posedge clk_i);
shared_exps0 = 8'd118;
shared_exps1 = 8'd151;
a_mant0 = 8'd101; a_mant1 = 8'd186; a_mant2 = 8'd99; a_mant3 = 8'd57;
b_mant0 = 8'd126; b_mant1 = 8'd74; b_mant2 = 8'd32; b_mant3 = 8'd115;
a_exp0 = 10'd487; a_exp1 = 10'd371; a_exp2 = 10'd570; a_exp3 = 10'd346;
b_exp0 = 10'd0; b_exp1 = 10'd206; b_exp2 = 10'd815; b_exp3 = 10'd223;
a_sign0 = 4'd7; a_sign1 = 4'd12; a_sign2 = 4'd7; a_sign3 = 4'd4;
b_sign0 = 4'd5; b_sign1 = 4'd10; b_sign2 = 4'd14; b_sign3 = 4'd12;
@(posedge clk_i);
a_mant0 = 8'd168; a_mant1 = 8'd70; a_mant2 = 8'd132; a_mant3 = 8'd225;
b_mant0 = 8'd52; b_mant1 = 8'd254; b_mant2 = 8'd223; b_mant3 = 8'd208;
a_exp0 = 10'd565; a_exp1 = 10'd757; a_exp2 = 10'd55; a_exp3 = 10'd975;
b_exp0 = 10'd689; b_exp1 = 10'd648; b_exp2 = 10'd108; b_exp3 = 10'd420;
a_sign0 = 4'd3; a_sign1 = 4'd6; a_sign2 = 4'd1; a_sign3 = 4'd4;
b_sign0 = 4'd14; b_sign1 = 4'd6; b_sign2 = 4'd0; b_sign3 = 4'd12;
@(posedge clk_i);
a_mant0 = 8'd136; a_mant1 = 8'd120; a_mant2 = 8'd2; a_mant3 = 8'd33;
b_mant0 = 8'd33; b_mant1 = 8'd149; b_mant2 = 8'd56; b_mant3 = 8'd167;
a_exp0 = 10'd149; a_exp1 = 10'd987; a_exp2 = 10'd107; a_exp3 = 10'd901;
b_exp0 = 10'd211; b_exp1 = 10'd486; b_exp2 = 10'd941; b_exp3 = 10'd458;
a_sign0 = 4'd9; a_sign1 = 4'd12; a_sign2 = 4'd13; a_sign3 = 4'd5;
b_sign0 = 4'd6; b_sign1 = 4'd9; b_sign2 = 4'd4; b_sign3 = 4'd7;
@(posedge clk_i);
a_mant0 = 8'd255; a_mant1 = 8'd85; a_mant2 = 8'd48; a_mant3 = 8'd219;
b_mant0 = 8'd221; b_mant1 = 8'd151; b_mant2 = 8'd56; b_mant3 = 8'd14;
a_exp0 = 10'd543; a_exp1 = 10'd536; a_exp2 = 10'd831; a_exp3 = 10'd6;
b_exp0 = 10'd600; b_exp1 = 10'd857; b_exp2 = 10'd285; b_exp3 = 10'd1016;
a_sign0 = 4'd14; a_sign1 = 4'd7; a_sign2 = 4'd11; a_sign3 = 4'd2;
b_sign0 = 4'd14; b_sign1 = 4'd12; b_sign2 = 4'd11; b_sign3 = 4'd9;
@(posedge clk_i);
a_mant0 = 8'd21; a_mant1 = 8'd120; a_mant2 = 8'd106; a_mant3 = 8'd51;
b_mant0 = 8'd134; b_mant1 = 8'd26; b_mant2 = 8'd44; b_mant3 = 8'd67;
a_exp0 = 10'd895; a_exp1 = 10'd745; a_exp2 = 10'd461; a_exp3 = 10'd390;
b_exp0 = 10'd726; b_exp1 = 10'd676; b_exp2 = 10'd588; b_exp3 = 10'd57;
a_sign0 = 4'd9; a_sign1 = 4'd16; a_sign2 = 4'd4; a_sign3 = 4'd13;
b_sign0 = 4'd13; b_sign1 = 4'd6; b_sign2 = 4'd1; b_sign3 = 4'd5;
@(posedge clk_i);
a_mant0 = 8'd202; a_mant1 = 8'd152; a_mant2 = 8'd103; a_mant3 = 8'd208;
b_mant0 = 8'd238; b_mant1 = 8'd76; b_mant2 = 8'd188; b_mant3 = 8'd169;
a_exp0 = 10'd942; a_exp1 = 10'd668; a_exp2 = 10'd394; a_exp3 = 10'd948;
b_exp0 = 10'd693; b_exp1 = 10'd869; b_exp2 = 10'd538; b_exp3 = 10'd26;
a_sign0 = 4'd4; a_sign1 = 4'd15; a_sign2 = 4'd6; a_sign3 = 4'd2;
b_sign0 = 4'd8; b_sign1 = 4'd4; b_sign2 = 4'd1; b_sign3 = 4'd9;
@(posedge clk_i);
a_mant0 = 8'd194; a_mant1 = 8'd151; a_mant2 = 8'd144; a_mant3 = 8'd123;
b_mant0 = 8'd166; b_mant1 = 8'd101; b_mant2 = 8'd198; b_mant3 = 8'd108;
a_exp0 = 10'd94; a_exp1 = 10'd867; a_exp2 = 10'd736; a_exp3 = 10'd47;
b_exp0 = 10'd804; b_exp1 = 10'd68; b_exp2 = 10'd528; b_exp3 = 10'd4;
a_sign0 = 4'd6; a_sign1 = 4'd2; a_sign2 = 4'd1; a_sign3 = 4'd0;
b_sign0 = 4'd12; b_sign1 = 4'd12; b_sign2 = 4'd14; b_sign3 = 4'd15;
@(posedge clk_i);
a_mant0 = 8'd40; a_mant1 = 8'd83; a_mant2 = 8'd115; a_mant3 = 8'd195;
b_mant0 = 8'd114; b_mant1 = 8'd123; b_mant2 = 8'd192; b_mant3 = 8'd214;
a_exp0 = 10'd565; a_exp1 = 10'd723; a_exp2 = 10'd339; a_exp3 = 10'd310;
b_exp0 = 10'd257; b_exp1 = 10'd406; b_exp2 = 10'd834; b_exp3 = 10'd188;
a_sign0 = 4'd5; a_sign1 = 4'd2; a_sign2 = 4'd5; a_sign3 = 4'd16;
b_sign0 = 4'd8; b_sign1 = 4'd11; b_sign2 = 4'd6; b_sign3 = 4'd15;
@(posedge clk_i);
shared_exps0 = 8'd136;
shared_exps1 = 8'd119;
a_mant0 = 8'd225; a_mant1 = 8'd20; a_mant2 = 8'd226; a_mant3 = 8'd85;
b_mant0 = 8'd128; b_mant1 = 8'd218; b_mant2 = 8'd11; b_mant3 = 8'd134;
a_exp0 = 10'd23; a_exp1 = 10'd728; a_exp2 = 10'd528; a_exp3 = 10'd1017;
b_exp0 = 10'd27; b_exp1 = 10'd236; b_exp2 = 10'd102; b_exp3 = 10'd577;
a_sign0 = 4'd7; a_sign1 = 4'd15; a_sign2 = 4'd12; a_sign3 = 4'd14;
b_sign0 = 4'd15; b_sign1 = 4'd8; b_sign2 = 4'd15; b_sign3 = 4'd14;
@(posedge clk_i);
a_mant0 = 8'd163; a_mant1 = 8'd212; a_mant2 = 8'd88; a_mant3 = 8'd248;
b_mant0 = 8'd148; b_mant1 = 8'd223; b_mant2 = 8'd203; b_mant3 = 8'd109;
a_exp0 = 10'd1020; a_exp1 = 10'd62; a_exp2 = 10'd457; a_exp3 = 10'd781;
b_exp0 = 10'd717; b_exp1 = 10'd702; b_exp2 = 10'd851; b_exp3 = 10'd435;
a_sign0 = 4'd13; a_sign1 = 4'd5; a_sign2 = 4'd11; a_sign3 = 4'd3;
b_sign0 = 4'd4; b_sign1 = 4'd3; b_sign2 = 4'd8; b_sign3 = 4'd7;
@(posedge clk_i);
a_mant0 = 8'd104; a_mant1 = 8'd132; a_mant2 = 8'd194; a_mant3 = 8'd249;
b_mant0 = 8'd244; b_mant1 = 8'd88; b_mant2 = 8'd24; b_mant3 = 8'd19;
a_exp0 = 10'd488; a_exp1 = 10'd94; a_exp2 = 10'd164; a_exp3 = 10'd625;
b_exp0 = 10'd803; b_exp1 = 10'd298; b_exp2 = 10'd539; b_exp3 = 10'd108;
a_sign0 = 4'd12; a_sign1 = 4'd6; a_sign2 = 4'd15; a_sign3 = 4'd7;
b_sign0 = 4'd0; b_sign1 = 4'd11; b_sign2 = 4'd3; b_sign3 = 4'd1;
@(posedge clk_i);
a_mant0 = 8'd104; a_mant1 = 8'd42; a_mant2 = 8'd208; a_mant3 = 8'd178;
b_mant0 = 8'd101; b_mant1 = 8'd206; b_mant2 = 8'd83; b_mant3 = 8'd185;
a_exp0 = 10'd575; a_exp1 = 10'd466; a_exp2 = 10'd643; a_exp3 = 10'd355;
b_exp0 = 10'd659; b_exp1 = 10'd251; b_exp2 = 10'd84; b_exp3 = 10'd773;
a_sign0 = 4'd5; a_sign1 = 4'd13; a_sign2 = 4'd3; a_sign3 = 4'd1;
b_sign0 = 4'd7; b_sign1 = 4'd8; b_sign2 = 4'd8; b_sign3 = 4'd16;
@(posedge clk_i);
a_mant0 = 8'd211; a_mant1 = 8'd165; a_mant2 = 8'd231; a_mant3 = 8'd80;
b_mant0 = 8'd101; b_mant1 = 8'd245; b_mant2 = 8'd4; b_mant3 = 8'd55;
a_exp0 = 10'd552; a_exp1 = 10'd708; a_exp2 = 10'd934; a_exp3 = 10'd906;
b_exp0 = 10'd91; b_exp1 = 10'd179; b_exp2 = 10'd265; b_exp3 = 10'd271;
a_sign0 = 4'd6; a_sign1 = 4'd1; a_sign2 = 4'd15; a_sign3 = 4'd11;
b_sign0 = 4'd1; b_sign1 = 4'd9; b_sign2 = 4'd12; b_sign3 = 4'd2;
@(posedge clk_i);
a_mant0 = 8'd107; a_mant1 = 8'd158; a_mant2 = 8'd217; a_mant3 = 8'd240;
b_mant0 = 8'd15; b_mant1 = 8'd115; b_mant2 = 8'd20; b_mant3 = 8'd57;
a_exp0 = 10'd899; a_exp1 = 10'd228; a_exp2 = 10'd38; a_exp3 = 10'd810;
b_exp0 = 10'd14; b_exp1 = 10'd647; b_exp2 = 10'd500; b_exp3 = 10'd100;
a_sign0 = 4'd6; a_sign1 = 4'd6; a_sign2 = 4'd0; a_sign3 = 4'd4;
b_sign0 = 4'd13; b_sign1 = 4'd15; b_sign2 = 4'd14; b_sign3 = 4'd4;
@(posedge clk_i);
a_mant0 = 8'd181; a_mant1 = 8'd137; a_mant2 = 8'd166; a_mant3 = 8'd141;
b_mant0 = 8'd146; b_mant1 = 8'd111; b_mant2 = 8'd83; b_mant3 = 8'd156;
a_exp0 = 10'd320; a_exp1 = 10'd281; a_exp2 = 10'd83; a_exp3 = 10'd663;
b_exp0 = 10'd16; b_exp1 = 10'd723; b_exp2 = 10'd344; b_exp3 = 10'd1020;
a_sign0 = 4'd16; a_sign1 = 4'd9; a_sign2 = 4'd12; a_sign3 = 4'd15;
b_sign0 = 4'd0; b_sign1 = 4'd7; b_sign2 = 4'd12; b_sign3 = 4'd11;
@(posedge clk_i);
a_mant0 = 8'd187; a_mant1 = 8'd0; a_mant2 = 8'd149; a_mant3 = 8'd144;
b_mant0 = 8'd167; b_mant1 = 8'd209; b_mant2 = 8'd191; b_mant3 = 8'd1;
a_exp0 = 10'd964; a_exp1 = 10'd568; a_exp2 = 10'd161; a_exp3 = 10'd59;
b_exp0 = 10'd228; b_exp1 = 10'd919; b_exp2 = 10'd299; b_exp3 = 10'd885;
a_sign0 = 4'd13; a_sign1 = 4'd4; a_sign2 = 4'd1; a_sign3 = 4'd7;
b_sign0 = 4'd3; b_sign1 = 4'd10; b_sign2 = 4'd16; b_sign3 = 4'd15;
@(posedge clk_i);
shared_exps0 = 8'd134;
shared_exps1 = 8'd142;
a_mant0 = 8'd133; a_mant1 = 8'd239; a_mant2 = 8'd39; a_mant3 = 8'd206;
b_mant0 = 8'd207; b_mant1 = 8'd87; b_mant2 = 8'd46; b_mant3 = 8'd78;
a_exp0 = 10'd683; a_exp1 = 10'd666; a_exp2 = 10'd366; a_exp3 = 10'd372;
b_exp0 = 10'd905; b_exp1 = 10'd839; b_exp2 = 10'd402; b_exp3 = 10'd742;
a_sign0 = 4'd12; a_sign1 = 4'd5; a_sign2 = 4'd5; a_sign3 = 4'd8;
b_sign0 = 4'd3; b_sign1 = 4'd5; b_sign2 = 4'd11; b_sign3 = 4'd7;
@(posedge clk_i);
a_mant0 = 8'd108; a_mant1 = 8'd51; a_mant2 = 8'd166; a_mant3 = 8'd132;
b_mant0 = 8'd71; b_mant1 = 8'd244; b_mant2 = 8'd119; b_mant3 = 8'd240;
a_exp0 = 10'd211; a_exp1 = 10'd513; a_exp2 = 10'd981; a_exp3 = 10'd289;
b_exp0 = 10'd217; b_exp1 = 10'd263; b_exp2 = 10'd153; b_exp3 = 10'd865;
a_sign0 = 4'd15; a_sign1 = 4'd14; a_sign2 = 4'd1; a_sign3 = 4'd9;
b_sign0 = 4'd2; b_sign1 = 4'd3; b_sign2 = 4'd5; b_sign3 = 4'd9;
@(posedge clk_i);
a_mant0 = 8'd97; a_mant1 = 8'd23; a_mant2 = 8'd59; a_mant3 = 8'd213;
b_mant0 = 8'd112; b_mant1 = 8'd234; b_mant2 = 8'd72; b_mant3 = 8'd178;
a_exp0 = 10'd248; a_exp1 = 10'd725; a_exp2 = 10'd970; a_exp3 = 10'd564;
b_exp0 = 10'd196; b_exp1 = 10'd824; b_exp2 = 10'd109; b_exp3 = 10'd583;
a_sign0 = 4'd3; a_sign1 = 4'd1; a_sign2 = 4'd2; a_sign3 = 4'd8;
b_sign0 = 4'd8; b_sign1 = 4'd8; b_sign2 = 4'd9; b_sign3 = 4'd13;
@(posedge clk_i);
a_mant0 = 8'd198; a_mant1 = 8'd16; a_mant2 = 8'd93; a_mant3 = 8'd37;
b_mant0 = 8'd183; b_mant1 = 8'd183; b_mant2 = 8'd114; b_mant3 = 8'd19;
a_exp0 = 10'd233; a_exp1 = 10'd508; a_exp2 = 10'd65; a_exp3 = 10'd387;
b_exp0 = 10'd244; b_exp1 = 10'd523; b_exp2 = 10'd69; b_exp3 = 10'd347;
a_sign0 = 4'd2; a_sign1 = 4'd13; a_sign2 = 4'd10; a_sign3 = 4'd4;
b_sign0 = 4'd10; b_sign1 = 4'd10; b_sign2 = 4'd6; b_sign3 = 4'd0;
@(posedge clk_i);
a_mant0 = 8'd171; a_mant1 = 8'd108; a_mant2 = 8'd57; a_mant3 = 8'd95;
b_mant0 = 8'd44; b_mant1 = 8'd231; b_mant2 = 8'd202; b_mant3 = 8'd241;
a_exp0 = 10'd971; a_exp1 = 10'd839; a_exp2 = 10'd968; a_exp3 = 10'd783;
b_exp0 = 10'd265; b_exp1 = 10'd461; b_exp2 = 10'd694; b_exp3 = 10'd420;
a_sign0 = 4'd2; a_sign1 = 4'd4; a_sign2 = 4'd1; a_sign3 = 4'd3;
b_sign0 = 4'd5; b_sign1 = 4'd8; b_sign2 = 4'd0; b_sign3 = 4'd14;
@(posedge clk_i);
a_mant0 = 8'd97; a_mant1 = 8'd86; a_mant2 = 8'd181; a_mant3 = 8'd124;
b_mant0 = 8'd182; b_mant1 = 8'd20; b_mant2 = 8'd109; b_mant3 = 8'd199;
a_exp0 = 10'd438; a_exp1 = 10'd890; a_exp2 = 10'd811; a_exp3 = 10'd739;
b_exp0 = 10'd355; b_exp1 = 10'd499; b_exp2 = 10'd638; b_exp3 = 10'd496;
a_sign0 = 4'd6; a_sign1 = 4'd10; a_sign2 = 4'd16; a_sign3 = 4'd5;
b_sign0 = 4'd1; b_sign1 = 4'd11; b_sign2 = 4'd3; b_sign3 = 4'd15;
@(posedge clk_i);
a_mant0 = 8'd76; a_mant1 = 8'd136; a_mant2 = 8'd205; a_mant3 = 8'd76;
b_mant0 = 8'd243; b_mant1 = 8'd180; b_mant2 = 8'd61; b_mant3 = 8'd234;
a_exp0 = 10'd78; a_exp1 = 10'd1001; a_exp2 = 10'd318; a_exp3 = 10'd906;
b_exp0 = 10'd455; b_exp1 = 10'd891; b_exp2 = 10'd943; b_exp3 = 10'd481;
a_sign0 = 4'd13; a_sign1 = 4'd16; a_sign2 = 4'd3; a_sign3 = 4'd9;
b_sign0 = 4'd11; b_sign1 = 4'd1; b_sign2 = 4'd6; b_sign3 = 4'd14;
@(posedge clk_i);
a_mant0 = 8'd173; a_mant1 = 8'd203; a_mant2 = 8'd11; a_mant3 = 8'd27;
b_mant0 = 8'd200; b_mant1 = 8'd254; b_mant2 = 8'd201; b_mant3 = 8'd189;
a_exp0 = 10'd693; a_exp1 = 10'd788; a_exp2 = 10'd327; a_exp3 = 10'd404;
b_exp0 = 10'd489; b_exp1 = 10'd890; b_exp2 = 10'd389; b_exp3 = 10'd274;
a_sign0 = 4'd16; a_sign1 = 4'd10; a_sign2 = 4'd14; a_sign3 = 4'd9;
b_sign0 = 4'd4; b_sign1 = 4'd0; b_sign2 = 4'd6; b_sign3 = 4'd15;
@(posedge clk_i);
shared_exps0 = 8'd111;
shared_exps1 = 8'd118;
rstn = 0;
@(posedge clk_i);
rstn = 1;
a_mant0 = 8'd188; a_mant1 = 8'd167; a_mant2 = 8'd169; a_mant3 = 8'd71;
b_mant0 = 8'd186; b_mant1 = 8'd241; b_mant2 = 8'd77; b_mant3 = 8'd121;
a_exp0 = 10'd300; a_exp1 = 10'd665; a_exp2 = 10'd465; a_exp3 = 10'd502;
b_exp0 = 10'd193; b_exp1 = 10'd396; b_exp2 = 10'd272; b_exp3 = 10'd500;
a_sign0 = 4'd0; a_sign1 = 4'd5; a_sign2 = 4'd3; a_sign3 = 4'd11;
b_sign0 = 4'd4; b_sign1 = 4'd16; b_sign2 = 4'd14; b_sign3 = 4'd5;
@(posedge clk_i);
a_mant0 = 8'd229; a_mant1 = 8'd118; a_mant2 = 8'd159; a_mant3 = 8'd75;
b_mant0 = 8'd179; b_mant1 = 8'd107; b_mant2 = 8'd200; b_mant3 = 8'd201;
a_exp0 = 10'd310; a_exp1 = 10'd105; a_exp2 = 10'd253; a_exp3 = 10'd227;
b_exp0 = 10'd126; b_exp1 = 10'd307; b_exp2 = 10'd301; b_exp3 = 10'd305;
a_sign0 = 4'd10; a_sign1 = 4'd0; a_sign2 = 4'd5; a_sign3 = 4'd5;
b_sign0 = 4'd14; b_sign1 = 4'd13; b_sign2 = 4'd6; b_sign3 = 4'd8;
@(posedge clk_i);
a_mant0 = 8'd172; a_mant1 = 8'd111; a_mant2 = 8'd66; a_mant3 = 8'd4;
b_mant0 = 8'd212; b_mant1 = 8'd113; b_mant2 = 8'd101; b_mant3 = 8'd85;
a_exp0 = 10'd833; a_exp1 = 10'd185; a_exp2 = 10'd915; a_exp3 = 10'd927;
b_exp0 = 10'd44; b_exp1 = 10'd40; b_exp2 = 10'd823; b_exp3 = 10'd764;
a_sign0 = 4'd0; a_sign1 = 4'd6; a_sign2 = 4'd1; a_sign3 = 4'd3;
b_sign0 = 4'd10; b_sign1 = 4'd12; b_sign2 = 4'd12; b_sign3 = 4'd14;
@(posedge clk_i);
a_mant0 = 8'd183; a_mant1 = 8'd70; a_mant2 = 8'd241; a_mant3 = 8'd46;
b_mant0 = 8'd177; b_mant1 = 8'd210; b_mant2 = 8'd205; b_mant3 = 8'd226;
a_exp0 = 10'd578; a_exp1 = 10'd501; a_exp2 = 10'd910; a_exp3 = 10'd990;
b_exp0 = 10'd484; b_exp1 = 10'd1023; b_exp2 = 10'd928; b_exp3 = 10'd375;
a_sign0 = 4'd15; a_sign1 = 4'd14; a_sign2 = 4'd6; a_sign3 = 4'd8;
b_sign0 = 4'd2; b_sign1 = 4'd15; b_sign2 = 4'd5; b_sign3 = 4'd16;
@(posedge clk_i);
a_mant0 = 8'd169; a_mant1 = 8'd82; a_mant2 = 8'd29; a_mant3 = 8'd147;
b_mant0 = 8'd63; b_mant1 = 8'd80; b_mant2 = 8'd8; b_mant3 = 8'd12;
a_exp0 = 10'd854; a_exp1 = 10'd658; a_exp2 = 10'd168; a_exp3 = 10'd721;
b_exp0 = 10'd153; b_exp1 = 10'd353; b_exp2 = 10'd433; b_exp3 = 10'd478;
a_sign0 = 4'd1; a_sign1 = 4'd15; a_sign2 = 4'd5; a_sign3 = 4'd9;
b_sign0 = 4'd8; b_sign1 = 4'd9; b_sign2 = 4'd4; b_sign3 = 4'd5;
@(posedge clk_i);
a_mant0 = 8'd47; a_mant1 = 8'd242; a_mant2 = 8'd88; a_mant3 = 8'd36;
b_mant0 = 8'd158; b_mant1 = 8'd67; b_mant2 = 8'd227; b_mant3 = 8'd233;
a_exp0 = 10'd1010; a_exp1 = 10'd598; a_exp2 = 10'd48; a_exp3 = 10'd122;
b_exp0 = 10'd117; b_exp1 = 10'd472; b_exp2 = 10'd679; b_exp3 = 10'd780;
a_sign0 = 4'd12; a_sign1 = 4'd7; a_sign2 = 4'd10; a_sign3 = 4'd14;
b_sign0 = 4'd11; b_sign1 = 4'd15; b_sign2 = 4'd11; b_sign3 = 4'd12;
@(posedge clk_i);
a_mant0 = 8'd100; a_mant1 = 8'd138; a_mant2 = 8'd153; a_mant3 = 8'd1;
b_mant0 = 8'd191; b_mant1 = 8'd12; b_mant2 = 8'd11; b_mant3 = 8'd165;
a_exp0 = 10'd219; a_exp1 = 10'd986; a_exp2 = 10'd273; a_exp3 = 10'd242;
b_exp0 = 10'd461; b_exp1 = 10'd777; b_exp2 = 10'd724; b_exp3 = 10'd48;
a_sign0 = 4'd5; a_sign1 = 4'd9; a_sign2 = 4'd15; a_sign3 = 4'd12;
b_sign0 = 4'd0; b_sign1 = 4'd7; b_sign2 = 4'd14; b_sign3 = 4'd8;
@(posedge clk_i);
shared_exps0 = 8'd133;
shared_exps1 = 8'd123;
a_mant0 = 8'd96; a_mant1 = 8'd205; a_mant2 = 8'd119; a_mant3 = 8'd141;
b_mant0 = 8'd63; b_mant1 = 8'd192; b_mant2 = 8'd45; b_mant3 = 8'd160;
a_exp0 = 10'd810; a_exp1 = 10'd149; a_exp2 = 10'd300; a_exp3 = 10'd505;
b_exp0 = 10'd838; b_exp1 = 10'd312; b_exp2 = 10'd78; b_exp3 = 10'd121;
a_sign0 = 4'd12; a_sign1 = 4'd9; a_sign2 = 4'd13; a_sign3 = 4'd9;
b_sign0 = 4'd9; b_sign1 = 4'd12; b_sign2 = 4'd8; b_sign3 = 4'd10;
@(posedge clk_i);
a_mant0 = 8'd121; a_mant1 = 8'd46; a_mant2 = 8'd52; a_mant3 = 8'd160;
b_mant0 = 8'd189; b_mant1 = 8'd186; b_mant2 = 8'd91; b_mant3 = 8'd215;
a_exp0 = 10'd174; a_exp1 = 10'd457; a_exp2 = 10'd695; a_exp3 = 10'd651;
b_exp0 = 10'd20; b_exp1 = 10'd524; b_exp2 = 10'd753; b_exp3 = 10'd676;
a_sign0 = 4'd9; a_sign1 = 4'd12; a_sign2 = 4'd7; a_sign3 = 4'd14;
b_sign0 = 4'd15; b_sign1 = 4'd8; b_sign2 = 4'd1; b_sign3 = 4'd15;
@(posedge clk_i);
a_mant0 = 8'd92; a_mant1 = 8'd203; a_mant2 = 8'd93; a_mant3 = 8'd80;
b_mant0 = 8'd90; b_mant1 = 8'd231; b_mant2 = 8'd23; b_mant3 = 8'd213;
a_exp0 = 10'd657; a_exp1 = 10'd853; a_exp2 = 10'd621; a_exp3 = 10'd976;
b_exp0 = 10'd739; b_exp1 = 10'd938; b_exp2 = 10'd227; b_exp3 = 10'd751;
a_sign0 = 4'd14; a_sign1 = 4'd11; a_sign2 = 4'd10; a_sign3 = 4'd12;
b_sign0 = 4'd15; b_sign1 = 4'd2; b_sign2 = 4'd9; b_sign3 = 4'd16;
@(posedge clk_i);
a_mant0 = 8'd31; a_mant1 = 8'd171; a_mant2 = 8'd244; a_mant3 = 8'd10;
b_mant0 = 8'd163; b_mant1 = 8'd91; b_mant2 = 8'd62; b_mant3 = 8'd253;
a_exp0 = 10'd235; a_exp1 = 10'd684; a_exp2 = 10'd572; a_exp3 = 10'd86;
b_exp0 = 10'd271; b_exp1 = 10'd734; b_exp2 = 10'd689; b_exp3 = 10'd557;
a_sign0 = 4'd2; a_sign1 = 4'd9; a_sign2 = 4'd1; a_sign3 = 4'd6;
b_sign0 = 4'd16; b_sign1 = 4'd14; b_sign2 = 4'd15; b_sign3 = 4'd5;
@(posedge clk_i);
a_mant0 = 8'd121; a_mant1 = 8'd89; a_mant2 = 8'd151; a_mant3 = 8'd72;
b_mant0 = 8'd104; b_mant1 = 8'd166; b_mant2 = 8'd111; b_mant3 = 8'd186;
a_exp0 = 10'd319; a_exp1 = 10'd962; a_exp2 = 10'd270; a_exp3 = 10'd64;
b_exp0 = 10'd364; b_exp1 = 10'd720; b_exp2 = 10'd300; b_exp3 = 10'd125;
a_sign0 = 4'd1; a_sign1 = 4'd0; a_sign2 = 4'd5; a_sign3 = 4'd9;
b_sign0 = 4'd16; b_sign1 = 4'd2; b_sign2 = 4'd15; b_sign3 = 4'd8;
@(posedge clk_i);
a_mant0 = 8'd176; a_mant1 = 8'd75; a_mant2 = 8'd159; a_mant3 = 8'd186;
b_mant0 = 8'd132; b_mant1 = 8'd31; b_mant2 = 8'd18; b_mant3 = 8'd181;
a_exp0 = 10'd726; a_exp1 = 10'd946; a_exp2 = 10'd785; a_exp3 = 10'd655;
b_exp0 = 10'd984; b_exp1 = 10'd997; b_exp2 = 10'd432; b_exp3 = 10'd1018;
a_sign0 = 4'd16; a_sign1 = 4'd6; a_sign2 = 4'd4; a_sign3 = 4'd11;
b_sign0 = 4'd15; b_sign1 = 4'd9; b_sign2 = 4'd14; b_sign3 = 4'd14;
@(posedge clk_i);
a_mant0 = 8'd219; a_mant1 = 8'd228; a_mant2 = 8'd166; a_mant3 = 8'd148;
b_mant0 = 8'd135; b_mant1 = 8'd50; b_mant2 = 8'd210; b_mant3 = 8'd249;
a_exp0 = 10'd834; a_exp1 = 10'd786; a_exp2 = 10'd743; a_exp3 = 10'd63;
b_exp0 = 10'd863; b_exp1 = 10'd1009; b_exp2 = 10'd42; b_exp3 = 10'd829;
a_sign0 = 4'd0; a_sign1 = 4'd8; a_sign2 = 4'd10; a_sign3 = 4'd14;
b_sign0 = 4'd9; b_sign1 = 4'd5; b_sign2 = 4'd13; b_sign3 = 4'd9;
@(posedge clk_i);
a_mant0 = 8'd44; a_mant1 = 8'd184; a_mant2 = 8'd158; a_mant3 = 8'd191;
b_mant0 = 8'd111; b_mant1 = 8'd44; b_mant2 = 8'd1; b_mant3 = 8'd96;
a_exp0 = 10'd151; a_exp1 = 10'd130; a_exp2 = 10'd204; a_exp3 = 10'd795;
b_exp0 = 10'd423; b_exp1 = 10'd305; b_exp2 = 10'd913; b_exp3 = 10'd876;
a_sign0 = 4'd14; a_sign1 = 4'd7; a_sign2 = 4'd8; a_sign3 = 4'd15;
b_sign0 = 4'd0; b_sign1 = 4'd13; b_sign2 = 4'd9; b_sign3 = 4'd9;
@(posedge clk_i);
shared_exps0 = 8'd134;
shared_exps1 = 8'd127;
a_mant0 = 8'd77; a_mant1 = 8'd192; a_mant2 = 8'd9; a_mant3 = 8'd184;
b_mant0 = 8'd146; b_mant1 = 8'd48; b_mant2 = 8'd178; b_mant3 = 8'd43;
a_exp0 = 10'd886; a_exp1 = 10'd834; a_exp2 = 10'd925; a_exp3 = 10'd323;
b_exp0 = 10'd686; b_exp1 = 10'd932; b_exp2 = 10'd585; b_exp3 = 10'd546;
a_sign0 = 4'd8; a_sign1 = 4'd15; a_sign2 = 4'd2; a_sign3 = 4'd10;
b_sign0 = 4'd14; b_sign1 = 4'd14; b_sign2 = 4'd6; b_sign3 = 4'd7;
@(posedge clk_i);
a_mant0 = 8'd71; a_mant1 = 8'd243; a_mant2 = 8'd170; a_mant3 = 8'd198;
b_mant0 = 8'd113; b_mant1 = 8'd5; b_mant2 = 8'd161; b_mant3 = 8'd186;
a_exp0 = 10'd991; a_exp1 = 10'd687; a_exp2 = 10'd326; a_exp3 = 10'd534;
b_exp0 = 10'd396; b_exp1 = 10'd431; b_exp2 = 10'd922; b_exp3 = 10'd499;
a_sign0 = 4'd11; a_sign1 = 4'd14; a_sign2 = 4'd14; a_sign3 = 4'd12;
b_sign0 = 4'd14; b_sign1 = 4'd12; b_sign2 = 4'd13; b_sign3 = 4'd4;
@(posedge clk_i);
a_mant0 = 8'd173; a_mant1 = 8'd21; a_mant2 = 8'd223; a_mant3 = 8'd254;
b_mant0 = 8'd4; b_mant1 = 8'd205; b_mant2 = 8'd12; b_mant3 = 8'd175;
a_exp0 = 10'd856; a_exp1 = 10'd317; a_exp2 = 10'd1014; a_exp3 = 10'd260;
b_exp0 = 10'd810; b_exp1 = 10'd788; b_exp2 = 10'd531; b_exp3 = 10'd54;
a_sign0 = 4'd8; a_sign1 = 4'd6; a_sign2 = 4'd16; a_sign3 = 4'd8;
b_sign0 = 4'd12; b_sign1 = 4'd7; b_sign2 = 4'd9; b_sign3 = 4'd3;
@(posedge clk_i);
a_mant0 = 8'd104; a_mant1 = 8'd202; a_mant2 = 8'd123; a_mant3 = 8'd119;
b_mant0 = 8'd24; b_mant1 = 8'd144; b_mant2 = 8'd138; b_mant3 = 8'd131;
a_exp0 = 10'd439; a_exp1 = 10'd421; a_exp2 = 10'd211; a_exp3 = 10'd126;
b_exp0 = 10'd893; b_exp1 = 10'd1009; b_exp2 = 10'd241; b_exp3 = 10'd986;
a_sign0 = 4'd9; a_sign1 = 4'd10; a_sign2 = 4'd12; a_sign3 = 4'd12;
b_sign0 = 4'd1; b_sign1 = 4'd12; b_sign2 = 4'd3; b_sign3 = 4'd6;
@(posedge clk_i);
a_mant0 = 8'd198; a_mant1 = 8'd154; a_mant2 = 8'd126; a_mant3 = 8'd215;
b_mant0 = 8'd44; b_mant1 = 8'd209; b_mant2 = 8'd158; b_mant3 = 8'd173;
a_exp0 = 10'd717; a_exp1 = 10'd610; a_exp2 = 10'd7; a_exp3 = 10'd413;
b_exp0 = 10'd342; b_exp1 = 10'd338; b_exp2 = 10'd646; b_exp3 = 10'd1001;
a_sign0 = 4'd6; a_sign1 = 4'd12; a_sign2 = 4'd14; a_sign3 = 4'd2;
b_sign0 = 4'd3; b_sign1 = 4'd1; b_sign2 = 4'd0; b_sign3 = 4'd12;
@(posedge clk_i);
a_mant0 = 8'd182; a_mant1 = 8'd4; a_mant2 = 8'd85; a_mant3 = 8'd86;
b_mant0 = 8'd31; b_mant1 = 8'd207; b_mant2 = 8'd208; b_mant3 = 8'd93;
a_exp0 = 10'd774; a_exp1 = 10'd470; a_exp2 = 10'd994; a_exp3 = 10'd114;
b_exp0 = 10'd894; b_exp1 = 10'd704; b_exp2 = 10'd890; b_exp3 = 10'd818;
a_sign0 = 4'd11; a_sign1 = 4'd2; a_sign2 = 4'd8; a_sign3 = 4'd6;
b_sign0 = 4'd3; b_sign1 = 4'd4; b_sign2 = 4'd11; b_sign3 = 4'd2;
@(posedge clk_i);
a_mant0 = 8'd36; a_mant1 = 8'd35; a_mant2 = 8'd229; a_mant3 = 8'd60;
b_mant0 = 8'd168; b_mant1 = 8'd104; b_mant2 = 8'd196; b_mant3 = 8'd144;
a_exp0 = 10'd733; a_exp1 = 10'd684; a_exp2 = 10'd199; a_exp3 = 10'd716;
b_exp0 = 10'd926; b_exp1 = 10'd157; b_exp2 = 10'd948; b_exp3 = 10'd844;
a_sign0 = 4'd8; a_sign1 = 4'd14; a_sign2 = 4'd2; a_sign3 = 4'd3;
b_sign0 = 4'd10; b_sign1 = 4'd1; b_sign2 = 4'd3; b_sign3 = 4'd5;
@(posedge clk_i);
a_mant0 = 8'd245; a_mant1 = 8'd28; a_mant2 = 8'd180; a_mant3 = 8'd198;
b_mant0 = 8'd46; b_mant1 = 8'd249; b_mant2 = 8'd230; b_mant3 = 8'd23;
a_exp0 = 10'd122; a_exp1 = 10'd202; a_exp2 = 10'd766; a_exp3 = 10'd563;
b_exp0 = 10'd659; b_exp1 = 10'd28; b_exp2 = 10'd424; b_exp3 = 10'd430;
a_sign0 = 4'd0; a_sign1 = 4'd11; a_sign2 = 4'd6; a_sign3 = 4'd7;
b_sign0 = 4'd1; b_sign1 = 4'd15; b_sign2 = 4'd0; b_sign3 = 4'd16;
@(posedge clk_i);
shared_exps0 = 8'd133;
shared_exps1 = 8'd141;
a_mant0 = 8'd141; a_mant1 = 8'd120; a_mant2 = 8'd79; a_mant3 = 8'd214;
b_mant0 = 8'd123; b_mant1 = 8'd178; b_mant2 = 8'd252; b_mant3 = 8'd231;
a_exp0 = 10'd87; a_exp1 = 10'd981; a_exp2 = 10'd931; a_exp3 = 10'd672;
b_exp0 = 10'd834; b_exp1 = 10'd595; b_exp2 = 10'd57; b_exp3 = 10'd470;
a_sign0 = 4'd6; a_sign1 = 4'd11; a_sign2 = 4'd14; a_sign3 = 4'd15;
b_sign0 = 4'd9; b_sign1 = 4'd1; b_sign2 = 4'd12; b_sign3 = 4'd15;
@(posedge clk_i);
a_mant0 = 8'd112; a_mant1 = 8'd87; a_mant2 = 8'd170; a_mant3 = 8'd99;
b_mant0 = 8'd146; b_mant1 = 8'd249; b_mant2 = 8'd53; b_mant3 = 8'd91;
a_exp0 = 10'd841; a_exp1 = 10'd365; a_exp2 = 10'd71; a_exp3 = 10'd113;
b_exp0 = 10'd646; b_exp1 = 10'd986; b_exp2 = 10'd255; b_exp3 = 10'd989;
a_sign0 = 4'd13; a_sign1 = 4'd14; a_sign2 = 4'd16; a_sign3 = 4'd2;
b_sign0 = 4'd10; b_sign1 = 4'd14; b_sign2 = 4'd0; b_sign3 = 4'd15;
@(posedge clk_i);
a_mant0 = 8'd79; a_mant1 = 8'd52; a_mant2 = 8'd69; a_mant3 = 8'd192;
b_mant0 = 8'd140; b_mant1 = 8'd242; b_mant2 = 8'd129; b_mant3 = 8'd5;
a_exp0 = 10'd273; a_exp1 = 10'd650; a_exp2 = 10'd356; a_exp3 = 10'd818;
b_exp0 = 10'd1003; b_exp1 = 10'd749; b_exp2 = 10'd39; b_exp3 = 10'd402;
a_sign0 = 4'd10; a_sign1 = 4'd14; a_sign2 = 4'd3; a_sign3 = 4'd7;
b_sign0 = 4'd16; b_sign1 = 4'd8; b_sign2 = 4'd7; b_sign3 = 4'd16;
@(posedge clk_i);
a_mant0 = 8'd220; a_mant1 = 8'd192; a_mant2 = 8'd87; a_mant3 = 8'd80;
b_mant0 = 8'd227; b_mant1 = 8'd197; b_mant2 = 8'd138; b_mant3 = 8'd35;
a_exp0 = 10'd21; a_exp1 = 10'd384; a_exp2 = 10'd20; a_exp3 = 10'd415;
b_exp0 = 10'd476; b_exp1 = 10'd923; b_exp2 = 10'd45; b_exp3 = 10'd369;
a_sign0 = 4'd14; a_sign1 = 4'd15; a_sign2 = 4'd7; a_sign3 = 4'd0;
b_sign0 = 4'd4; b_sign1 = 4'd2; b_sign2 = 4'd16; b_sign3 = 4'd4;
@(posedge clk_i);
a_mant0 = 8'd165; a_mant1 = 8'd202; a_mant2 = 8'd139; a_mant3 = 8'd234;
b_mant0 = 8'd37; b_mant1 = 8'd54; b_mant2 = 8'd129; b_mant3 = 8'd149;
a_exp0 = 10'd750; a_exp1 = 10'd499; a_exp2 = 10'd777; a_exp3 = 10'd30;
b_exp0 = 10'd817; b_exp1 = 10'd681; b_exp2 = 10'd264; b_exp3 = 10'd282;
a_sign0 = 4'd2; a_sign1 = 4'd3; a_sign2 = 4'd1; a_sign3 = 4'd10;
b_sign0 = 4'd3; b_sign1 = 4'd2; b_sign2 = 4'd13; b_sign3 = 4'd5;
@(posedge clk_i);
a_mant0 = 8'd118; a_mant1 = 8'd55; a_mant2 = 8'd19; a_mant3 = 8'd240;
b_mant0 = 8'd83; b_mant1 = 8'd171; b_mant2 = 8'd116; b_mant3 = 8'd213;
a_exp0 = 10'd243; a_exp1 = 10'd205; a_exp2 = 10'd589; a_exp3 = 10'd129;
b_exp0 = 10'd231; b_exp1 = 10'd856; b_exp2 = 10'd693; b_exp3 = 10'd1016;
a_sign0 = 4'd9; a_sign1 = 4'd8; a_sign2 = 4'd14; a_sign3 = 4'd6;
b_sign0 = 4'd14; b_sign1 = 4'd13; b_sign2 = 4'd6; b_sign3 = 4'd10;
@(posedge clk_i);
a_mant0 = 8'd70; a_mant1 = 8'd60; a_mant2 = 8'd99; a_mant3 = 8'd145;
b_mant0 = 8'd128; b_mant1 = 8'd104; b_mant2 = 8'd120; b_mant3 = 8'd207;
a_exp0 = 10'd958; a_exp1 = 10'd338; a_exp2 = 10'd289; a_exp3 = 10'd206;
b_exp0 = 10'd699; b_exp1 = 10'd856; b_exp2 = 10'd126; b_exp3 = 10'd7;
a_sign0 = 4'd11; a_sign1 = 4'd14; a_sign2 = 4'd4; a_sign3 = 4'd16;
b_sign0 = 4'd5; b_sign1 = 4'd4; b_sign2 = 4'd0; b_sign3 = 4'd8;
@(posedge clk_i);
a_mant0 = 8'd138; a_mant1 = 8'd7; a_mant2 = 8'd164; a_mant3 = 8'd28;
b_mant0 = 8'd86; b_mant1 = 8'd157; b_mant2 = 8'd234; b_mant3 = 8'd117;
a_exp0 = 10'd650; a_exp1 = 10'd846; a_exp2 = 10'd806; a_exp3 = 10'd852;
b_exp0 = 10'd687; b_exp1 = 10'd234; b_exp2 = 10'd941; b_exp3 = 10'd51;
a_sign0 = 4'd8; a_sign1 = 4'd8; a_sign2 = 4'd2; a_sign3 = 4'd8;
b_sign0 = 4'd8; b_sign1 = 4'd12; b_sign2 = 4'd12; b_sign3 = 4'd15;
@(posedge clk_i);
shared_exps0 = 8'd156;
shared_exps1 = 8'd134;
rstn = 0;
@(posedge clk_i);
rstn = 1;
a_mant0 = 8'd126; a_mant1 = 8'd197; a_mant2 = 8'd106; a_mant3 = 8'd147;
b_mant0 = 8'd122; b_mant1 = 8'd150; b_mant2 = 8'd67; b_mant3 = 8'd24;
a_exp0 = 10'd622; a_exp1 = 10'd823; a_exp2 = 10'd863; a_exp3 = 10'd154;
b_exp0 = 10'd70; b_exp1 = 10'd104; b_exp2 = 10'd917; b_exp3 = 10'd459;
a_sign0 = 4'd3; a_sign1 = 4'd7; a_sign2 = 4'd1; a_sign3 = 4'd3;
b_sign0 = 4'd4; b_sign1 = 4'd12; b_sign2 = 4'd10; b_sign3 = 4'd14;
@(posedge clk_i);
a_mant0 = 8'd185; a_mant1 = 8'd237; a_mant2 = 8'd229; a_mant3 = 8'd137;
b_mant0 = 8'd156; b_mant1 = 8'd188; b_mant2 = 8'd184; b_mant3 = 8'd53;
a_exp0 = 10'd697; a_exp1 = 10'd793; a_exp2 = 10'd1010; a_exp3 = 10'd887;
b_exp0 = 10'd325; b_exp1 = 10'd584; b_exp2 = 10'd905; b_exp3 = 10'd413;
a_sign0 = 4'd9; a_sign1 = 4'd0; a_sign2 = 4'd10; a_sign3 = 4'd1;
b_sign0 = 4'd6; b_sign1 = 4'd6; b_sign2 = 4'd10; b_sign3 = 4'd13;
@(posedge clk_i);
a_mant0 = 8'd23; a_mant1 = 8'd41; a_mant2 = 8'd120; a_mant3 = 8'd96;
b_mant0 = 8'd225; b_mant1 = 8'd40; b_mant2 = 8'd212; b_mant3 = 8'd249;
a_exp0 = 10'd681; a_exp1 = 10'd867; a_exp2 = 10'd159; a_exp3 = 10'd60;
b_exp0 = 10'd324; b_exp1 = 10'd882; b_exp2 = 10'd503; b_exp3 = 10'd990;
a_sign0 = 4'd9; a_sign1 = 4'd14; a_sign2 = 4'd2; a_sign3 = 4'd2;
b_sign0 = 4'd12; b_sign1 = 4'd11; b_sign2 = 4'd12; b_sign3 = 4'd7;
@(posedge clk_i);
a_mant0 = 8'd89; a_mant1 = 8'd13; a_mant2 = 8'd204; a_mant3 = 8'd34;
b_mant0 = 8'd6; b_mant1 = 8'd65; b_mant2 = 8'd217; b_mant3 = 8'd252;
a_exp0 = 10'd685; a_exp1 = 10'd201; a_exp2 = 10'd643; a_exp3 = 10'd723;
b_exp0 = 10'd894; b_exp1 = 10'd369; b_exp2 = 10'd93; b_exp3 = 10'd780;
a_sign0 = 4'd6; a_sign1 = 4'd15; a_sign2 = 4'd3; a_sign3 = 4'd14;
b_sign0 = 4'd6; b_sign1 = 4'd14; b_sign2 = 4'd10; b_sign3 = 4'd15;
@(posedge clk_i);
a_mant0 = 8'd130; a_mant1 = 8'd105; a_mant2 = 8'd61; a_mant3 = 8'd52;
b_mant0 = 8'd252; b_mant1 = 8'd23; b_mant2 = 8'd83; b_mant3 = 8'd189;
a_exp0 = 10'd700; a_exp1 = 10'd893; a_exp2 = 10'd523; a_exp3 = 10'd184;
b_exp0 = 10'd136; b_exp1 = 10'd100; b_exp2 = 10'd250; b_exp3 = 10'd202;
a_sign0 = 4'd5; a_sign1 = 4'd12; a_sign2 = 4'd0; a_sign3 = 4'd2;
b_sign0 = 4'd6; b_sign1 = 4'd8; b_sign2 = 4'd5; b_sign3 = 4'd3;
@(posedge clk_i);
a_mant0 = 8'd56; a_mant1 = 8'd237; a_mant2 = 8'd193; a_mant3 = 8'd66;
b_mant0 = 8'd34; b_mant1 = 8'd22; b_mant2 = 8'd201; b_mant3 = 8'd74;
a_exp0 = 10'd203; a_exp1 = 10'd168; a_exp2 = 10'd706; a_exp3 = 10'd619;
b_exp0 = 10'd375; b_exp1 = 10'd812; b_exp2 = 10'd568; b_exp3 = 10'd822;
a_sign0 = 4'd2; a_sign1 = 4'd11; a_sign2 = 4'd11; a_sign3 = 4'd8;
b_sign0 = 4'd15; b_sign1 = 4'd11; b_sign2 = 4'd2; b_sign3 = 4'd5;
@(posedge clk_i);
a_mant0 = 8'd244; a_mant1 = 8'd166; a_mant2 = 8'd26; a_mant3 = 8'd237;
b_mant0 = 8'd178; b_mant1 = 8'd97; b_mant2 = 8'd77; b_mant3 = 8'd84;
a_exp0 = 10'd587; a_exp1 = 10'd278; a_exp2 = 10'd11; a_exp3 = 10'd698;
b_exp0 = 10'd69; b_exp1 = 10'd502; b_exp2 = 10'd423; b_exp3 = 10'd317;
a_sign0 = 4'd2; a_sign1 = 4'd0; a_sign2 = 4'd10; a_sign3 = 4'd13;
b_sign0 = 4'd7; b_sign1 = 4'd3; b_sign2 = 4'd0; b_sign3 = 4'd1;
@(posedge clk_i);
shared_exps0 = 8'd133;
shared_exps1 = 8'd162;
a_mant0 = 8'd25; a_mant1 = 8'd211; a_mant2 = 8'd117; a_mant3 = 8'd3;
b_mant0 = 8'd93; b_mant1 = 8'd203; b_mant2 = 8'd78; b_mant3 = 8'd110;
a_exp0 = 10'd825; a_exp1 = 10'd359; a_exp2 = 10'd130; a_exp3 = 10'd857;
b_exp0 = 10'd87; b_exp1 = 10'd445; b_exp2 = 10'd152; b_exp3 = 10'd224;
a_sign0 = 4'd7; a_sign1 = 4'd2; a_sign2 = 4'd8; a_sign3 = 4'd15;
b_sign0 = 4'd3; b_sign1 = 4'd10; b_sign2 = 4'd1; b_sign3 = 4'd16;
@(posedge clk_i);
a_mant0 = 8'd34; a_mant1 = 8'd117; a_mant2 = 8'd28; a_mant3 = 8'd142;
b_mant0 = 8'd244; b_mant1 = 8'd7; b_mant2 = 8'd121; b_mant3 = 8'd193;
a_exp0 = 10'd815; a_exp1 = 10'd58; a_exp2 = 10'd717; a_exp3 = 10'd832;
b_exp0 = 10'd196; b_exp1 = 10'd954; b_exp2 = 10'd952; b_exp3 = 10'd194;
a_sign0 = 4'd3; a_sign1 = 4'd6; a_sign2 = 4'd14; a_sign3 = 4'd10;
b_sign0 = 4'd13; b_sign1 = 4'd11; b_sign2 = 4'd1; b_sign3 = 4'd10;
@(posedge clk_i);
a_mant0 = 8'd82; a_mant1 = 8'd64; a_mant2 = 8'd37; a_mant3 = 8'd25;
b_mant0 = 8'd26; b_mant1 = 8'd0; b_mant2 = 8'd178; b_mant3 = 8'd160;
a_exp0 = 10'd12; a_exp1 = 10'd347; a_exp2 = 10'd92; a_exp3 = 10'd330;
b_exp0 = 10'd725; b_exp1 = 10'd90; b_exp2 = 10'd314; b_exp3 = 10'd919;
a_sign0 = 4'd12; a_sign1 = 4'd7; a_sign2 = 4'd4; a_sign3 = 4'd9;
b_sign0 = 4'd2; b_sign1 = 4'd10; b_sign2 = 4'd4; b_sign3 = 4'd11;
@(posedge clk_i);
a_mant0 = 8'd155; a_mant1 = 8'd246; a_mant2 = 8'd227; a_mant3 = 8'd108;
b_mant0 = 8'd36; b_mant1 = 8'd210; b_mant2 = 8'd179; b_mant3 = 8'd210;
a_exp0 = 10'd121; a_exp1 = 10'd394; a_exp2 = 10'd267; a_exp3 = 10'd185;
b_exp0 = 10'd895; b_exp1 = 10'd456; b_exp2 = 10'd494; b_exp3 = 10'd961;
a_sign0 = 4'd9; a_sign1 = 4'd16; a_sign2 = 4'd10; a_sign3 = 4'd11;
b_sign0 = 4'd8; b_sign1 = 4'd10; b_sign2 = 4'd9; b_sign3 = 4'd11;
@(posedge clk_i);
a_mant0 = 8'd170; a_mant1 = 8'd186; a_mant2 = 8'd72; a_mant3 = 8'd116;
b_mant0 = 8'd12; b_mant1 = 8'd156; b_mant2 = 8'd181; b_mant3 = 8'd251;
a_exp0 = 10'd164; a_exp1 = 10'd608; a_exp2 = 10'd937; a_exp3 = 10'd861;
b_exp0 = 10'd496; b_exp1 = 10'd925; b_exp2 = 10'd90; b_exp3 = 10'd699;
a_sign0 = 4'd7; a_sign1 = 4'd12; a_sign2 = 4'd14; a_sign3 = 4'd14;
b_sign0 = 4'd14; b_sign1 = 4'd2; b_sign2 = 4'd7; b_sign3 = 4'd12;
@(posedge clk_i);
a_mant0 = 8'd50; a_mant1 = 8'd85; a_mant2 = 8'd243; a_mant3 = 8'd8;
b_mant0 = 8'd42; b_mant1 = 8'd169; b_mant2 = 8'd60; b_mant3 = 8'd239;
a_exp0 = 10'd537; a_exp1 = 10'd884; a_exp2 = 10'd400; a_exp3 = 10'd321;
b_exp0 = 10'd838; b_exp1 = 10'd726; b_exp2 = 10'd478; b_exp3 = 10'd859;
a_sign0 = 4'd9; a_sign1 = 4'd9; a_sign2 = 4'd2; a_sign3 = 4'd7;
b_sign0 = 4'd12; b_sign1 = 4'd8; b_sign2 = 4'd5; b_sign3 = 4'd2;
@(posedge clk_i);
a_mant0 = 8'd78; a_mant1 = 8'd30; a_mant2 = 8'd187; a_mant3 = 8'd31;
b_mant0 = 8'd164; b_mant1 = 8'd80; b_mant2 = 8'd195; b_mant3 = 8'd84;
a_exp0 = 10'd518; a_exp1 = 10'd404; a_exp2 = 10'd42; a_exp3 = 10'd500;
b_exp0 = 10'd551; b_exp1 = 10'd166; b_exp2 = 10'd375; b_exp3 = 10'd624;
a_sign0 = 4'd9; a_sign1 = 4'd5; a_sign2 = 4'd12; a_sign3 = 4'd8;
b_sign0 = 4'd10; b_sign1 = 4'd1; b_sign2 = 4'd12; b_sign3 = 4'd15;
@(posedge clk_i);
a_mant0 = 8'd60; a_mant1 = 8'd243; a_mant2 = 8'd193; a_mant3 = 8'd7;
b_mant0 = 8'd160; b_mant1 = 8'd172; b_mant2 = 8'd134; b_mant3 = 8'd206;
a_exp0 = 10'd526; a_exp1 = 10'd747; a_exp2 = 10'd312; a_exp3 = 10'd587;
b_exp0 = 10'd444; b_exp1 = 10'd1021; b_exp2 = 10'd323; b_exp3 = 10'd899;
a_sign0 = 4'd5; a_sign1 = 4'd5; a_sign2 = 4'd14; a_sign3 = 4'd11;
b_sign0 = 4'd16; b_sign1 = 4'd10; b_sign2 = 4'd1; b_sign3 = 4'd5;
@(posedge clk_i);
shared_exps0 = 8'd131;
shared_exps1 = 8'd135;
a_mant0 = 8'd191; a_mant1 = 8'd152; a_mant2 = 8'd16; a_mant3 = 8'd219;
b_mant0 = 8'd138; b_mant1 = 8'd91; b_mant2 = 8'd218; b_mant3 = 8'd104;
a_exp0 = 10'd993; a_exp1 = 10'd752; a_exp2 = 10'd99; a_exp3 = 10'd237;
b_exp0 = 10'd1015; b_exp1 = 10'd969; b_exp2 = 10'd233; b_exp3 = 10'd936;
a_sign0 = 4'd5; a_sign1 = 4'd3; a_sign2 = 4'd6; a_sign3 = 4'd11;
b_sign0 = 4'd1; b_sign1 = 4'd4; b_sign2 = 4'd14; b_sign3 = 4'd15;
@(posedge clk_i);
a_mant0 = 8'd143; a_mant1 = 8'd107; a_mant2 = 8'd216; a_mant3 = 8'd30;
b_mant0 = 8'd68; b_mant1 = 8'd25; b_mant2 = 8'd178; b_mant3 = 8'd153;
a_exp0 = 10'd851; a_exp1 = 10'd188; a_exp2 = 10'd685; a_exp3 = 10'd498;
b_exp0 = 10'd720; b_exp1 = 10'd604; b_exp2 = 10'd697; b_exp3 = 10'd593;
a_sign0 = 4'd3; a_sign1 = 4'd9; a_sign2 = 4'd2; a_sign3 = 4'd12;
b_sign0 = 4'd8; b_sign1 = 4'd8; b_sign2 = 4'd14; b_sign3 = 4'd11;
@(posedge clk_i);
a_mant0 = 8'd51; a_mant1 = 8'd44; a_mant2 = 8'd157; a_mant3 = 8'd11;
b_mant0 = 8'd114; b_mant1 = 8'd57; b_mant2 = 8'd191; b_mant3 = 8'd243;
a_exp0 = 10'd984; a_exp1 = 10'd262; a_exp2 = 10'd358; a_exp3 = 10'd639;
b_exp0 = 10'd170; b_exp1 = 10'd220; b_exp2 = 10'd244; b_exp3 = 10'd906;
a_sign0 = 4'd9; a_sign1 = 4'd0; a_sign2 = 4'd0; a_sign3 = 4'd6;
b_sign0 = 4'd10; b_sign1 = 4'd12; b_sign2 = 4'd12; b_sign3 = 4'd14;
@(posedge clk_i);
a_mant0 = 8'd129; a_mant1 = 8'd191; a_mant2 = 8'd119; a_mant3 = 8'd3;
b_mant0 = 8'd40; b_mant1 = 8'd252; b_mant2 = 8'd9; b_mant3 = 8'd24;
a_exp0 = 10'd406; a_exp1 = 10'd151; a_exp2 = 10'd146; a_exp3 = 10'd225;
b_exp0 = 10'd465; b_exp1 = 10'd1020; b_exp2 = 10'd532; b_exp3 = 10'd990;
a_sign0 = 4'd0; a_sign1 = 4'd9; a_sign2 = 4'd4; a_sign3 = 4'd10;
b_sign0 = 4'd13; b_sign1 = 4'd0; b_sign2 = 4'd15; b_sign3 = 4'd16;
@(posedge clk_i);
a_mant0 = 8'd237; a_mant1 = 8'd176; a_mant2 = 8'd155; a_mant3 = 8'd193;
b_mant0 = 8'd189; b_mant1 = 8'd29; b_mant2 = 8'd99; b_mant3 = 8'd188;
a_exp0 = 10'd726; a_exp1 = 10'd175; a_exp2 = 10'd577; a_exp3 = 10'd286;
b_exp0 = 10'd510; b_exp1 = 10'd225; b_exp2 = 10'd407; b_exp3 = 10'd125;
a_sign0 = 4'd16; a_sign1 = 4'd10; a_sign2 = 4'd15; a_sign3 = 4'd7;
b_sign0 = 4'd9; b_sign1 = 4'd6; b_sign2 = 4'd4; b_sign3 = 4'd7;
@(posedge clk_i);
a_mant0 = 8'd113; a_mant1 = 8'd107; a_mant2 = 8'd189; a_mant3 = 8'd17;
b_mant0 = 8'd8; b_mant1 = 8'd148; b_mant2 = 8'd119; b_mant3 = 8'd98;
a_exp0 = 10'd22; a_exp1 = 10'd178; a_exp2 = 10'd495; a_exp3 = 10'd623;
b_exp0 = 10'd791; b_exp1 = 10'd447; b_exp2 = 10'd692; b_exp3 = 10'd723;
a_sign0 = 4'd9; a_sign1 = 4'd0; a_sign2 = 4'd3; a_sign3 = 4'd12;
b_sign0 = 4'd16; b_sign1 = 4'd12; b_sign2 = 4'd14; b_sign3 = 4'd15;
@(posedge clk_i);
a_mant0 = 8'd103; a_mant1 = 8'd106; a_mant2 = 8'd253; a_mant3 = 8'd149;
b_mant0 = 8'd49; b_mant1 = 8'd177; b_mant2 = 8'd28; b_mant3 = 8'd158;
a_exp0 = 10'd164; a_exp1 = 10'd384; a_exp2 = 10'd483; a_exp3 = 10'd191;
b_exp0 = 10'd484; b_exp1 = 10'd843; b_exp2 = 10'd894; b_exp3 = 10'd396;
a_sign0 = 4'd15; a_sign1 = 4'd2; a_sign2 = 4'd13; a_sign3 = 4'd0;
b_sign0 = 4'd9; b_sign1 = 4'd11; b_sign2 = 4'd5; b_sign3 = 4'd12;
@(posedge clk_i);
a_mant0 = 8'd196; a_mant1 = 8'd224; a_mant2 = 8'd69; a_mant3 = 8'd219;
b_mant0 = 8'd129; b_mant1 = 8'd41; b_mant2 = 8'd59; b_mant3 = 8'd95;
a_exp0 = 10'd259; a_exp1 = 10'd963; a_exp2 = 10'd604; a_exp3 = 10'd869;
b_exp0 = 10'd6; b_exp1 = 10'd54; b_exp2 = 10'd553; b_exp3 = 10'd643;
a_sign0 = 4'd7; a_sign1 = 4'd12; a_sign2 = 4'd11; a_sign3 = 4'd6;
b_sign0 = 4'd8; b_sign1 = 4'd8; b_sign2 = 4'd4; b_sign3 = 4'd1;
@(posedge clk_i);
shared_exps0 = 8'd141;
shared_exps1 = 8'd135;
a_mant0 = 8'd82; a_mant1 = 8'd56; a_mant2 = 8'd47; a_mant3 = 8'd216;
b_mant0 = 8'd109; b_mant1 = 8'd3; b_mant2 = 8'd168; b_mant3 = 8'd29;
a_exp0 = 10'd16; a_exp1 = 10'd171; a_exp2 = 10'd682; a_exp3 = 10'd202;
b_exp0 = 10'd912; b_exp1 = 10'd445; b_exp2 = 10'd781; b_exp3 = 10'd986;
a_sign0 = 4'd8; a_sign1 = 4'd8; a_sign2 = 4'd6; a_sign3 = 4'd12;
b_sign0 = 4'd10; b_sign1 = 4'd14; b_sign2 = 4'd3; b_sign3 = 4'd2;
@(posedge clk_i);
a_mant0 = 8'd151; a_mant1 = 8'd91; a_mant2 = 8'd47; a_mant3 = 8'd189;
b_mant0 = 8'd66; b_mant1 = 8'd250; b_mant2 = 8'd111; b_mant3 = 8'd32;
a_exp0 = 10'd194; a_exp1 = 10'd276; a_exp2 = 10'd777; a_exp3 = 10'd254;
b_exp0 = 10'd351; b_exp1 = 10'd230; b_exp2 = 10'd504; b_exp3 = 10'd1022;
a_sign0 = 4'd12; a_sign1 = 4'd13; a_sign2 = 4'd5; a_sign3 = 4'd12;
b_sign0 = 4'd15; b_sign1 = 4'd9; b_sign2 = 4'd2; b_sign3 = 4'd12;
@(posedge clk_i);
a_mant0 = 8'd62; a_mant1 = 8'd50; a_mant2 = 8'd54; a_mant3 = 8'd43;
b_mant0 = 8'd135; b_mant1 = 8'd220; b_mant2 = 8'd72; b_mant3 = 8'd247;
a_exp0 = 10'd323; a_exp1 = 10'd214; a_exp2 = 10'd422; a_exp3 = 10'd793;
b_exp0 = 10'd583; b_exp1 = 10'd439; b_exp2 = 10'd928; b_exp3 = 10'd302;
a_sign0 = 4'd4; a_sign1 = 4'd16; a_sign2 = 4'd14; a_sign3 = 4'd16;
b_sign0 = 4'd7; b_sign1 = 4'd13; b_sign2 = 4'd7; b_sign3 = 4'd4;
@(posedge clk_i);
a_mant0 = 8'd204; a_mant1 = 8'd163; a_mant2 = 8'd60; a_mant3 = 8'd44;
b_mant0 = 8'd171; b_mant1 = 8'd94; b_mant2 = 8'd140; b_mant3 = 8'd162;
a_exp0 = 10'd338; a_exp1 = 10'd946; a_exp2 = 10'd379; a_exp3 = 10'd409;
b_exp0 = 10'd520; b_exp1 = 10'd371; b_exp2 = 10'd906; b_exp3 = 10'd14;
a_sign0 = 4'd13; a_sign1 = 4'd2; a_sign2 = 4'd10; a_sign3 = 4'd0;
b_sign0 = 4'd8; b_sign1 = 4'd13; b_sign2 = 4'd12; b_sign3 = 4'd2;
@(posedge clk_i);
a_mant0 = 8'd155; a_mant1 = 8'd111; a_mant2 = 8'd139; a_mant3 = 8'd31;
b_mant0 = 8'd138; b_mant1 = 8'd229; b_mant2 = 8'd228; b_mant3 = 8'd129;
a_exp0 = 10'd933; a_exp1 = 10'd615; a_exp2 = 10'd710; a_exp3 = 10'd176;
b_exp0 = 10'd535; b_exp1 = 10'd470; b_exp2 = 10'd286; b_exp3 = 10'd523;
a_sign0 = 4'd14; a_sign1 = 4'd1; a_sign2 = 4'd10; a_sign3 = 4'd3;
b_sign0 = 4'd10; b_sign1 = 4'd1; b_sign2 = 4'd5; b_sign3 = 4'd14;
@(posedge clk_i);
a_mant0 = 8'd111; a_mant1 = 8'd94; a_mant2 = 8'd10; a_mant3 = 8'd181;
b_mant0 = 8'd125; b_mant1 = 8'd37; b_mant2 = 8'd200; b_mant3 = 8'd137;
a_exp0 = 10'd679; a_exp1 = 10'd991; a_exp2 = 10'd41; a_exp3 = 10'd172;
b_exp0 = 10'd11; b_exp1 = 10'd32; b_exp2 = 10'd468; b_exp3 = 10'd411;
a_sign0 = 4'd2; a_sign1 = 4'd1; a_sign2 = 4'd8; a_sign3 = 4'd12;
b_sign0 = 4'd5; b_sign1 = 4'd13; b_sign2 = 4'd13; b_sign3 = 4'd9;
@(posedge clk_i);
a_mant0 = 8'd29; a_mant1 = 8'd29; a_mant2 = 8'd203; a_mant3 = 8'd106;
b_mant0 = 8'd36; b_mant1 = 8'd45; b_mant2 = 8'd104; b_mant3 = 8'd3;
a_exp0 = 10'd670; a_exp1 = 10'd609; a_exp2 = 10'd856; a_exp3 = 10'd75;
b_exp0 = 10'd587; b_exp1 = 10'd637; b_exp2 = 10'd606; b_exp3 = 10'd515;
a_sign0 = 4'd1; a_sign1 = 4'd10; a_sign2 = 4'd6; a_sign3 = 4'd16;
b_sign0 = 4'd5; b_sign1 = 4'd6; b_sign2 = 4'd6; b_sign3 = 4'd7;
@(posedge clk_i);
a_mant0 = 8'd250; a_mant1 = 8'd246; a_mant2 = 8'd134; a_mant3 = 8'd68;
b_mant0 = 8'd103; b_mant1 = 8'd161; b_mant2 = 8'd63; b_mant3 = 8'd42;
a_exp0 = 10'd221; a_exp1 = 10'd183; a_exp2 = 10'd66; a_exp3 = 10'd458;
b_exp0 = 10'd487; b_exp1 = 10'd790; b_exp2 = 10'd855; b_exp3 = 10'd583;
a_sign0 = 4'd16; a_sign1 = 4'd2; a_sign2 = 4'd14; a_sign3 = 4'd4;
b_sign0 = 4'd5; b_sign1 = 4'd13; b_sign2 = 4'd0; b_sign3 = 4'd7;
@(posedge clk_i);
shared_exps0 = 8'd118;
shared_exps1 = 8'd120;
rstn = 0;
@(posedge clk_i);
rstn = 1;
a_mant0 = 8'd8; a_mant1 = 8'd121; a_mant2 = 8'd140; a_mant3 = 8'd237;
b_mant0 = 8'd209; b_mant1 = 8'd173; b_mant2 = 8'd170; b_mant3 = 8'd81;
a_exp0 = 10'd415; a_exp1 = 10'd66; a_exp2 = 10'd562; a_exp3 = 10'd581;
b_exp0 = 10'd485; b_exp1 = 10'd858; b_exp2 = 10'd619; b_exp3 = 10'd621;
a_sign0 = 4'd2; a_sign1 = 4'd14; a_sign2 = 4'd8; a_sign3 = 4'd15;
b_sign0 = 4'd0; b_sign1 = 4'd8; b_sign2 = 4'd12; b_sign3 = 4'd12;
@(posedge clk_i);
a_mant0 = 8'd136; a_mant1 = 8'd157; a_mant2 = 8'd253; a_mant3 = 8'd229;
b_mant0 = 8'd224; b_mant1 = 8'd54; b_mant2 = 8'd193; b_mant3 = 8'd16;
a_exp0 = 10'd810; a_exp1 = 10'd789; a_exp2 = 10'd524; a_exp3 = 10'd125;
b_exp0 = 10'd612; b_exp1 = 10'd746; b_exp2 = 10'd150; b_exp3 = 10'd914;
a_sign0 = 4'd3; a_sign1 = 4'd11; a_sign2 = 4'd13; a_sign3 = 4'd4;
b_sign0 = 4'd7; b_sign1 = 4'd14; b_sign2 = 4'd16; b_sign3 = 4'd14;
@(posedge clk_i);
a_mant0 = 8'd142; a_mant1 = 8'd50; a_mant2 = 8'd237; a_mant3 = 8'd168;
b_mant0 = 8'd192; b_mant1 = 8'd27; b_mant2 = 8'd188; b_mant3 = 8'd102;
a_exp0 = 10'd397; a_exp1 = 10'd525; a_exp2 = 10'd823; a_exp3 = 10'd240;
b_exp0 = 10'd482; b_exp1 = 10'd325; b_exp2 = 10'd93; b_exp3 = 10'd630;
a_sign0 = 4'd2; a_sign1 = 4'd4; a_sign2 = 4'd10; a_sign3 = 4'd3;
b_sign0 = 4'd2; b_sign1 = 4'd2; b_sign2 = 4'd9; b_sign3 = 4'd9;
@(posedge clk_i);
a_mant0 = 8'd124; a_mant1 = 8'd84; a_mant2 = 8'd10; a_mant3 = 8'd137;
b_mant0 = 8'd36; b_mant1 = 8'd235; b_mant2 = 8'd59; b_mant3 = 8'd35;
a_exp0 = 10'd114; a_exp1 = 10'd703; a_exp2 = 10'd282; a_exp3 = 10'd908;
b_exp0 = 10'd220; b_exp1 = 10'd145; b_exp2 = 10'd739; b_exp3 = 10'd543;
a_sign0 = 4'd1; a_sign1 = 4'd3; a_sign2 = 4'd0; a_sign3 = 4'd3;
b_sign0 = 4'd14; b_sign1 = 4'd10; b_sign2 = 4'd16; b_sign3 = 4'd4;
@(posedge clk_i);
a_mant0 = 8'd177; a_mant1 = 8'd19; a_mant2 = 8'd1; a_mant3 = 8'd119;
b_mant0 = 8'd170; b_mant1 = 8'd120; b_mant2 = 8'd183; b_mant3 = 8'd253;
a_exp0 = 10'd519; a_exp1 = 10'd49; a_exp2 = 10'd311; a_exp3 = 10'd855;
b_exp0 = 10'd870; b_exp1 = 10'd159; b_exp2 = 10'd402; b_exp3 = 10'd844;
a_sign0 = 4'd8; a_sign1 = 4'd7; a_sign2 = 4'd3; a_sign3 = 4'd1;
b_sign0 = 4'd5; b_sign1 = 4'd4; b_sign2 = 4'd6; b_sign3 = 4'd9;
@(posedge clk_i);
a_mant0 = 8'd159; a_mant1 = 8'd207; a_mant2 = 8'd142; a_mant3 = 8'd55;
b_mant0 = 8'd208; b_mant1 = 8'd185; b_mant2 = 8'd143; b_mant3 = 8'd150;
a_exp0 = 10'd256; a_exp1 = 10'd142; a_exp2 = 10'd88; a_exp3 = 10'd515;
b_exp0 = 10'd616; b_exp1 = 10'd340; b_exp2 = 10'd41; b_exp3 = 10'd552;
a_sign0 = 4'd12; a_sign1 = 4'd13; a_sign2 = 4'd0; a_sign3 = 4'd5;
b_sign0 = 4'd4; b_sign1 = 4'd11; b_sign2 = 4'd12; b_sign3 = 4'd2;
@(posedge clk_i);
a_mant0 = 8'd115; a_mant1 = 8'd46; a_mant2 = 8'd137; a_mant3 = 8'd106;
b_mant0 = 8'd224; b_mant1 = 8'd255; b_mant2 = 8'd11; b_mant3 = 8'd7;
a_exp0 = 10'd879; a_exp1 = 10'd173; a_exp2 = 10'd391; a_exp3 = 10'd244;
b_exp0 = 10'd546; b_exp1 = 10'd154; b_exp2 = 10'd213; b_exp3 = 10'd637;
a_sign0 = 4'd9; a_sign1 = 4'd13; a_sign2 = 4'd11; a_sign3 = 4'd0;
b_sign0 = 4'd11; b_sign1 = 4'd14; b_sign2 = 4'd13; b_sign3 = 4'd8;
@(posedge clk_i);
shared_exps0 = 8'd135;
shared_exps1 = 8'd122;
a_mant0 = 8'd126; a_mant1 = 8'd186; a_mant2 = 8'd158; a_mant3 = 8'd254;
b_mant0 = 8'd199; b_mant1 = 8'd244; b_mant2 = 8'd78; b_mant3 = 8'd221;
a_exp0 = 10'd646; a_exp1 = 10'd901; a_exp2 = 10'd229; a_exp3 = 10'd599;
b_exp0 = 10'd138; b_exp1 = 10'd96; b_exp2 = 10'd30; b_exp3 = 10'd10;
a_sign0 = 4'd6; a_sign1 = 4'd0; a_sign2 = 4'd14; a_sign3 = 4'd0;
b_sign0 = 4'd11; b_sign1 = 4'd11; b_sign2 = 4'd7; b_sign3 = 4'd5;
@(posedge clk_i);
a_mant0 = 8'd163; a_mant1 = 8'd121; a_mant2 = 8'd241; a_mant3 = 8'd155;
b_mant0 = 8'd34; b_mant1 = 8'd189; b_mant2 = 8'd138; b_mant3 = 8'd20;
a_exp0 = 10'd656; a_exp1 = 10'd781; a_exp2 = 10'd489; a_exp3 = 10'd6;
b_exp0 = 10'd134; b_exp1 = 10'd144; b_exp2 = 10'd682; b_exp3 = 10'd307;
a_sign0 = 4'd11; a_sign1 = 4'd1; a_sign2 = 4'd11; a_sign3 = 4'd3;
b_sign0 = 4'd5; b_sign1 = 4'd1; b_sign2 = 4'd0; b_sign3 = 4'd5;
@(posedge clk_i);
a_mant0 = 8'd8; a_mant1 = 8'd100; a_mant2 = 8'd61; a_mant3 = 8'd34;
b_mant0 = 8'd253; b_mant1 = 8'd2; b_mant2 = 8'd8; b_mant3 = 8'd244;
a_exp0 = 10'd945; a_exp1 = 10'd248; a_exp2 = 10'd889; a_exp3 = 10'd173;
b_exp0 = 10'd785; b_exp1 = 10'd452; b_exp2 = 10'd628; b_exp3 = 10'd566;
a_sign0 = 4'd4; a_sign1 = 4'd12; a_sign2 = 4'd16; a_sign3 = 4'd13;
b_sign0 = 4'd14; b_sign1 = 4'd8; b_sign2 = 4'd0; b_sign3 = 4'd13;
@(posedge clk_i);
a_mant0 = 8'd240; a_mant1 = 8'd12; a_mant2 = 8'd231; a_mant3 = 8'd2;
b_mant0 = 8'd44; b_mant1 = 8'd115; b_mant2 = 8'd35; b_mant3 = 8'd224;
a_exp0 = 10'd276; a_exp1 = 10'd508; a_exp2 = 10'd868; a_exp3 = 10'd279;
b_exp0 = 10'd785; b_exp1 = 10'd849; b_exp2 = 10'd1; b_exp3 = 10'd1019;
a_sign0 = 4'd5; a_sign1 = 4'd9; a_sign2 = 4'd13; a_sign3 = 4'd9;
b_sign0 = 4'd8; b_sign1 = 4'd8; b_sign2 = 4'd11; b_sign3 = 4'd15;
@(posedge clk_i);
a_mant0 = 8'd194; a_mant1 = 8'd239; a_mant2 = 8'd182; a_mant3 = 8'd71;
b_mant0 = 8'd22; b_mant1 = 8'd28; b_mant2 = 8'd179; b_mant3 = 8'd77;
a_exp0 = 10'd307; a_exp1 = 10'd622; a_exp2 = 10'd521; a_exp3 = 10'd837;
b_exp0 = 10'd818; b_exp1 = 10'd153; b_exp2 = 10'd197; b_exp3 = 10'd605;
a_sign0 = 4'd15; a_sign1 = 4'd12; a_sign2 = 4'd0; a_sign3 = 4'd15;
b_sign0 = 4'd7; b_sign1 = 4'd12; b_sign2 = 4'd15; b_sign3 = 4'd0;
@(posedge clk_i);
a_mant0 = 8'd253; a_mant1 = 8'd246; a_mant2 = 8'd204; a_mant3 = 8'd215;
b_mant0 = 8'd102; b_mant1 = 8'd206; b_mant2 = 8'd212; b_mant3 = 8'd61;
a_exp0 = 10'd436; a_exp1 = 10'd918; a_exp2 = 10'd55; a_exp3 = 10'd365;
b_exp0 = 10'd1017; b_exp1 = 10'd138; b_exp2 = 10'd674; b_exp3 = 10'd785;
a_sign0 = 4'd2; a_sign1 = 4'd5; a_sign2 = 4'd4; a_sign3 = 4'd14;
b_sign0 = 4'd3; b_sign1 = 4'd8; b_sign2 = 4'd1; b_sign3 = 4'd13;
@(posedge clk_i);
a_mant0 = 8'd163; a_mant1 = 8'd116; a_mant2 = 8'd125; a_mant3 = 8'd203;
b_mant0 = 8'd240; b_mant1 = 8'd112; b_mant2 = 8'd204; b_mant3 = 8'd233;
a_exp0 = 10'd994; a_exp1 = 10'd173; a_exp2 = 10'd336; a_exp3 = 10'd1006;
b_exp0 = 10'd536; b_exp1 = 10'd924; b_exp2 = 10'd957; b_exp3 = 10'd583;
a_sign0 = 4'd7; a_sign1 = 4'd8; a_sign2 = 4'd11; a_sign3 = 4'd11;
b_sign0 = 4'd8; b_sign1 = 4'd2; b_sign2 = 4'd4; b_sign3 = 4'd13;
@(posedge clk_i);
a_mant0 = 8'd162; a_mant1 = 8'd101; a_mant2 = 8'd62; a_mant3 = 8'd237;
b_mant0 = 8'd228; b_mant1 = 8'd231; b_mant2 = 8'd145; b_mant3 = 8'd122;
a_exp0 = 10'd850; a_exp1 = 10'd263; a_exp2 = 10'd1000; a_exp3 = 10'd906;
b_exp0 = 10'd192; b_exp1 = 10'd470; b_exp2 = 10'd944; b_exp3 = 10'd774;
a_sign0 = 4'd13; a_sign1 = 4'd10; a_sign2 = 4'd3; a_sign3 = 4'd4;
b_sign0 = 4'd10; b_sign1 = 4'd3; b_sign2 = 4'd9; b_sign3 = 4'd10;
@(posedge clk_i);
shared_exps0 = 8'd152;
shared_exps1 = 8'd115;
a_mant0 = 8'd79; a_mant1 = 8'd106; a_mant2 = 8'd38; a_mant3 = 8'd232;
b_mant0 = 8'd81; b_mant1 = 8'd163; b_mant2 = 8'd109; b_mant3 = 8'd49;
a_exp0 = 10'd255; a_exp1 = 10'd368; a_exp2 = 10'd484; a_exp3 = 10'd118;
b_exp0 = 10'd358; b_exp1 = 10'd332; b_exp2 = 10'd802; b_exp3 = 10'd238;
a_sign0 = 4'd4; a_sign1 = 4'd0; a_sign2 = 4'd1; a_sign3 = 4'd4;
b_sign0 = 4'd4; b_sign1 = 4'd3; b_sign2 = 4'd0; b_sign3 = 4'd3;
@(posedge clk_i);
a_mant0 = 8'd78; a_mant1 = 8'd42; a_mant2 = 8'd95; a_mant3 = 8'd20;
b_mant0 = 8'd222; b_mant1 = 8'd235; b_mant2 = 8'd147; b_mant3 = 8'd241;
a_exp0 = 10'd1004; a_exp1 = 10'd664; a_exp2 = 10'd285; a_exp3 = 10'd289;
b_exp0 = 10'd282; b_exp1 = 10'd600; b_exp2 = 10'd928; b_exp3 = 10'd137;
a_sign0 = 4'd5; a_sign1 = 4'd16; a_sign2 = 4'd13; a_sign3 = 4'd10;
b_sign0 = 4'd10; b_sign1 = 4'd13; b_sign2 = 4'd15; b_sign3 = 4'd10;
@(posedge clk_i);
a_mant0 = 8'd166; a_mant1 = 8'd87; a_mant2 = 8'd243; a_mant3 = 8'd109;
b_mant0 = 8'd165; b_mant1 = 8'd113; b_mant2 = 8'd35; b_mant3 = 8'd179;
a_exp0 = 10'd821; a_exp1 = 10'd794; a_exp2 = 10'd367; a_exp3 = 10'd210;
b_exp0 = 10'd216; b_exp1 = 10'd120; b_exp2 = 10'd117; b_exp3 = 10'd516;
a_sign0 = 4'd12; a_sign1 = 4'd7; a_sign2 = 4'd4; a_sign3 = 4'd9;
b_sign0 = 4'd14; b_sign1 = 4'd0; b_sign2 = 4'd0; b_sign3 = 4'd16;
@(posedge clk_i);
a_mant0 = 8'd174; a_mant1 = 8'd199; a_mant2 = 8'd240; a_mant3 = 8'd4;
b_mant0 = 8'd174; b_mant1 = 8'd90; b_mant2 = 8'd215; b_mant3 = 8'd147;
a_exp0 = 10'd121; a_exp1 = 10'd261; a_exp2 = 10'd309; a_exp3 = 10'd850;
b_exp0 = 10'd21; b_exp1 = 10'd144; b_exp2 = 10'd313; b_exp3 = 10'd11;
a_sign0 = 4'd2; a_sign1 = 4'd16; a_sign2 = 4'd13; a_sign3 = 4'd2;
b_sign0 = 4'd13; b_sign1 = 4'd12; b_sign2 = 4'd11; b_sign3 = 4'd5;
@(posedge clk_i);
a_mant0 = 8'd50; a_mant1 = 8'd38; a_mant2 = 8'd200; a_mant3 = 8'd180;
b_mant0 = 8'd46; b_mant1 = 8'd65; b_mant2 = 8'd199; b_mant3 = 8'd115;
a_exp0 = 10'd379; a_exp1 = 10'd187; a_exp2 = 10'd716; a_exp3 = 10'd752;
b_exp0 = 10'd347; b_exp1 = 10'd171; b_exp2 = 10'd267; b_exp3 = 10'd538;
a_sign0 = 4'd5; a_sign1 = 4'd13; a_sign2 = 4'd9; a_sign3 = 4'd0;
b_sign0 = 4'd1; b_sign1 = 4'd16; b_sign2 = 4'd3; b_sign3 = 4'd2;
@(posedge clk_i);
a_mant0 = 8'd12; a_mant1 = 8'd65; a_mant2 = 8'd135; a_mant3 = 8'd161;
b_mant0 = 8'd6; b_mant1 = 8'd175; b_mant2 = 8'd98; b_mant3 = 8'd254;
a_exp0 = 10'd180; a_exp1 = 10'd620; a_exp2 = 10'd943; a_exp3 = 10'd940;
b_exp0 = 10'd185; b_exp1 = 10'd761; b_exp2 = 10'd1001; b_exp3 = 10'd831;
a_sign0 = 4'd1; a_sign1 = 4'd3; a_sign2 = 4'd4; a_sign3 = 4'd4;
b_sign0 = 4'd15; b_sign1 = 4'd13; b_sign2 = 4'd3; b_sign3 = 4'd15;
@(posedge clk_i);
a_mant0 = 8'd121; a_mant1 = 8'd80; a_mant2 = 8'd126; a_mant3 = 8'd176;
b_mant0 = 8'd145; b_mant1 = 8'd50; b_mant2 = 8'd105; b_mant3 = 8'd125;
a_exp0 = 10'd236; a_exp1 = 10'd728; a_exp2 = 10'd840; a_exp3 = 10'd40;
b_exp0 = 10'd892; b_exp1 = 10'd55; b_exp2 = 10'd236; b_exp3 = 10'd143;
a_sign0 = 4'd4; a_sign1 = 4'd10; a_sign2 = 4'd5; a_sign3 = 4'd10;
b_sign0 = 4'd8; b_sign1 = 4'd5; b_sign2 = 4'd14; b_sign3 = 4'd13;
@(posedge clk_i);
a_mant0 = 8'd73; a_mant1 = 8'd162; a_mant2 = 8'd236; a_mant3 = 8'd55;
b_mant0 = 8'd31; b_mant1 = 8'd128; b_mant2 = 8'd155; b_mant3 = 8'd15;
a_exp0 = 10'd564; a_exp1 = 10'd49; a_exp2 = 10'd333; a_exp3 = 10'd882;
b_exp0 = 10'd679; b_exp1 = 10'd773; b_exp2 = 10'd579; b_exp3 = 10'd365;
a_sign0 = 4'd4; a_sign1 = 4'd6; a_sign2 = 4'd4; a_sign3 = 4'd11;
b_sign0 = 4'd4; b_sign1 = 4'd9; b_sign2 = 4'd7; b_sign3 = 4'd3;
@(posedge clk_i);
shared_exps0 = 8'd143;
shared_exps1 = 8'd121;
a_mant0 = 8'd231; a_mant1 = 8'd192; a_mant2 = 8'd33; a_mant3 = 8'd183;
b_mant0 = 8'd147; b_mant1 = 8'd227; b_mant2 = 8'd30; b_mant3 = 8'd161;
a_exp0 = 10'd872; a_exp1 = 10'd75; a_exp2 = 10'd62; a_exp3 = 10'd423;
b_exp0 = 10'd859; b_exp1 = 10'd844; b_exp2 = 10'd200; b_exp3 = 10'd138;
a_sign0 = 4'd2; a_sign1 = 4'd14; a_sign2 = 4'd7; a_sign3 = 4'd8;
b_sign0 = 4'd7; b_sign1 = 4'd11; b_sign2 = 4'd6; b_sign3 = 4'd8;
@(posedge clk_i);
a_mant0 = 8'd12; a_mant1 = 8'd164; a_mant2 = 8'd164; a_mant3 = 8'd68;
b_mant0 = 8'd81; b_mant1 = 8'd155; b_mant2 = 8'd129; b_mant3 = 8'd203;
a_exp0 = 10'd531; a_exp1 = 10'd457; a_exp2 = 10'd227; a_exp3 = 10'd750;
b_exp0 = 10'd734; b_exp1 = 10'd308; b_exp2 = 10'd294; b_exp3 = 10'd332;
a_sign0 = 4'd8; a_sign1 = 4'd6; a_sign2 = 4'd12; a_sign3 = 4'd16;
b_sign0 = 4'd5; b_sign1 = 4'd2; b_sign2 = 4'd9; b_sign3 = 4'd6;
@(posedge clk_i);
a_mant0 = 8'd99; a_mant1 = 8'd104; a_mant2 = 8'd92; a_mant3 = 8'd186;
b_mant0 = 8'd126; b_mant1 = 8'd24; b_mant2 = 8'd96; b_mant3 = 8'd30;
a_exp0 = 10'd620; a_exp1 = 10'd408; a_exp2 = 10'd470; a_exp3 = 10'd479;
b_exp0 = 10'd1020; b_exp1 = 10'd97; b_exp2 = 10'd687; b_exp3 = 10'd218;
a_sign0 = 4'd1; a_sign1 = 4'd3; a_sign2 = 4'd4; a_sign3 = 4'd0;
b_sign0 = 4'd9; b_sign1 = 4'd6; b_sign2 = 4'd12; b_sign3 = 4'd16;
@(posedge clk_i);
a_mant0 = 8'd58; a_mant1 = 8'd173; a_mant2 = 8'd24; a_mant3 = 8'd232;
b_mant0 = 8'd247; b_mant1 = 8'd202; b_mant2 = 8'd107; b_mant3 = 8'd216;
a_exp0 = 10'd232; a_exp1 = 10'd433; a_exp2 = 10'd215; a_exp3 = 10'd379;
b_exp0 = 10'd659; b_exp1 = 10'd51; b_exp2 = 10'd587; b_exp3 = 10'd1007;
a_sign0 = 4'd3; a_sign1 = 4'd11; a_sign2 = 4'd11; a_sign3 = 4'd10;
b_sign0 = 4'd15; b_sign1 = 4'd14; b_sign2 = 4'd2; b_sign3 = 4'd16;
@(posedge clk_i);
a_mant0 = 8'd206; a_mant1 = 8'd9; a_mant2 = 8'd53; a_mant3 = 8'd9;
b_mant0 = 8'd74; b_mant1 = 8'd165; b_mant2 = 8'd58; b_mant3 = 8'd8;
a_exp0 = 10'd161; a_exp1 = 10'd141; a_exp2 = 10'd1021; a_exp3 = 10'd353;
b_exp0 = 10'd412; b_exp1 = 10'd981; b_exp2 = 10'd541; b_exp3 = 10'd254;
a_sign0 = 4'd13; a_sign1 = 4'd9; a_sign2 = 4'd16; a_sign3 = 4'd13;
b_sign0 = 4'd8; b_sign1 = 4'd6; b_sign2 = 4'd9; b_sign3 = 4'd10;
@(posedge clk_i);
a_mant0 = 8'd94; a_mant1 = 8'd154; a_mant2 = 8'd94; a_mant3 = 8'd152;
b_mant0 = 8'd29; b_mant1 = 8'd75; b_mant2 = 8'd16; b_mant3 = 8'd68;
a_exp0 = 10'd304; a_exp1 = 10'd844; a_exp2 = 10'd651; a_exp3 = 10'd879;
b_exp0 = 10'd972; b_exp1 = 10'd466; b_exp2 = 10'd47; b_exp3 = 10'd85;
a_sign0 = 4'd4; a_sign1 = 4'd0; a_sign2 = 4'd4; a_sign3 = 4'd6;
b_sign0 = 4'd9; b_sign1 = 4'd9; b_sign2 = 4'd13; b_sign3 = 4'd5;
@(posedge clk_i);
a_mant0 = 8'd215; a_mant1 = 8'd164; a_mant2 = 8'd12; a_mant3 = 8'd121;
b_mant0 = 8'd207; b_mant1 = 8'd51; b_mant2 = 8'd170; b_mant3 = 8'd97;
a_exp0 = 10'd471; a_exp1 = 10'd427; a_exp2 = 10'd246; a_exp3 = 10'd11;
b_exp0 = 10'd676; b_exp1 = 10'd110; b_exp2 = 10'd792; b_exp3 = 10'd400;
a_sign0 = 4'd9; a_sign1 = 4'd8; a_sign2 = 4'd12; a_sign3 = 4'd6;
b_sign0 = 4'd15; b_sign1 = 4'd12; b_sign2 = 4'd15; b_sign3 = 4'd15;
@(posedge clk_i);
a_mant0 = 8'd54; a_mant1 = 8'd88; a_mant2 = 8'd193; a_mant3 = 8'd215;
b_mant0 = 8'd47; b_mant1 = 8'd139; b_mant2 = 8'd195; b_mant3 = 8'd194;
a_exp0 = 10'd156; a_exp1 = 10'd364; a_exp2 = 10'd936; a_exp3 = 10'd559;
b_exp0 = 10'd503; b_exp1 = 10'd831; b_exp2 = 10'd664; b_exp3 = 10'd296;
a_sign0 = 4'd8; a_sign1 = 4'd11; a_sign2 = 4'd3; a_sign3 = 4'd7;
b_sign0 = 4'd6; b_sign1 = 4'd15; b_sign2 = 4'd11; b_sign3 = 4'd14;
@(posedge clk_i);
shared_exps0 = 8'd110;
shared_exps1 = 8'd100;
rstn = 0;
@(posedge clk_i);
rstn = 1;
a_mant0 = 8'd179; a_mant1 = 8'd89; a_mant2 = 8'd47; a_mant3 = 8'd180;
b_mant0 = 8'd29; b_mant1 = 8'd193; b_mant2 = 8'd192; b_mant3 = 8'd11;
a_exp0 = 10'd244; a_exp1 = 10'd72; a_exp2 = 10'd63; a_exp3 = 10'd120;
b_exp0 = 10'd887; b_exp1 = 10'd105; b_exp2 = 10'd499; b_exp3 = 10'd728;
a_sign0 = 4'd3; a_sign1 = 4'd15; a_sign2 = 4'd1; a_sign3 = 4'd6;
b_sign0 = 4'd8; b_sign1 = 4'd4; b_sign2 = 4'd1; b_sign3 = 4'd3;
@(posedge clk_i);
a_mant0 = 8'd68; a_mant1 = 8'd16; a_mant2 = 8'd168; a_mant3 = 8'd16;
b_mant0 = 8'd137; b_mant1 = 8'd237; b_mant2 = 8'd83; b_mant3 = 8'd87;
a_exp0 = 10'd530; a_exp1 = 10'd783; a_exp2 = 10'd954; a_exp3 = 10'd689;
b_exp0 = 10'd442; b_exp1 = 10'd875; b_exp2 = 10'd757; b_exp3 = 10'd944;
a_sign0 = 4'd6; a_sign1 = 4'd9; a_sign2 = 4'd5; a_sign3 = 4'd10;
b_sign0 = 4'd9; b_sign1 = 4'd2; b_sign2 = 4'd3; b_sign3 = 4'd3;
@(posedge clk_i);
a_mant0 = 8'd25; a_mant1 = 8'd174; a_mant2 = 8'd77; a_mant3 = 8'd226;
b_mant0 = 8'd133; b_mant1 = 8'd227; b_mant2 = 8'd61; b_mant3 = 8'd155;
a_exp0 = 10'd507; a_exp1 = 10'd522; a_exp2 = 10'd188; a_exp3 = 10'd344;
b_exp0 = 10'd418; b_exp1 = 10'd978; b_exp2 = 10'd274; b_exp3 = 10'd685;
a_sign0 = 4'd12; a_sign1 = 4'd4; a_sign2 = 4'd10; a_sign3 = 4'd13;
b_sign0 = 4'd5; b_sign1 = 4'd2; b_sign2 = 4'd0; b_sign3 = 4'd15;
@(posedge clk_i);
a_mant0 = 8'd155; a_mant1 = 8'd245; a_mant2 = 8'd220; a_mant3 = 8'd122;
b_mant0 = 8'd220; b_mant1 = 8'd71; b_mant2 = 8'd126; b_mant3 = 8'd162;
a_exp0 = 10'd871; a_exp1 = 10'd806; a_exp2 = 10'd47; a_exp3 = 10'd353;
b_exp0 = 10'd293; b_exp1 = 10'd742; b_exp2 = 10'd495; b_exp3 = 10'd124;
a_sign0 = 4'd2; a_sign1 = 4'd8; a_sign2 = 4'd11; a_sign3 = 4'd4;
b_sign0 = 4'd10; b_sign1 = 4'd12; b_sign2 = 4'd6; b_sign3 = 4'd15;
@(posedge clk_i);
a_mant0 = 8'd28; a_mant1 = 8'd32; a_mant2 = 8'd115; a_mant3 = 8'd92;
b_mant0 = 8'd235; b_mant1 = 8'd47; b_mant2 = 8'd107; b_mant3 = 8'd248;
a_exp0 = 10'd118; a_exp1 = 10'd398; a_exp2 = 10'd789; a_exp3 = 10'd811;
b_exp0 = 10'd723; b_exp1 = 10'd231; b_exp2 = 10'd709; b_exp3 = 10'd578;
a_sign0 = 4'd7; a_sign1 = 4'd12; a_sign2 = 4'd15; a_sign3 = 4'd16;
b_sign0 = 4'd4; b_sign1 = 4'd8; b_sign2 = 4'd3; b_sign3 = 4'd12;
@(posedge clk_i);
a_mant0 = 8'd73; a_mant1 = 8'd57; a_mant2 = 8'd12; a_mant3 = 8'd33;
b_mant0 = 8'd45; b_mant1 = 8'd6; b_mant2 = 8'd171; b_mant3 = 8'd248;
a_exp0 = 10'd781; a_exp1 = 10'd457; a_exp2 = 10'd738; a_exp3 = 10'd60;
b_exp0 = 10'd746; b_exp1 = 10'd251; b_exp2 = 10'd457; b_exp3 = 10'd39;
a_sign0 = 4'd4; a_sign1 = 4'd3; a_sign2 = 4'd9; a_sign3 = 4'd6;
b_sign0 = 4'd9; b_sign1 = 4'd7; b_sign2 = 4'd7; b_sign3 = 4'd3;
@(posedge clk_i);
a_mant0 = 8'd182; a_mant1 = 8'd171; a_mant2 = 8'd77; a_mant3 = 8'd65;
b_mant0 = 8'd56; b_mant1 = 8'd216; b_mant2 = 8'd236; b_mant3 = 8'd228;
a_exp0 = 10'd342; a_exp1 = 10'd667; a_exp2 = 10'd71; a_exp3 = 10'd267;
b_exp0 = 10'd646; b_exp1 = 10'd833; b_exp2 = 10'd661; b_exp3 = 10'd652;
a_sign0 = 4'd11; a_sign1 = 4'd13; a_sign2 = 4'd11; a_sign3 = 4'd10;
b_sign0 = 4'd2; b_sign1 = 4'd0; b_sign2 = 4'd6; b_sign3 = 4'd9;
@(posedge clk_i);
shared_exps0 = 8'd109;
shared_exps1 = 8'd136;
a_mant0 = 8'd16; a_mant1 = 8'd5; a_mant2 = 8'd0; a_mant3 = 8'd158;
b_mant0 = 8'd71; b_mant1 = 8'd17; b_mant2 = 8'd178; b_mant3 = 8'd149;
a_exp0 = 10'd573; a_exp1 = 10'd129; a_exp2 = 10'd910; a_exp3 = 10'd342;
b_exp0 = 10'd289; b_exp1 = 10'd733; b_exp2 = 10'd102; b_exp3 = 10'd258;
a_sign0 = 4'd4; a_sign1 = 4'd11; a_sign2 = 4'd8; a_sign3 = 4'd6;
b_sign0 = 4'd7; b_sign1 = 4'd2; b_sign2 = 4'd13; b_sign3 = 4'd10;
@(posedge clk_i);
a_mant0 = 8'd244; a_mant1 = 8'd199; a_mant2 = 8'd255; a_mant3 = 8'd227;
b_mant0 = 8'd155; b_mant1 = 8'd10; b_mant2 = 8'd153; b_mant3 = 8'd66;
a_exp0 = 10'd1000; a_exp1 = 10'd863; a_exp2 = 10'd423; a_exp3 = 10'd710;
b_exp0 = 10'd327; b_exp1 = 10'd498; b_exp2 = 10'd29; b_exp3 = 10'd329;
a_sign0 = 4'd4; a_sign1 = 4'd10; a_sign2 = 4'd0; a_sign3 = 4'd9;
b_sign0 = 4'd12; b_sign1 = 4'd14; b_sign2 = 4'd10; b_sign3 = 4'd13;
@(posedge clk_i);
a_mant0 = 8'd0; a_mant1 = 8'd74; a_mant2 = 8'd198; a_mant3 = 8'd244;
b_mant0 = 8'd112; b_mant1 = 8'd243; b_mant2 = 8'd7; b_mant3 = 8'd99;
a_exp0 = 10'd559; a_exp1 = 10'd786; a_exp2 = 10'd948; a_exp3 = 10'd171;
b_exp0 = 10'd541; b_exp1 = 10'd1021; b_exp2 = 10'd218; b_exp3 = 10'd581;
a_sign0 = 4'd0; a_sign1 = 4'd4; a_sign2 = 4'd9; a_sign3 = 4'd8;
b_sign0 = 4'd10; b_sign1 = 4'd8; b_sign2 = 4'd1; b_sign3 = 4'd5;
@(posedge clk_i);
a_mant0 = 8'd175; a_mant1 = 8'd198; a_mant2 = 8'd254; a_mant3 = 8'd169;
b_mant0 = 8'd124; b_mant1 = 8'd162; b_mant2 = 8'd38; b_mant3 = 8'd17;
a_exp0 = 10'd935; a_exp1 = 10'd728; a_exp2 = 10'd774; a_exp3 = 10'd764;
b_exp0 = 10'd398; b_exp1 = 10'd865; b_exp2 = 10'd491; b_exp3 = 10'd843;
a_sign0 = 4'd5; a_sign1 = 4'd12; a_sign2 = 4'd15; a_sign3 = 4'd14;
b_sign0 = 4'd7; b_sign1 = 4'd3; b_sign2 = 4'd7; b_sign3 = 4'd8;
@(posedge clk_i);
a_mant0 = 8'd4; a_mant1 = 8'd230; a_mant2 = 8'd204; a_mant3 = 8'd82;
b_mant0 = 8'd24; b_mant1 = 8'd73; b_mant2 = 8'd182; b_mant3 = 8'd65;
a_exp0 = 10'd2; a_exp1 = 10'd721; a_exp2 = 10'd752; a_exp3 = 10'd564;
b_exp0 = 10'd724; b_exp1 = 10'd586; b_exp2 = 10'd742; b_exp3 = 10'd78;
a_sign0 = 4'd16; a_sign1 = 4'd13; a_sign2 = 4'd10; a_sign3 = 4'd0;
b_sign0 = 4'd9; b_sign1 = 4'd1; b_sign2 = 4'd8; b_sign3 = 4'd2;
@(posedge clk_i);
a_mant0 = 8'd165; a_mant1 = 8'd10; a_mant2 = 8'd22; a_mant3 = 8'd113;
b_mant0 = 8'd140; b_mant1 = 8'd221; b_mant2 = 8'd214; b_mant3 = 8'd123;
a_exp0 = 10'd471; a_exp1 = 10'd820; a_exp2 = 10'd840; a_exp3 = 10'd648;
b_exp0 = 10'd109; b_exp1 = 10'd993; b_exp2 = 10'd548; b_exp3 = 10'd618;
a_sign0 = 4'd14; a_sign1 = 4'd15; a_sign2 = 4'd4; a_sign3 = 4'd3;
b_sign0 = 4'd10; b_sign1 = 4'd12; b_sign2 = 4'd11; b_sign3 = 4'd7;
@(posedge clk_i);
a_mant0 = 8'd69; a_mant1 = 8'd237; a_mant2 = 8'd75; a_mant3 = 8'd157;
b_mant0 = 8'd42; b_mant1 = 8'd183; b_mant2 = 8'd129; b_mant3 = 8'd58;
a_exp0 = 10'd431; a_exp1 = 10'd753; a_exp2 = 10'd166; a_exp3 = 10'd42;
b_exp0 = 10'd997; b_exp1 = 10'd727; b_exp2 = 10'd648; b_exp3 = 10'd238;
a_sign0 = 4'd15; a_sign1 = 4'd14; a_sign2 = 4'd6; a_sign3 = 4'd13;
b_sign0 = 4'd14; b_sign1 = 4'd2; b_sign2 = 4'd5; b_sign3 = 4'd10;
@(posedge clk_i);
a_mant0 = 8'd62; a_mant1 = 8'd107; a_mant2 = 8'd215; a_mant3 = 8'd105;
b_mant0 = 8'd222; b_mant1 = 8'd82; b_mant2 = 8'd251; b_mant3 = 8'd24;
a_exp0 = 10'd346; a_exp1 = 10'd547; a_exp2 = 10'd420; a_exp3 = 10'd741;
b_exp0 = 10'd725; b_exp1 = 10'd1014; b_exp2 = 10'd805; b_exp3 = 10'd623;
a_sign0 = 4'd16; a_sign1 = 4'd11; a_sign2 = 4'd6; a_sign3 = 4'd3;
b_sign0 = 4'd16; b_sign1 = 4'd5; b_sign2 = 4'd2; b_sign3 = 4'd14;
@(posedge clk_i);
shared_exps0 = 8'd119;
shared_exps1 = 8'd154;
a_mant0 = 8'd46; a_mant1 = 8'd224; a_mant2 = 8'd83; a_mant3 = 8'd236;
b_mant0 = 8'd155; b_mant1 = 8'd99; b_mant2 = 8'd83; b_mant3 = 8'd62;
a_exp0 = 10'd139; a_exp1 = 10'd630; a_exp2 = 10'd206; a_exp3 = 10'd730;
b_exp0 = 10'd349; b_exp1 = 10'd687; b_exp2 = 10'd421; b_exp3 = 10'd891;
a_sign0 = 4'd7; a_sign1 = 4'd12; a_sign2 = 4'd3; a_sign3 = 4'd7;
b_sign0 = 4'd15; b_sign1 = 4'd6; b_sign2 = 4'd14; b_sign3 = 4'd2;
@(posedge clk_i);
a_mant0 = 8'd133; a_mant1 = 8'd156; a_mant2 = 8'd98; a_mant3 = 8'd106;
b_mant0 = 8'd136; b_mant1 = 8'd56; b_mant2 = 8'd131; b_mant3 = 8'd16;
a_exp0 = 10'd283; a_exp1 = 10'd547; a_exp2 = 10'd904; a_exp3 = 10'd151;
b_exp0 = 10'd945; b_exp1 = 10'd468; b_exp2 = 10'd140; b_exp3 = 10'd400;
a_sign0 = 4'd14; a_sign1 = 4'd14; a_sign2 = 4'd0; a_sign3 = 4'd2;
b_sign0 = 4'd0; b_sign1 = 4'd14; b_sign2 = 4'd10; b_sign3 = 4'd2;
@(posedge clk_i);
a_mant0 = 8'd64; a_mant1 = 8'd115; a_mant2 = 8'd73; a_mant3 = 8'd29;
b_mant0 = 8'd64; b_mant1 = 8'd122; b_mant2 = 8'd43; b_mant3 = 8'd214;
a_exp0 = 10'd987; a_exp1 = 10'd313; a_exp2 = 10'd344; a_exp3 = 10'd142;
b_exp0 = 10'd818; b_exp1 = 10'd160; b_exp2 = 10'd549; b_exp3 = 10'd99;
a_sign0 = 4'd14; a_sign1 = 4'd2; a_sign2 = 4'd1; a_sign3 = 4'd14;
b_sign0 = 4'd12; b_sign1 = 4'd16; b_sign2 = 4'd9; b_sign3 = 4'd7;
@(posedge clk_i);
a_mant0 = 8'd110; a_mant1 = 8'd143; a_mant2 = 8'd43; a_mant3 = 8'd235;
b_mant0 = 8'd24; b_mant1 = 8'd217; b_mant2 = 8'd209; b_mant3 = 8'd113;
a_exp0 = 10'd227; a_exp1 = 10'd282; a_exp2 = 10'd810; a_exp3 = 10'd407;
b_exp0 = 10'd253; b_exp1 = 10'd330; b_exp2 = 10'd332; b_exp3 = 10'd306;
a_sign0 = 4'd15; a_sign1 = 4'd16; a_sign2 = 4'd5; a_sign3 = 4'd14;
b_sign0 = 4'd13; b_sign1 = 4'd12; b_sign2 = 4'd0; b_sign3 = 4'd6;
@(posedge clk_i);
a_mant0 = 8'd227; a_mant1 = 8'd236; a_mant2 = 8'd54; a_mant3 = 8'd237;
b_mant0 = 8'd9; b_mant1 = 8'd72; b_mant2 = 8'd27; b_mant3 = 8'd26;
a_exp0 = 10'd147; a_exp1 = 10'd809; a_exp2 = 10'd876; a_exp3 = 10'd501;
b_exp0 = 10'd187; b_exp1 = 10'd417; b_exp2 = 10'd426; b_exp3 = 10'd3;
a_sign0 = 4'd11; a_sign1 = 4'd5; a_sign2 = 4'd6; a_sign3 = 4'd15;
b_sign0 = 4'd13; b_sign1 = 4'd7; b_sign2 = 4'd5; b_sign3 = 4'd4;
@(posedge clk_i);
a_mant0 = 8'd140; a_mant1 = 8'd227; a_mant2 = 8'd42; a_mant3 = 8'd99;
b_mant0 = 8'd62; b_mant1 = 8'd21; b_mant2 = 8'd74; b_mant3 = 8'd66;
a_exp0 = 10'd747; a_exp1 = 10'd102; a_exp2 = 10'd282; a_exp3 = 10'd158;
b_exp0 = 10'd318; b_exp1 = 10'd569; b_exp2 = 10'd382; b_exp3 = 10'd582;
a_sign0 = 4'd13; a_sign1 = 4'd11; a_sign2 = 4'd13; a_sign3 = 4'd7;
b_sign0 = 4'd9; b_sign1 = 4'd7; b_sign2 = 4'd0; b_sign3 = 4'd15;
@(posedge clk_i);
a_mant0 = 8'd128; a_mant1 = 8'd53; a_mant2 = 8'd26; a_mant3 = 8'd81;
b_mant0 = 8'd83; b_mant1 = 8'd203; b_mant2 = 8'd12; b_mant3 = 8'd245;
a_exp0 = 10'd220; a_exp1 = 10'd720; a_exp2 = 10'd325; a_exp3 = 10'd554;
b_exp0 = 10'd99; b_exp1 = 10'd510; b_exp2 = 10'd922; b_exp3 = 10'd671;
a_sign0 = 4'd9; a_sign1 = 4'd6; a_sign2 = 4'd7; a_sign3 = 4'd13;
b_sign0 = 4'd12; b_sign1 = 4'd16; b_sign2 = 4'd5; b_sign3 = 4'd16;
@(posedge clk_i);
a_mant0 = 8'd110; a_mant1 = 8'd34; a_mant2 = 8'd236; a_mant3 = 8'd134;
b_mant0 = 8'd64; b_mant1 = 8'd109; b_mant2 = 8'd88; b_mant3 = 8'd221;
a_exp0 = 10'd655; a_exp1 = 10'd807; a_exp2 = 10'd795; a_exp3 = 10'd744;
b_exp0 = 10'd790; b_exp1 = 10'd998; b_exp2 = 10'd530; b_exp3 = 10'd268;
a_sign0 = 4'd8; a_sign1 = 4'd14; a_sign2 = 4'd5; a_sign3 = 4'd15;
b_sign0 = 4'd8; b_sign1 = 4'd9; b_sign2 = 4'd4; b_sign3 = 4'd2;
@(posedge clk_i);
shared_exps0 = 8'd122;
shared_exps1 = 8'd114;
a_mant0 = 8'd143; a_mant1 = 8'd76; a_mant2 = 8'd102; a_mant3 = 8'd37;
b_mant0 = 8'd31; b_mant1 = 8'd34; b_mant2 = 8'd7; b_mant3 = 8'd170;
a_exp0 = 10'd778; a_exp1 = 10'd133; a_exp2 = 10'd965; a_exp3 = 10'd914;
b_exp0 = 10'd445; b_exp1 = 10'd491; b_exp2 = 10'd761; b_exp3 = 10'd616;
a_sign0 = 4'd14; a_sign1 = 4'd0; a_sign2 = 4'd10; a_sign3 = 4'd0;
b_sign0 = 4'd5; b_sign1 = 4'd8; b_sign2 = 4'd15; b_sign3 = 4'd15;
@(posedge clk_i);
a_mant0 = 8'd189; a_mant1 = 8'd59; a_mant2 = 8'd249; a_mant3 = 8'd0;
b_mant0 = 8'd108; b_mant1 = 8'd44; b_mant2 = 8'd39; b_mant3 = 8'd203;
a_exp0 = 10'd430; a_exp1 = 10'd181; a_exp2 = 10'd725; a_exp3 = 10'd241;
b_exp0 = 10'd987; b_exp1 = 10'd394; b_exp2 = 10'd301; b_exp3 = 10'd295;
a_sign0 = 4'd6; a_sign1 = 4'd1; a_sign2 = 4'd13; a_sign3 = 4'd0;
b_sign0 = 4'd0; b_sign1 = 4'd13; b_sign2 = 4'd16; b_sign3 = 4'd8;
@(posedge clk_i);
a_mant0 = 8'd202; a_mant1 = 8'd185; a_mant2 = 8'd246; a_mant3 = 8'd29;
b_mant0 = 8'd22; b_mant1 = 8'd25; b_mant2 = 8'd28; b_mant3 = 8'd169;
a_exp0 = 10'd732; a_exp1 = 10'd669; a_exp2 = 10'd746; a_exp3 = 10'd629;
b_exp0 = 10'd21; b_exp1 = 10'd568; b_exp2 = 10'd953; b_exp3 = 10'd761;
a_sign0 = 4'd8; a_sign1 = 4'd16; a_sign2 = 4'd14; a_sign3 = 4'd14;
b_sign0 = 4'd14; b_sign1 = 4'd7; b_sign2 = 4'd12; b_sign3 = 4'd2;
@(posedge clk_i);
a_mant0 = 8'd102; a_mant1 = 8'd51; a_mant2 = 8'd55; a_mant3 = 8'd126;
b_mant0 = 8'd243; b_mant1 = 8'd190; b_mant2 = 8'd158; b_mant3 = 8'd89;
a_exp0 = 10'd135; a_exp1 = 10'd864; a_exp2 = 10'd747; a_exp3 = 10'd129;
b_exp0 = 10'd46; b_exp1 = 10'd756; b_exp2 = 10'd628; b_exp3 = 10'd766;
a_sign0 = 4'd8; a_sign1 = 4'd7; a_sign2 = 4'd10; a_sign3 = 4'd3;
b_sign0 = 4'd10; b_sign1 = 4'd2; b_sign2 = 4'd9; b_sign3 = 4'd13;
@(posedge clk_i);
a_mant0 = 8'd124; a_mant1 = 8'd135; a_mant2 = 8'd243; a_mant3 = 8'd55;
b_mant0 = 8'd130; b_mant1 = 8'd76; b_mant2 = 8'd168; b_mant3 = 8'd72;
a_exp0 = 10'd487; a_exp1 = 10'd567; a_exp2 = 10'd753; a_exp3 = 10'd504;
b_exp0 = 10'd69; b_exp1 = 10'd735; b_exp2 = 10'd299; b_exp3 = 10'd651;
a_sign0 = 4'd1; a_sign1 = 4'd8; a_sign2 = 4'd3; a_sign3 = 4'd6;
b_sign0 = 4'd1; b_sign1 = 4'd13; b_sign2 = 4'd2; b_sign3 = 4'd3;
@(posedge clk_i);
a_mant0 = 8'd206; a_mant1 = 8'd15; a_mant2 = 8'd92; a_mant3 = 8'd255;
b_mant0 = 8'd39; b_mant1 = 8'd168; b_mant2 = 8'd231; b_mant3 = 8'd189;
a_exp0 = 10'd169; a_exp1 = 10'd669; a_exp2 = 10'd350; a_exp3 = 10'd767;
b_exp0 = 10'd236; b_exp1 = 10'd1016; b_exp2 = 10'd757; b_exp3 = 10'd502;
a_sign0 = 4'd10; a_sign1 = 4'd9; a_sign2 = 4'd3; a_sign3 = 4'd11;
b_sign0 = 4'd3; b_sign1 = 4'd1; b_sign2 = 4'd16; b_sign3 = 4'd11;
@(posedge clk_i);
a_mant0 = 8'd218; a_mant1 = 8'd144; a_mant2 = 8'd96; a_mant3 = 8'd133;
b_mant0 = 8'd24; b_mant1 = 8'd94; b_mant2 = 8'd65; b_mant3 = 8'd200;
a_exp0 = 10'd259; a_exp1 = 10'd757; a_exp2 = 10'd637; a_exp3 = 10'd990;
b_exp0 = 10'd822; b_exp1 = 10'd261; b_exp2 = 10'd470; b_exp3 = 10'd916;
a_sign0 = 4'd8; a_sign1 = 4'd5; a_sign2 = 4'd2; a_sign3 = 4'd0;
b_sign0 = 4'd3; b_sign1 = 4'd3; b_sign2 = 4'd14; b_sign3 = 4'd14;
@(posedge clk_i);
a_mant0 = 8'd186; a_mant1 = 8'd37; a_mant2 = 8'd166; a_mant3 = 8'd174;
b_mant0 = 8'd74; b_mant1 = 8'd82; b_mant2 = 8'd175; b_mant3 = 8'd218;
a_exp0 = 10'd998; a_exp1 = 10'd148; a_exp2 = 10'd546; a_exp3 = 10'd22;
b_exp0 = 10'd171; b_exp1 = 10'd1017; b_exp2 = 10'd465; b_exp3 = 10'd837;
a_sign0 = 4'd9; a_sign1 = 4'd13; a_sign2 = 4'd5; a_sign3 = 4'd8;
b_sign0 = 4'd16; b_sign1 = 4'd5; b_sign2 = 4'd1; b_sign3 = 4'd11;
@(posedge clk_i);
shared_exps0 = 8'd121;
shared_exps1 = 8'd106;
rstn = 0;
@(posedge clk_i);
rstn = 1;
a_mant0 = 8'd192; a_mant1 = 8'd163; a_mant2 = 8'd90; a_mant3 = 8'd238;
b_mant0 = 8'd250; b_mant1 = 8'd171; b_mant2 = 8'd132; b_mant3 = 8'd26;
a_exp0 = 10'd987; a_exp1 = 10'd505; a_exp2 = 10'd702; a_exp3 = 10'd270;
b_exp0 = 10'd324; b_exp1 = 10'd938; b_exp2 = 10'd971; b_exp3 = 10'd330;
a_sign0 = 4'd7; a_sign1 = 4'd15; a_sign2 = 4'd9; a_sign3 = 4'd4;
b_sign0 = 4'd1; b_sign1 = 4'd13; b_sign2 = 4'd12; b_sign3 = 4'd7;
@(posedge clk_i);
a_mant0 = 8'd57; a_mant1 = 8'd92; a_mant2 = 8'd55; a_mant3 = 8'd201;
b_mant0 = 8'd34; b_mant1 = 8'd236; b_mant2 = 8'd91; b_mant3 = 8'd1;
a_exp0 = 10'd475; a_exp1 = 10'd953; a_exp2 = 10'd865; a_exp3 = 10'd562;
b_exp0 = 10'd301; b_exp1 = 10'd251; b_exp2 = 10'd401; b_exp3 = 10'd74;
a_sign0 = 4'd8; a_sign1 = 4'd9; a_sign2 = 4'd16; a_sign3 = 4'd0;
b_sign0 = 4'd10; b_sign1 = 4'd7; b_sign2 = 4'd4; b_sign3 = 4'd11;
@(posedge clk_i);
a_mant0 = 8'd167; a_mant1 = 8'd165; a_mant2 = 8'd110; a_mant3 = 8'd123;
b_mant0 = 8'd187; b_mant1 = 8'd207; b_mant2 = 8'd78; b_mant3 = 8'd51;
a_exp0 = 10'd81; a_exp1 = 10'd978; a_exp2 = 10'd925; a_exp3 = 10'd185;
b_exp0 = 10'd1003; b_exp1 = 10'd204; b_exp2 = 10'd338; b_exp3 = 10'd205;
a_sign0 = 4'd5; a_sign1 = 4'd7; a_sign2 = 4'd14; a_sign3 = 4'd15;
b_sign0 = 4'd10; b_sign1 = 4'd15; b_sign2 = 4'd11; b_sign3 = 4'd0;
@(posedge clk_i);
a_mant0 = 8'd178; a_mant1 = 8'd228; a_mant2 = 8'd4; a_mant3 = 8'd57;
b_mant0 = 8'd156; b_mant1 = 8'd78; b_mant2 = 8'd13; b_mant3 = 8'd1;
a_exp0 = 10'd302; a_exp1 = 10'd780; a_exp2 = 10'd795; a_exp3 = 10'd14;
b_exp0 = 10'd930; b_exp1 = 10'd173; b_exp2 = 10'd657; b_exp3 = 10'd1018;
a_sign0 = 4'd8; a_sign1 = 4'd5; a_sign2 = 4'd2; a_sign3 = 4'd16;
b_sign0 = 4'd15; b_sign1 = 4'd2; b_sign2 = 4'd13; b_sign3 = 4'd14;
@(posedge clk_i);
a_mant0 = 8'd29; a_mant1 = 8'd148; a_mant2 = 8'd232; a_mant3 = 8'd96;
b_mant0 = 8'd53; b_mant1 = 8'd189; b_mant2 = 8'd10; b_mant3 = 8'd189;
a_exp0 = 10'd82; a_exp1 = 10'd952; a_exp2 = 10'd770; a_exp3 = 10'd66;
b_exp0 = 10'd753; b_exp1 = 10'd918; b_exp2 = 10'd662; b_exp3 = 10'd454;
a_sign0 = 4'd7; a_sign1 = 4'd16; a_sign2 = 4'd14; a_sign3 = 4'd12;
b_sign0 = 4'd2; b_sign1 = 4'd2; b_sign2 = 4'd2; b_sign3 = 4'd11;
@(posedge clk_i);
a_mant0 = 8'd45; a_mant1 = 8'd41; a_mant2 = 8'd95; a_mant3 = 8'd90;
b_mant0 = 8'd147; b_mant1 = 8'd121; b_mant2 = 8'd156; b_mant3 = 8'd31;
a_exp0 = 10'd63; a_exp1 = 10'd828; a_exp2 = 10'd861; a_exp3 = 10'd154;
b_exp0 = 10'd865; b_exp1 = 10'd424; b_exp2 = 10'd468; b_exp3 = 10'd655;
a_sign0 = 4'd5; a_sign1 = 4'd5; a_sign2 = 4'd0; a_sign3 = 4'd10;
b_sign0 = 4'd13; b_sign1 = 4'd2; b_sign2 = 4'd0; b_sign3 = 4'd13;
@(posedge clk_i);
a_mant0 = 8'd205; a_mant1 = 8'd40; a_mant2 = 8'd126; a_mant3 = 8'd141;
b_mant0 = 8'd247; b_mant1 = 8'd231; b_mant2 = 8'd72; b_mant3 = 8'd13;
a_exp0 = 10'd514; a_exp1 = 10'd665; a_exp2 = 10'd236; a_exp3 = 10'd961;
b_exp0 = 10'd247; b_exp1 = 10'd194; b_exp2 = 10'd831; b_exp3 = 10'd328;
a_sign0 = 4'd1; a_sign1 = 4'd5; a_sign2 = 4'd5; a_sign3 = 4'd9;
b_sign0 = 4'd10; b_sign1 = 4'd13; b_sign2 = 4'd13; b_sign3 = 4'd7;
@(posedge clk_i);
shared_exps0 = 8'd127;
shared_exps1 = 8'd148;
a_mant0 = 8'd78; a_mant1 = 8'd77; a_mant2 = 8'd46; a_mant3 = 8'd179;
b_mant0 = 8'd205; b_mant1 = 8'd104; b_mant2 = 8'd187; b_mant3 = 8'd183;
a_exp0 = 10'd952; a_exp1 = 10'd752; a_exp2 = 10'd203; a_exp3 = 10'd254;
b_exp0 = 10'd996; b_exp1 = 10'd491; b_exp2 = 10'd855; b_exp3 = 10'd23;
a_sign0 = 4'd11; a_sign1 = 4'd3; a_sign2 = 4'd8; a_sign3 = 4'd1;
b_sign0 = 4'd9; b_sign1 = 4'd11; b_sign2 = 4'd0; b_sign3 = 4'd6;
@(posedge clk_i);
a_mant0 = 8'd203; a_mant1 = 8'd75; a_mant2 = 8'd202; a_mant3 = 8'd13;
b_mant0 = 8'd198; b_mant1 = 8'd89; b_mant2 = 8'd169; b_mant3 = 8'd165;
a_exp0 = 10'd929; a_exp1 = 10'd1006; a_exp2 = 10'd511; a_exp3 = 10'd723;
b_exp0 = 10'd134; b_exp1 = 10'd229; b_exp2 = 10'd341; b_exp3 = 10'd465;
a_sign0 = 4'd7; a_sign1 = 4'd15; a_sign2 = 4'd15; a_sign3 = 4'd8;
b_sign0 = 4'd8; b_sign1 = 4'd3; b_sign2 = 4'd12; b_sign3 = 4'd1;
@(posedge clk_i);
a_mant0 = 8'd231; a_mant1 = 8'd122; a_mant2 = 8'd220; a_mant3 = 8'd170;
b_mant0 = 8'd45; b_mant1 = 8'd165; b_mant2 = 8'd117; b_mant3 = 8'd138;
a_exp0 = 10'd172; a_exp1 = 10'd800; a_exp2 = 10'd286; a_exp3 = 10'd592;
b_exp0 = 10'd825; b_exp1 = 10'd768; b_exp2 = 10'd968; b_exp3 = 10'd626;
a_sign0 = 4'd13; a_sign1 = 4'd14; a_sign2 = 4'd8; a_sign3 = 4'd4;
b_sign0 = 4'd11; b_sign1 = 4'd16; b_sign2 = 4'd14; b_sign3 = 4'd12;
@(posedge clk_i);
a_mant0 = 8'd232; a_mant1 = 8'd201; a_mant2 = 8'd209; a_mant3 = 8'd203;
b_mant0 = 8'd33; b_mant1 = 8'd139; b_mant2 = 8'd253; b_mant3 = 8'd14;
a_exp0 = 10'd280; a_exp1 = 10'd485; a_exp2 = 10'd950; a_exp3 = 10'd205;
b_exp0 = 10'd665; b_exp1 = 10'd746; b_exp2 = 10'd320; b_exp3 = 10'd668;
a_sign0 = 4'd5; a_sign1 = 4'd8; a_sign2 = 4'd6; a_sign3 = 4'd12;
b_sign0 = 4'd8; b_sign1 = 4'd0; b_sign2 = 4'd0; b_sign3 = 4'd8;
@(posedge clk_i);
a_mant0 = 8'd71; a_mant1 = 8'd214; a_mant2 = 8'd223; a_mant3 = 8'd142;
b_mant0 = 8'd175; b_mant1 = 8'd75; b_mant2 = 8'd66; b_mant3 = 8'd25;
a_exp0 = 10'd28; a_exp1 = 10'd548; a_exp2 = 10'd811; a_exp3 = 10'd1000;
b_exp0 = 10'd855; b_exp1 = 10'd630; b_exp2 = 10'd968; b_exp3 = 10'd332;
a_sign0 = 4'd11; a_sign1 = 4'd8; a_sign2 = 4'd4; a_sign3 = 4'd7;
b_sign0 = 4'd4; b_sign1 = 4'd6; b_sign2 = 4'd11; b_sign3 = 4'd10;
@(posedge clk_i);
a_mant0 = 8'd9; a_mant1 = 8'd176; a_mant2 = 8'd103; a_mant3 = 8'd30;
b_mant0 = 8'd199; b_mant1 = 8'd225; b_mant2 = 8'd202; b_mant3 = 8'd105;
a_exp0 = 10'd751; a_exp1 = 10'd1013; a_exp2 = 10'd7; a_exp3 = 10'd332;
b_exp0 = 10'd730; b_exp1 = 10'd126; b_exp2 = 10'd575; b_exp3 = 10'd887;
a_sign0 = 4'd16; a_sign1 = 4'd11; a_sign2 = 4'd11; a_sign3 = 4'd6;
b_sign0 = 4'd2; b_sign1 = 4'd15; b_sign2 = 4'd8; b_sign3 = 4'd16;
@(posedge clk_i);
a_mant0 = 8'd185; a_mant1 = 8'd38; a_mant2 = 8'd129; a_mant3 = 8'd96;
b_mant0 = 8'd62; b_mant1 = 8'd149; b_mant2 = 8'd141; b_mant3 = 8'd212;
a_exp0 = 10'd49; a_exp1 = 10'd58; a_exp2 = 10'd593; a_exp3 = 10'd320;
b_exp0 = 10'd79; b_exp1 = 10'd832; b_exp2 = 10'd73; b_exp3 = 10'd14;
a_sign0 = 4'd12; a_sign1 = 4'd6; a_sign2 = 4'd0; a_sign3 = 4'd4;
b_sign0 = 4'd9; b_sign1 = 4'd0; b_sign2 = 4'd10; b_sign3 = 4'd3;
@(posedge clk_i);
a_mant0 = 8'd108; a_mant1 = 8'd131; a_mant2 = 8'd80; a_mant3 = 8'd60;
b_mant0 = 8'd82; b_mant1 = 8'd191; b_mant2 = 8'd141; b_mant3 = 8'd34;
a_exp0 = 10'd118; a_exp1 = 10'd715; a_exp2 = 10'd19; a_exp3 = 10'd101;
b_exp0 = 10'd141; b_exp1 = 10'd688; b_exp2 = 10'd664; b_exp3 = 10'd959;
a_sign0 = 4'd7; a_sign1 = 4'd13; a_sign2 = 4'd5; a_sign3 = 4'd14;
b_sign0 = 4'd1; b_sign1 = 4'd7; b_sign2 = 4'd1; b_sign3 = 4'd13;
@(posedge clk_i);
shared_exps0 = 8'd118;
shared_exps1 = 8'd146;
a_mant0 = 8'd154; a_mant1 = 8'd172; a_mant2 = 8'd157; a_mant3 = 8'd221;
b_mant0 = 8'd68; b_mant1 = 8'd100; b_mant2 = 8'd154; b_mant3 = 8'd61;
a_exp0 = 10'd616; a_exp1 = 10'd149; a_exp2 = 10'd775; a_exp3 = 10'd178;
b_exp0 = 10'd545; b_exp1 = 10'd151; b_exp2 = 10'd607; b_exp3 = 10'd823;
a_sign0 = 4'd0; a_sign1 = 4'd4; a_sign2 = 4'd10; a_sign3 = 4'd16;
b_sign0 = 4'd0; b_sign1 = 4'd11; b_sign2 = 4'd11; b_sign3 = 4'd4;
@(posedge clk_i);
a_mant0 = 8'd36; a_mant1 = 8'd40; a_mant2 = 8'd239; a_mant3 = 8'd87;
b_mant0 = 8'd41; b_mant1 = 8'd44; b_mant2 = 8'd223; b_mant3 = 8'd177;
a_exp0 = 10'd412; a_exp1 = 10'd584; a_exp2 = 10'd758; a_exp3 = 10'd252;
b_exp0 = 10'd914; b_exp1 = 10'd605; b_exp2 = 10'd154; b_exp3 = 10'd895;
a_sign0 = 4'd15; a_sign1 = 4'd8; a_sign2 = 4'd4; a_sign3 = 4'd8;
b_sign0 = 4'd9; b_sign1 = 4'd16; b_sign2 = 4'd8; b_sign3 = 4'd16;
@(posedge clk_i);
a_mant0 = 8'd250; a_mant1 = 8'd171; a_mant2 = 8'd88; a_mant3 = 8'd214;
b_mant0 = 8'd37; b_mant1 = 8'd238; b_mant2 = 8'd146; b_mant3 = 8'd135;
a_exp0 = 10'd172; a_exp1 = 10'd232; a_exp2 = 10'd201; a_exp3 = 10'd93;
b_exp0 = 10'd133; b_exp1 = 10'd181; b_exp2 = 10'd268; b_exp3 = 10'd993;
a_sign0 = 4'd0; a_sign1 = 4'd3; a_sign2 = 4'd13; a_sign3 = 4'd4;
b_sign0 = 4'd10; b_sign1 = 4'd5; b_sign2 = 4'd2; b_sign3 = 4'd9;
@(posedge clk_i);
a_mant0 = 8'd52; a_mant1 = 8'd125; a_mant2 = 8'd222; a_mant3 = 8'd105;
b_mant0 = 8'd82; b_mant1 = 8'd171; b_mant2 = 8'd24; b_mant3 = 8'd227;
a_exp0 = 10'd644; a_exp1 = 10'd949; a_exp2 = 10'd882; a_exp3 = 10'd513;
b_exp0 = 10'd935; b_exp1 = 10'd254; b_exp2 = 10'd642; b_exp3 = 10'd106;
a_sign0 = 4'd8; a_sign1 = 4'd2; a_sign2 = 4'd8; a_sign3 = 4'd5;
b_sign0 = 4'd7; b_sign1 = 4'd0; b_sign2 = 4'd14; b_sign3 = 4'd7;
@(posedge clk_i);
a_mant0 = 8'd34; a_mant1 = 8'd44; a_mant2 = 8'd210; a_mant3 = 8'd226;
b_mant0 = 8'd18; b_mant1 = 8'd219; b_mant2 = 8'd66; b_mant3 = 8'd166;
a_exp0 = 10'd908; a_exp1 = 10'd71; a_exp2 = 10'd755; a_exp3 = 10'd20;
b_exp0 = 10'd686; b_exp1 = 10'd913; b_exp2 = 10'd332; b_exp3 = 10'd46;
a_sign0 = 4'd16; a_sign1 = 4'd14; a_sign2 = 4'd13; a_sign3 = 4'd0;
b_sign0 = 4'd5; b_sign1 = 4'd3; b_sign2 = 4'd13; b_sign3 = 4'd2;
@(posedge clk_i);
a_mant0 = 8'd46; a_mant1 = 8'd134; a_mant2 = 8'd165; a_mant3 = 8'd79;
b_mant0 = 8'd103; b_mant1 = 8'd60; b_mant2 = 8'd249; b_mant3 = 8'd26;
a_exp0 = 10'd688; a_exp1 = 10'd595; a_exp2 = 10'd910; a_exp3 = 10'd696;
b_exp0 = 10'd908; b_exp1 = 10'd125; b_exp2 = 10'd251; b_exp3 = 10'd761;
a_sign0 = 4'd9; a_sign1 = 4'd11; a_sign2 = 4'd6; a_sign3 = 4'd11;
b_sign0 = 4'd5; b_sign1 = 4'd5; b_sign2 = 4'd0; b_sign3 = 4'd2;
@(posedge clk_i);
a_mant0 = 8'd11; a_mant1 = 8'd193; a_mant2 = 8'd125; a_mant3 = 8'd164;
b_mant0 = 8'd19; b_mant1 = 8'd128; b_mant2 = 8'd42; b_mant3 = 8'd28;
a_exp0 = 10'd672; a_exp1 = 10'd918; a_exp2 = 10'd628; a_exp3 = 10'd49;
b_exp0 = 10'd667; b_exp1 = 10'd851; b_exp2 = 10'd53; b_exp3 = 10'd394;
a_sign0 = 4'd1; a_sign1 = 4'd12; a_sign2 = 4'd8; a_sign3 = 4'd16;
b_sign0 = 4'd10; b_sign1 = 4'd3; b_sign2 = 4'd5; b_sign3 = 4'd5;
@(posedge clk_i);
a_mant0 = 8'd141; a_mant1 = 8'd156; a_mant2 = 8'd236; a_mant3 = 8'd239;
b_mant0 = 8'd71; b_mant1 = 8'd186; b_mant2 = 8'd235; b_mant3 = 8'd12;
a_exp0 = 10'd339; a_exp1 = 10'd177; a_exp2 = 10'd234; a_exp3 = 10'd33;
b_exp0 = 10'd872; b_exp1 = 10'd763; b_exp2 = 10'd593; b_exp3 = 10'd955;
a_sign0 = 4'd7; a_sign1 = 4'd9; a_sign2 = 4'd6; a_sign3 = 4'd3;
b_sign0 = 4'd4; b_sign1 = 4'd13; b_sign2 = 4'd7; b_sign3 = 4'd5;
@(posedge clk_i);
shared_exps0 = 8'd126;
shared_exps1 = 8'd126;
a_mant0 = 8'd144; a_mant1 = 8'd13; a_mant2 = 8'd232; a_mant3 = 8'd150;
b_mant0 = 8'd181; b_mant1 = 8'd19; b_mant2 = 8'd70; b_mant3 = 8'd212;
a_exp0 = 10'd588; a_exp1 = 10'd458; a_exp2 = 10'd54; a_exp3 = 10'd36;
b_exp0 = 10'd139; b_exp1 = 10'd4; b_exp2 = 10'd749; b_exp3 = 10'd764;
a_sign0 = 4'd14; a_sign1 = 4'd8; a_sign2 = 4'd9; a_sign3 = 4'd1;
b_sign0 = 4'd9; b_sign1 = 4'd4; b_sign2 = 4'd10; b_sign3 = 4'd3;
@(posedge clk_i);
a_mant0 = 8'd75; a_mant1 = 8'd55; a_mant2 = 8'd201; a_mant3 = 8'd120;
b_mant0 = 8'd79; b_mant1 = 8'd10; b_mant2 = 8'd5; b_mant3 = 8'd156;
a_exp0 = 10'd208; a_exp1 = 10'd769; a_exp2 = 10'd417; a_exp3 = 10'd398;
b_exp0 = 10'd623; b_exp1 = 10'd338; b_exp2 = 10'd130; b_exp3 = 10'd676;
a_sign0 = 4'd1; a_sign1 = 4'd15; a_sign2 = 4'd8; a_sign3 = 4'd6;
b_sign0 = 4'd0; b_sign1 = 4'd5; b_sign2 = 4'd14; b_sign3 = 4'd15;
@(posedge clk_i);
a_mant0 = 8'd15; a_mant1 = 8'd23; a_mant2 = 8'd173; a_mant3 = 8'd50;
b_mant0 = 8'd31; b_mant1 = 8'd89; b_mant2 = 8'd190; b_mant3 = 8'd119;
a_exp0 = 10'd2; a_exp1 = 10'd524; a_exp2 = 10'd680; a_exp3 = 10'd40;
b_exp0 = 10'd878; b_exp1 = 10'd620; b_exp2 = 10'd835; b_exp3 = 10'd93;
a_sign0 = 4'd11; a_sign1 = 4'd10; a_sign2 = 4'd2; a_sign3 = 4'd8;
b_sign0 = 4'd12; b_sign1 = 4'd3; b_sign2 = 4'd14; b_sign3 = 4'd12;
@(posedge clk_i);
a_mant0 = 8'd55; a_mant1 = 8'd74; a_mant2 = 8'd118; a_mant3 = 8'd239;
b_mant0 = 8'd95; b_mant1 = 8'd6; b_mant2 = 8'd253; b_mant3 = 8'd162;
a_exp0 = 10'd679; a_exp1 = 10'd577; a_exp2 = 10'd122; a_exp3 = 10'd903;
b_exp0 = 10'd77; b_exp1 = 10'd230; b_exp2 = 10'd577; b_exp3 = 10'd383;
a_sign0 = 4'd8; a_sign1 = 4'd12; a_sign2 = 4'd16; a_sign3 = 4'd14;
b_sign0 = 4'd2; b_sign1 = 4'd6; b_sign2 = 4'd7; b_sign3 = 4'd11;
@(posedge clk_i);
a_mant0 = 8'd74; a_mant1 = 8'd122; a_mant2 = 8'd87; a_mant3 = 8'd211;
b_mant0 = 8'd86; b_mant1 = 8'd25; b_mant2 = 8'd201; b_mant3 = 8'd40;
a_exp0 = 10'd845; a_exp1 = 10'd163; a_exp2 = 10'd122; a_exp3 = 10'd178;
b_exp0 = 10'd804; b_exp1 = 10'd358; b_exp2 = 10'd574; b_exp3 = 10'd505;
a_sign0 = 4'd16; a_sign1 = 4'd9; a_sign2 = 4'd7; a_sign3 = 4'd16;
b_sign0 = 4'd14; b_sign1 = 4'd10; b_sign2 = 4'd0; b_sign3 = 4'd15;
@(posedge clk_i);
a_mant0 = 8'd117; a_mant1 = 8'd64; a_mant2 = 8'd11; a_mant3 = 8'd224;
b_mant0 = 8'd33; b_mant1 = 8'd99; b_mant2 = 8'd122; b_mant3 = 8'd72;
a_exp0 = 10'd798; a_exp1 = 10'd920; a_exp2 = 10'd41; a_exp3 = 10'd821;
b_exp0 = 10'd753; b_exp1 = 10'd231; b_exp2 = 10'd603; b_exp3 = 10'd444;
a_sign0 = 4'd12; a_sign1 = 4'd7; a_sign2 = 4'd0; a_sign3 = 4'd1;
b_sign0 = 4'd0; b_sign1 = 4'd0; b_sign2 = 4'd15; b_sign3 = 4'd9;
@(posedge clk_i);
a_mant0 = 8'd208; a_mant1 = 8'd48; a_mant2 = 8'd39; a_mant3 = 8'd0;
b_mant0 = 8'd56; b_mant1 = 8'd152; b_mant2 = 8'd141; b_mant3 = 8'd45;
a_exp0 = 10'd819; a_exp1 = 10'd572; a_exp2 = 10'd755; a_exp3 = 10'd37;
b_exp0 = 10'd852; b_exp1 = 10'd366; b_exp2 = 10'd885; b_exp3 = 10'd942;
a_sign0 = 4'd3; a_sign1 = 4'd15; a_sign2 = 4'd9; a_sign3 = 4'd6;
b_sign0 = 4'd0; b_sign1 = 4'd14; b_sign2 = 4'd9; b_sign3 = 4'd16;
@(posedge clk_i);
a_mant0 = 8'd203; a_mant1 = 8'd221; a_mant2 = 8'd94; a_mant3 = 8'd200;
b_mant0 = 8'd140; b_mant1 = 8'd206; b_mant2 = 8'd199; b_mant3 = 8'd101;
a_exp0 = 10'd399; a_exp1 = 10'd375; a_exp2 = 10'd230; a_exp3 = 10'd791;
b_exp0 = 10'd188; b_exp1 = 10'd205; b_exp2 = 10'd704; b_exp3 = 10'd312;
a_sign0 = 4'd10; a_sign1 = 4'd3; a_sign2 = 4'd14; a_sign3 = 4'd0;
b_sign0 = 4'd2; b_sign1 = 4'd16; b_sign2 = 4'd12; b_sign3 = 4'd0;
@(posedge clk_i);
shared_exps0 = 8'd128;
shared_exps1 = 8'd108;
rstn = 0;
@(posedge clk_i);
rstn = 1;
a_mant0 = 8'd184; a_mant1 = 8'd113; a_mant2 = 8'd111; a_mant3 = 8'd39;
b_mant0 = 8'd253; b_mant1 = 8'd135; b_mant2 = 8'd51; b_mant3 = 8'd36;
a_exp0 = 10'd1010; a_exp1 = 10'd330; a_exp2 = 10'd680; a_exp3 = 10'd385;
b_exp0 = 10'd448; b_exp1 = 10'd561; b_exp2 = 10'd835; b_exp3 = 10'd707;
a_sign0 = 4'd1; a_sign1 = 4'd9; a_sign2 = 4'd2; a_sign3 = 4'd16;
b_sign0 = 4'd14; b_sign1 = 4'd1; b_sign2 = 4'd14; b_sign3 = 4'd12;
@(posedge clk_i);
a_mant0 = 8'd179; a_mant1 = 8'd101; a_mant2 = 8'd76; a_mant3 = 8'd52;
b_mant0 = 8'd216; b_mant1 = 8'd226; b_mant2 = 8'd111; b_mant3 = 8'd35;
a_exp0 = 10'd668; a_exp1 = 10'd901; a_exp2 = 10'd936; a_exp3 = 10'd331;
b_exp0 = 10'd812; b_exp1 = 10'd844; b_exp2 = 10'd340; b_exp3 = 10'd299;
a_sign0 = 4'd14; a_sign1 = 4'd3; a_sign2 = 4'd13; a_sign3 = 4'd7;
b_sign0 = 4'd16; b_sign1 = 4'd4; b_sign2 = 4'd5; b_sign3 = 4'd5;
@(posedge clk_i);
a_mant0 = 8'd128; a_mant1 = 8'd191; a_mant2 = 8'd87; a_mant3 = 8'd233;
b_mant0 = 8'd97; b_mant1 = 8'd42; b_mant2 = 8'd107; b_mant3 = 8'd180;
a_exp0 = 10'd203; a_exp1 = 10'd350; a_exp2 = 10'd749; a_exp3 = 10'd720;
b_exp0 = 10'd367; b_exp1 = 10'd564; b_exp2 = 10'd891; b_exp3 = 10'd118;
a_sign0 = 4'd4; a_sign1 = 4'd9; a_sign2 = 4'd15; a_sign3 = 4'd5;
b_sign0 = 4'd9; b_sign1 = 4'd14; b_sign2 = 4'd6; b_sign3 = 4'd7;
@(posedge clk_i);
a_mant0 = 8'd51; a_mant1 = 8'd86; a_mant2 = 8'd181; a_mant3 = 8'd148;
b_mant0 = 8'd182; b_mant1 = 8'd197; b_mant2 = 8'd98; b_mant3 = 8'd142;
a_exp0 = 10'd887; a_exp1 = 10'd277; a_exp2 = 10'd195; a_exp3 = 10'd600;
b_exp0 = 10'd721; b_exp1 = 10'd455; b_exp2 = 10'd299; b_exp3 = 10'd392;
a_sign0 = 4'd12; a_sign1 = 4'd7; a_sign2 = 4'd1; a_sign3 = 4'd13;
b_sign0 = 4'd7; b_sign1 = 4'd4; b_sign2 = 4'd10; b_sign3 = 4'd11;
@(posedge clk_i);
a_mant0 = 8'd48; a_mant1 = 8'd186; a_mant2 = 8'd234; a_mant3 = 8'd33;
b_mant0 = 8'd224; b_mant1 = 8'd215; b_mant2 = 8'd69; b_mant3 = 8'd150;
a_exp0 = 10'd17; a_exp1 = 10'd744; a_exp2 = 10'd286; a_exp3 = 10'd999;
b_exp0 = 10'd220; b_exp1 = 10'd543; b_exp2 = 10'd635; b_exp3 = 10'd757;
a_sign0 = 4'd3; a_sign1 = 4'd12; a_sign2 = 4'd2; a_sign3 = 4'd8;
b_sign0 = 4'd1; b_sign1 = 4'd4; b_sign2 = 4'd13; b_sign3 = 4'd14;
@(posedge clk_i);
a_mant0 = 8'd160; a_mant1 = 8'd126; a_mant2 = 8'd225; a_mant3 = 8'd206;
b_mant0 = 8'd192; b_mant1 = 8'd21; b_mant2 = 8'd210; b_mant3 = 8'd115;
a_exp0 = 10'd864; a_exp1 = 10'd296; a_exp2 = 10'd747; a_exp3 = 10'd423;
b_exp0 = 10'd1016; b_exp1 = 10'd902; b_exp2 = 10'd101; b_exp3 = 10'd959;
a_sign0 = 4'd15; a_sign1 = 4'd15; a_sign2 = 4'd6; a_sign3 = 4'd1;
b_sign0 = 4'd1; b_sign1 = 4'd14; b_sign2 = 4'd15; b_sign3 = 4'd10;
@(posedge clk_i);
a_mant0 = 8'd126; a_mant1 = 8'd139; a_mant2 = 8'd115; a_mant3 = 8'd151;
b_mant0 = 8'd69; b_mant1 = 8'd47; b_mant2 = 8'd186; b_mant3 = 8'd84;
a_exp0 = 10'd654; a_exp1 = 10'd844; a_exp2 = 10'd619; a_exp3 = 10'd856;
b_exp0 = 10'd583; b_exp1 = 10'd736; b_exp2 = 10'd578; b_exp3 = 10'd926;
a_sign0 = 4'd16; a_sign1 = 4'd6; a_sign2 = 4'd9; a_sign3 = 4'd9;
b_sign0 = 4'd8; b_sign1 = 4'd9; b_sign2 = 4'd0; b_sign3 = 4'd7;
@(posedge clk_i);
shared_exps0 = 8'd145;
shared_exps1 = 8'd117;
a_mant0 = 8'd58; a_mant1 = 8'd31; a_mant2 = 8'd17; a_mant3 = 8'd250;
b_mant0 = 8'd185; b_mant1 = 8'd12; b_mant2 = 8'd175; b_mant3 = 8'd221;
a_exp0 = 10'd913; a_exp1 = 10'd721; a_exp2 = 10'd365; a_exp3 = 10'd677;
b_exp0 = 10'd923; b_exp1 = 10'd5; b_exp2 = 10'd409; b_exp3 = 10'd795;
a_sign0 = 4'd11; a_sign1 = 4'd12; a_sign2 = 4'd4; a_sign3 = 4'd16;
b_sign0 = 4'd14; b_sign1 = 4'd11; b_sign2 = 4'd14; b_sign3 = 4'd16;
@(posedge clk_i);
a_mant0 = 8'd23; a_mant1 = 8'd169; a_mant2 = 8'd201; a_mant3 = 8'd192;
b_mant0 = 8'd138; b_mant1 = 8'd51; b_mant2 = 8'd8; b_mant3 = 8'd27;
a_exp0 = 10'd668; a_exp1 = 10'd345; a_exp2 = 10'd445; a_exp3 = 10'd95;
b_exp0 = 10'd322; b_exp1 = 10'd625; b_exp2 = 10'd539; b_exp3 = 10'd338;
a_sign0 = 4'd7; a_sign1 = 4'd14; a_sign2 = 4'd14; a_sign3 = 4'd2;
b_sign0 = 4'd9; b_sign1 = 4'd11; b_sign2 = 4'd6; b_sign3 = 4'd11;
@(posedge clk_i);
a_mant0 = 8'd171; a_mant1 = 8'd30; a_mant2 = 8'd97; a_mant3 = 8'd120;
b_mant0 = 8'd27; b_mant1 = 8'd212; b_mant2 = 8'd254; b_mant3 = 8'd143;
a_exp0 = 10'd256; a_exp1 = 10'd884; a_exp2 = 10'd134; a_exp3 = 10'd970;
b_exp0 = 10'd1000; b_exp1 = 10'd807; b_exp2 = 10'd644; b_exp3 = 10'd254;
a_sign0 = 4'd3; a_sign1 = 4'd5; a_sign2 = 4'd2; a_sign3 = 4'd6;
b_sign0 = 4'd2; b_sign1 = 4'd12; b_sign2 = 4'd13; b_sign3 = 4'd3;
@(posedge clk_i);
a_mant0 = 8'd241; a_mant1 = 8'd160; a_mant2 = 8'd177; a_mant3 = 8'd111;
b_mant0 = 8'd28; b_mant1 = 8'd24; b_mant2 = 8'd34; b_mant3 = 8'd71;
a_exp0 = 10'd476; a_exp1 = 10'd445; a_exp2 = 10'd103; a_exp3 = 10'd316;
b_exp0 = 10'd372; b_exp1 = 10'd834; b_exp2 = 10'd100; b_exp3 = 10'd257;
a_sign0 = 4'd13; a_sign1 = 4'd10; a_sign2 = 4'd12; a_sign3 = 4'd14;
b_sign0 = 4'd11; b_sign1 = 4'd13; b_sign2 = 4'd16; b_sign3 = 4'd3;
@(posedge clk_i);
a_mant0 = 8'd57; a_mant1 = 8'd33; a_mant2 = 8'd154; a_mant3 = 8'd161;
b_mant0 = 8'd16; b_mant1 = 8'd67; b_mant2 = 8'd180; b_mant3 = 8'd90;
a_exp0 = 10'd319; a_exp1 = 10'd1021; a_exp2 = 10'd618; a_exp3 = 10'd830;
b_exp0 = 10'd848; b_exp1 = 10'd553; b_exp2 = 10'd754; b_exp3 = 10'd559;
a_sign0 = 4'd12; a_sign1 = 4'd8; a_sign2 = 4'd8; a_sign3 = 4'd15;
b_sign0 = 4'd14; b_sign1 = 4'd4; b_sign2 = 4'd8; b_sign3 = 4'd3;
@(posedge clk_i);
a_mant0 = 8'd163; a_mant1 = 8'd39; a_mant2 = 8'd185; a_mant3 = 8'd61;
b_mant0 = 8'd132; b_mant1 = 8'd240; b_mant2 = 8'd150; b_mant3 = 8'd113;
a_exp0 = 10'd687; a_exp1 = 10'd443; a_exp2 = 10'd232; a_exp3 = 10'd191;
b_exp0 = 10'd509; b_exp1 = 10'd579; b_exp2 = 10'd631; b_exp3 = 10'd533;
a_sign0 = 4'd12; a_sign1 = 4'd10; a_sign2 = 4'd6; a_sign3 = 4'd5;
b_sign0 = 4'd7; b_sign1 = 4'd3; b_sign2 = 4'd7; b_sign3 = 4'd10;
@(posedge clk_i);
a_mant0 = 8'd48; a_mant1 = 8'd107; a_mant2 = 8'd75; a_mant3 = 8'd53;
b_mant0 = 8'd19; b_mant1 = 8'd117; b_mant2 = 8'd169; b_mant3 = 8'd1;
a_exp0 = 10'd96; a_exp1 = 10'd989; a_exp2 = 10'd578; a_exp3 = 10'd826;
b_exp0 = 10'd402; b_exp1 = 10'd759; b_exp2 = 10'd744; b_exp3 = 10'd317;
a_sign0 = 4'd13; a_sign1 = 4'd9; a_sign2 = 4'd11; a_sign3 = 4'd13;
b_sign0 = 4'd5; b_sign1 = 4'd2; b_sign2 = 4'd13; b_sign3 = 4'd3;
@(posedge clk_i);
a_mant0 = 8'd97; a_mant1 = 8'd27; a_mant2 = 8'd119; a_mant3 = 8'd228;
b_mant0 = 8'd225; b_mant1 = 8'd97; b_mant2 = 8'd50; b_mant3 = 8'd72;
a_exp0 = 10'd991; a_exp1 = 10'd719; a_exp2 = 10'd252; a_exp3 = 10'd239;
b_exp0 = 10'd803; b_exp1 = 10'd520; b_exp2 = 10'd253; b_exp3 = 10'd722;
a_sign0 = 4'd0; a_sign1 = 4'd6; a_sign2 = 4'd3; a_sign3 = 4'd7;
b_sign0 = 4'd10; b_sign1 = 4'd0; b_sign2 = 4'd5; b_sign3 = 4'd7;
@(posedge clk_i);
shared_exps0 = 8'd117;
shared_exps1 = 8'd157;
a_mant0 = 8'd142; a_mant1 = 8'd147; a_mant2 = 8'd222; a_mant3 = 8'd201;
b_mant0 = 8'd80; b_mant1 = 8'd96; b_mant2 = 8'd0; b_mant3 = 8'd124;
a_exp0 = 10'd89; a_exp1 = 10'd430; a_exp2 = 10'd502; a_exp3 = 10'd959;
b_exp0 = 10'd37; b_exp1 = 10'd433; b_exp2 = 10'd105; b_exp3 = 10'd606;
a_sign0 = 4'd0; a_sign1 = 4'd0; a_sign2 = 4'd3; a_sign3 = 4'd2;
b_sign0 = 4'd16; b_sign1 = 4'd4; b_sign2 = 4'd14; b_sign3 = 4'd16;
@(posedge clk_i);
a_mant0 = 8'd39; a_mant1 = 8'd219; a_mant2 = 8'd201; a_mant3 = 8'd151;
b_mant0 = 8'd247; b_mant1 = 8'd5; b_mant2 = 8'd107; b_mant3 = 8'd69;
a_exp0 = 10'd797; a_exp1 = 10'd584; a_exp2 = 10'd742; a_exp3 = 10'd627;
b_exp0 = 10'd739; b_exp1 = 10'd168; b_exp2 = 10'd451; b_exp3 = 10'd715;
a_sign0 = 4'd12; a_sign1 = 4'd7; a_sign2 = 4'd11; a_sign3 = 4'd7;
b_sign0 = 4'd8; b_sign1 = 4'd15; b_sign2 = 4'd13; b_sign3 = 4'd16;
@(posedge clk_i);
a_mant0 = 8'd166; a_mant1 = 8'd110; a_mant2 = 8'd39; a_mant3 = 8'd58;
b_mant0 = 8'd2; b_mant1 = 8'd97; b_mant2 = 8'd53; b_mant3 = 8'd87;
a_exp0 = 10'd532; a_exp1 = 10'd983; a_exp2 = 10'd797; a_exp3 = 10'd969;
b_exp0 = 10'd365; b_exp1 = 10'd989; b_exp2 = 10'd978; b_exp3 = 10'd559;
a_sign0 = 4'd4; a_sign1 = 4'd14; a_sign2 = 4'd1; a_sign3 = 4'd7;
b_sign0 = 4'd15; b_sign1 = 4'd6; b_sign2 = 4'd3; b_sign3 = 4'd2;
@(posedge clk_i);
a_mant0 = 8'd167; a_mant1 = 8'd69; a_mant2 = 8'd110; a_mant3 = 8'd164;
b_mant0 = 8'd116; b_mant1 = 8'd18; b_mant2 = 8'd124; b_mant3 = 8'd216;
a_exp0 = 10'd380; a_exp1 = 10'd159; a_exp2 = 10'd657; a_exp3 = 10'd679;
b_exp0 = 10'd836; b_exp1 = 10'd188; b_exp2 = 10'd91; b_exp3 = 10'd1014;
a_sign0 = 4'd12; a_sign1 = 4'd16; a_sign2 = 4'd0; a_sign3 = 4'd13;
b_sign0 = 4'd2; b_sign1 = 4'd4; b_sign2 = 4'd4; b_sign3 = 4'd8;
@(posedge clk_i);
a_mant0 = 8'd2; a_mant1 = 8'd148; a_mant2 = 8'd135; a_mant3 = 8'd98;
b_mant0 = 8'd53; b_mant1 = 8'd74; b_mant2 = 8'd26; b_mant3 = 8'd146;
a_exp0 = 10'd786; a_exp1 = 10'd605; a_exp2 = 10'd807; a_exp3 = 10'd611;
b_exp0 = 10'd878; b_exp1 = 10'd476; b_exp2 = 10'd742; b_exp3 = 10'd108;
a_sign0 = 4'd5; a_sign1 = 4'd2; a_sign2 = 4'd9; a_sign3 = 4'd4;
b_sign0 = 4'd1; b_sign1 = 4'd1; b_sign2 = 4'd10; b_sign3 = 4'd2;
@(posedge clk_i);
a_mant0 = 8'd235; a_mant1 = 8'd77; a_mant2 = 8'd27; a_mant3 = 8'd17;
b_mant0 = 8'd28; b_mant1 = 8'd0; b_mant2 = 8'd13; b_mant3 = 8'd56;
a_exp0 = 10'd112; a_exp1 = 10'd285; a_exp2 = 10'd809; a_exp3 = 10'd14;
b_exp0 = 10'd720; b_exp1 = 10'd893; b_exp2 = 10'd152; b_exp3 = 10'd1009;
a_sign0 = 4'd8; a_sign1 = 4'd4; a_sign2 = 4'd14; a_sign3 = 4'd16;
b_sign0 = 4'd15; b_sign1 = 4'd1; b_sign2 = 4'd15; b_sign3 = 4'd11;
@(posedge clk_i);
a_mant0 = 8'd5; a_mant1 = 8'd89; a_mant2 = 8'd121; a_mant3 = 8'd238;
b_mant0 = 8'd60; b_mant1 = 8'd122; b_mant2 = 8'd179; b_mant3 = 8'd136;
a_exp0 = 10'd864; a_exp1 = 10'd501; a_exp2 = 10'd913; a_exp3 = 10'd818;
b_exp0 = 10'd284; b_exp1 = 10'd25; b_exp2 = 10'd947; b_exp3 = 10'd771;
a_sign0 = 4'd9; a_sign1 = 4'd8; a_sign2 = 4'd10; a_sign3 = 4'd5;
b_sign0 = 4'd7; b_sign1 = 4'd14; b_sign2 = 4'd13; b_sign3 = 4'd9;
@(posedge clk_i);
a_mant0 = 8'd57; a_mant1 = 8'd2; a_mant2 = 8'd73; a_mant3 = 8'd146;
b_mant0 = 8'd22; b_mant1 = 8'd206; b_mant2 = 8'd117; b_mant3 = 8'd81;
a_exp0 = 10'd695; a_exp1 = 10'd611; a_exp2 = 10'd770; a_exp3 = 10'd973;
b_exp0 = 10'd308; b_exp1 = 10'd9; b_exp2 = 10'd49; b_exp3 = 10'd292;
a_sign0 = 4'd14; a_sign1 = 4'd3; a_sign2 = 4'd15; a_sign3 = 4'd15;
b_sign0 = 4'd10; b_sign1 = 4'd10; b_sign2 = 4'd13; b_sign3 = 4'd3;
@(posedge clk_i);
shared_exps0 = 8'd124;
shared_exps1 = 8'd153;
a_mant0 = 8'd225; a_mant1 = 8'd5; a_mant2 = 8'd140; a_mant3 = 8'd92;
b_mant0 = 8'd116; b_mant1 = 8'd116; b_mant2 = 8'd31; b_mant3 = 8'd7;
a_exp0 = 10'd927; a_exp1 = 10'd591; a_exp2 = 10'd642; a_exp3 = 10'd378;
b_exp0 = 10'd136; b_exp1 = 10'd147; b_exp2 = 10'd315; b_exp3 = 10'd178;
a_sign0 = 4'd14; a_sign1 = 4'd4; a_sign2 = 4'd10; a_sign3 = 4'd7;
b_sign0 = 4'd14; b_sign1 = 4'd11; b_sign2 = 4'd8; b_sign3 = 4'd7;
@(posedge clk_i);
a_mant0 = 8'd84; a_mant1 = 8'd207; a_mant2 = 8'd65; a_mant3 = 8'd189;
b_mant0 = 8'd119; b_mant1 = 8'd224; b_mant2 = 8'd16; b_mant3 = 8'd224;
a_exp0 = 10'd29; a_exp1 = 10'd257; a_exp2 = 10'd476; a_exp3 = 10'd80;
b_exp0 = 10'd305; b_exp1 = 10'd464; b_exp2 = 10'd943; b_exp3 = 10'd1009;
a_sign0 = 4'd11; a_sign1 = 4'd2; a_sign2 = 4'd2; a_sign3 = 4'd16;
b_sign0 = 4'd15; b_sign1 = 4'd3; b_sign2 = 4'd12; b_sign3 = 4'd3;
@(posedge clk_i);
a_mant0 = 8'd55; a_mant1 = 8'd195; a_mant2 = 8'd127; a_mant3 = 8'd187;
b_mant0 = 8'd158; b_mant1 = 8'd174; b_mant2 = 8'd75; b_mant3 = 8'd222;
a_exp0 = 10'd719; a_exp1 = 10'd447; a_exp2 = 10'd131; a_exp3 = 10'd779;
b_exp0 = 10'd676; b_exp1 = 10'd761; b_exp2 = 10'd682; b_exp3 = 10'd990;
a_sign0 = 4'd15; a_sign1 = 4'd15; a_sign2 = 4'd0; a_sign3 = 4'd4;
b_sign0 = 4'd0; b_sign1 = 4'd11; b_sign2 = 4'd8; b_sign3 = 4'd3;
@(posedge clk_i);
a_mant0 = 8'd177; a_mant1 = 8'd43; a_mant2 = 8'd224; a_mant3 = 8'd9;
b_mant0 = 8'd42; b_mant1 = 8'd249; b_mant2 = 8'd174; b_mant3 = 8'd180;
a_exp0 = 10'd681; a_exp1 = 10'd493; a_exp2 = 10'd364; a_exp3 = 10'd745;
b_exp0 = 10'd340; b_exp1 = 10'd654; b_exp2 = 10'd631; b_exp3 = 10'd560;
a_sign0 = 4'd7; a_sign1 = 4'd8; a_sign2 = 4'd4; a_sign3 = 4'd3;
b_sign0 = 4'd13; b_sign1 = 4'd6; b_sign2 = 4'd2; b_sign3 = 4'd12;
@(posedge clk_i);
a_mant0 = 8'd122; a_mant1 = 8'd98; a_mant2 = 8'd143; a_mant3 = 8'd162;
b_mant0 = 8'd247; b_mant1 = 8'd142; b_mant2 = 8'd23; b_mant3 = 8'd87;
a_exp0 = 10'd209; a_exp1 = 10'd33; a_exp2 = 10'd525; a_exp3 = 10'd872;
b_exp0 = 10'd555; b_exp1 = 10'd185; b_exp2 = 10'd758; b_exp3 = 10'd907;
a_sign0 = 4'd6; a_sign1 = 4'd0; a_sign2 = 4'd13; a_sign3 = 4'd12;
b_sign0 = 4'd1; b_sign1 = 4'd1; b_sign2 = 4'd10; b_sign3 = 4'd13;
@(posedge clk_i);
a_mant0 = 8'd244; a_mant1 = 8'd201; a_mant2 = 8'd115; a_mant3 = 8'd171;
b_mant0 = 8'd98; b_mant1 = 8'd249; b_mant2 = 8'd129; b_mant3 = 8'd208;
a_exp0 = 10'd491; a_exp1 = 10'd501; a_exp2 = 10'd114; a_exp3 = 10'd56;
b_exp0 = 10'd802; b_exp1 = 10'd649; b_exp2 = 10'd800; b_exp3 = 10'd649;
a_sign0 = 4'd14; a_sign1 = 4'd7; a_sign2 = 4'd2; a_sign3 = 4'd8;
b_sign0 = 4'd9; b_sign1 = 4'd4; b_sign2 = 4'd16; b_sign3 = 4'd5;
@(posedge clk_i);
a_mant0 = 8'd25; a_mant1 = 8'd60; a_mant2 = 8'd17; a_mant3 = 8'd151;
b_mant0 = 8'd49; b_mant1 = 8'd25; b_mant2 = 8'd180; b_mant3 = 8'd131;
a_exp0 = 10'd306; a_exp1 = 10'd338; a_exp2 = 10'd729; a_exp3 = 10'd680;
b_exp0 = 10'd911; b_exp1 = 10'd273; b_exp2 = 10'd235; b_exp3 = 10'd105;
a_sign0 = 4'd0; a_sign1 = 4'd11; a_sign2 = 4'd11; a_sign3 = 4'd9;
b_sign0 = 4'd4; b_sign1 = 4'd6; b_sign2 = 4'd1; b_sign3 = 4'd4;
@(posedge clk_i);
a_mant0 = 8'd190; a_mant1 = 8'd51; a_mant2 = 8'd217; a_mant3 = 8'd33;
b_mant0 = 8'd124; b_mant1 = 8'd147; b_mant2 = 8'd234; b_mant3 = 8'd242;
a_exp0 = 10'd526; a_exp1 = 10'd337; a_exp2 = 10'd315; a_exp3 = 10'd255;
b_exp0 = 10'd273; b_exp1 = 10'd727; b_exp2 = 10'd744; b_exp3 = 10'd1020;
a_sign0 = 4'd6; a_sign1 = 4'd3; a_sign2 = 4'd11; a_sign3 = 4'd11;
b_sign0 = 4'd4; b_sign1 = 4'd14; b_sign2 = 4'd2; b_sign3 = 4'd11;
@(posedge clk_i);
shared_exps0 = 8'd105;
shared_exps1 = 8'd120;
rstn = 0;
@(posedge clk_i);
rstn = 1;
a_mant0 = 8'd69; a_mant1 = 8'd187; a_mant2 = 8'd157; a_mant3 = 8'd69;
b_mant0 = 8'd103; b_mant1 = 8'd245; b_mant2 = 8'd47; b_mant3 = 8'd0;
a_exp0 = 10'd603; a_exp1 = 10'd595; a_exp2 = 10'd819; a_exp3 = 10'd929;
b_exp0 = 10'd641; b_exp1 = 10'd120; b_exp2 = 10'd782; b_exp3 = 10'd252;
a_sign0 = 4'd9; a_sign1 = 4'd15; a_sign2 = 4'd2; a_sign3 = 4'd6;
b_sign0 = 4'd13; b_sign1 = 4'd9; b_sign2 = 4'd9; b_sign3 = 4'd11;
@(posedge clk_i);
a_mant0 = 8'd22; a_mant1 = 8'd141; a_mant2 = 8'd252; a_mant3 = 8'd37;
b_mant0 = 8'd199; b_mant1 = 8'd90; b_mant2 = 8'd153; b_mant3 = 8'd197;
a_exp0 = 10'd462; a_exp1 = 10'd825; a_exp2 = 10'd355; a_exp3 = 10'd480;
b_exp0 = 10'd128; b_exp1 = 10'd563; b_exp2 = 10'd307; b_exp3 = 10'd296;
a_sign0 = 4'd12; a_sign1 = 4'd7; a_sign2 = 4'd1; a_sign3 = 4'd3;
b_sign0 = 4'd3; b_sign1 = 4'd15; b_sign2 = 4'd9; b_sign3 = 4'd2;
@(posedge clk_i);
a_mant0 = 8'd135; a_mant1 = 8'd189; a_mant2 = 8'd184; a_mant3 = 8'd209;
b_mant0 = 8'd219; b_mant1 = 8'd86; b_mant2 = 8'd31; b_mant3 = 8'd44;
a_exp0 = 10'd441; a_exp1 = 10'd1001; a_exp2 = 10'd76; a_exp3 = 10'd1002;
b_exp0 = 10'd33; b_exp1 = 10'd429; b_exp2 = 10'd893; b_exp3 = 10'd293;
a_sign0 = 4'd6; a_sign1 = 4'd15; a_sign2 = 4'd2; a_sign3 = 4'd8;
b_sign0 = 4'd5; b_sign1 = 4'd0; b_sign2 = 4'd5; b_sign3 = 4'd6;
@(posedge clk_i);
a_mant0 = 8'd10; a_mant1 = 8'd110; a_mant2 = 8'd89; a_mant3 = 8'd38;
b_mant0 = 8'd173; b_mant1 = 8'd174; b_mant2 = 8'd5; b_mant3 = 8'd154;
a_exp0 = 10'd959; a_exp1 = 10'd338; a_exp2 = 10'd941; a_exp3 = 10'd810;
b_exp0 = 10'd970; b_exp1 = 10'd990; b_exp2 = 10'd84; b_exp3 = 10'd504;
a_sign0 = 4'd16; a_sign1 = 4'd6; a_sign2 = 4'd8; a_sign3 = 4'd5;
b_sign0 = 4'd4; b_sign1 = 4'd10; b_sign2 = 4'd9; b_sign3 = 4'd10;
@(posedge clk_i);
a_mant0 = 8'd143; a_mant1 = 8'd162; a_mant2 = 8'd35; a_mant3 = 8'd103;
b_mant0 = 8'd65; b_mant1 = 8'd102; b_mant2 = 8'd61; b_mant3 = 8'd164;
a_exp0 = 10'd426; a_exp1 = 10'd364; a_exp2 = 10'd1023; a_exp3 = 10'd736;
b_exp0 = 10'd59; b_exp1 = 10'd554; b_exp2 = 10'd529; b_exp3 = 10'd18;
a_sign0 = 4'd3; a_sign1 = 4'd4; a_sign2 = 4'd9; a_sign3 = 4'd4;
b_sign0 = 4'd15; b_sign1 = 4'd8; b_sign2 = 4'd2; b_sign3 = 4'd4;
@(posedge clk_i);
a_mant0 = 8'd56; a_mant1 = 8'd174; a_mant2 = 8'd79; a_mant3 = 8'd65;
b_mant0 = 8'd81; b_mant1 = 8'd9; b_mant2 = 8'd209; b_mant3 = 8'd205;
a_exp0 = 10'd882; a_exp1 = 10'd96; a_exp2 = 10'd582; a_exp3 = 10'd789;
b_exp0 = 10'd699; b_exp1 = 10'd488; b_exp2 = 10'd356; b_exp3 = 10'd48;
a_sign0 = 4'd3; a_sign1 = 4'd2; a_sign2 = 4'd2; a_sign3 = 4'd8;
b_sign0 = 4'd9; b_sign1 = 4'd10; b_sign2 = 4'd11; b_sign3 = 4'd11;
@(posedge clk_i);
a_mant0 = 8'd63; a_mant1 = 8'd97; a_mant2 = 8'd12; a_mant3 = 8'd122;
b_mant0 = 8'd62; b_mant1 = 8'd122; b_mant2 = 8'd154; b_mant3 = 8'd81;
a_exp0 = 10'd445; a_exp1 = 10'd74; a_exp2 = 10'd347; a_exp3 = 10'd184;
b_exp0 = 10'd494; b_exp1 = 10'd276; b_exp2 = 10'd317; b_exp3 = 10'd649;
a_sign0 = 4'd2; a_sign1 = 4'd16; a_sign2 = 4'd5; a_sign3 = 4'd10;
b_sign0 = 4'd10; b_sign1 = 4'd9; b_sign2 = 4'd9; b_sign3 = 4'd15;
@(posedge clk_i);
shared_exps0 = 8'd150;
shared_exps1 = 8'd120;
a_mant0 = 8'd13; a_mant1 = 8'd159; a_mant2 = 8'd83; a_mant3 = 8'd232;
b_mant0 = 8'd122; b_mant1 = 8'd127; b_mant2 = 8'd66; b_mant3 = 8'd212;
a_exp0 = 10'd808; a_exp1 = 10'd334; a_exp2 = 10'd852; a_exp3 = 10'd171;
b_exp0 = 10'd441; b_exp1 = 10'd345; b_exp2 = 10'd143; b_exp3 = 10'd461;
a_sign0 = 4'd13; a_sign1 = 4'd7; a_sign2 = 4'd7; a_sign3 = 4'd14;
b_sign0 = 4'd11; b_sign1 = 4'd1; b_sign2 = 4'd15; b_sign3 = 4'd11;
@(posedge clk_i);
a_mant0 = 8'd124; a_mant1 = 8'd33; a_mant2 = 8'd153; a_mant3 = 8'd155;
b_mant0 = 8'd41; b_mant1 = 8'd2; b_mant2 = 8'd67; b_mant3 = 8'd26;
a_exp0 = 10'd698; a_exp1 = 10'd159; a_exp2 = 10'd938; a_exp3 = 10'd724;
b_exp0 = 10'd43; b_exp1 = 10'd258; b_exp2 = 10'd535; b_exp3 = 10'd638;
a_sign0 = 4'd15; a_sign1 = 4'd8; a_sign2 = 4'd15; a_sign3 = 4'd14;
b_sign0 = 4'd10; b_sign1 = 4'd12; b_sign2 = 4'd13; b_sign3 = 4'd8;
@(posedge clk_i);
a_mant0 = 8'd78; a_mant1 = 8'd54; a_mant2 = 8'd65; a_mant3 = 8'd128;
b_mant0 = 8'd97; b_mant1 = 8'd3; b_mant2 = 8'd191; b_mant3 = 8'd221;
a_exp0 = 10'd763; a_exp1 = 10'd833; a_exp2 = 10'd625; a_exp3 = 10'd617;
b_exp0 = 10'd599; b_exp1 = 10'd74; b_exp2 = 10'd432; b_exp3 = 10'd374;
a_sign0 = 4'd3; a_sign1 = 4'd14; a_sign2 = 4'd15; a_sign3 = 4'd5;
b_sign0 = 4'd16; b_sign1 = 4'd8; b_sign2 = 4'd4; b_sign3 = 4'd11;
@(posedge clk_i);
a_mant0 = 8'd119; a_mant1 = 8'd162; a_mant2 = 8'd148; a_mant3 = 8'd149;
b_mant0 = 8'd126; b_mant1 = 8'd251; b_mant2 = 8'd186; b_mant3 = 8'd202;
a_exp0 = 10'd549; a_exp1 = 10'd894; a_exp2 = 10'd313; a_exp3 = 10'd153;
b_exp0 = 10'd76; b_exp1 = 10'd383; b_exp2 = 10'd559; b_exp3 = 10'd921;
a_sign0 = 4'd16; a_sign1 = 4'd2; a_sign2 = 4'd12; a_sign3 = 4'd0;
b_sign0 = 4'd14; b_sign1 = 4'd8; b_sign2 = 4'd13; b_sign3 = 4'd14;
@(posedge clk_i);
a_mant0 = 8'd115; a_mant1 = 8'd128; a_mant2 = 8'd84; a_mant3 = 8'd151;
b_mant0 = 8'd113; b_mant1 = 8'd58; b_mant2 = 8'd219; b_mant3 = 8'd96;
a_exp0 = 10'd657; a_exp1 = 10'd514; a_exp2 = 10'd717; a_exp3 = 10'd746;
b_exp0 = 10'd250; b_exp1 = 10'd722; b_exp2 = 10'd751; b_exp3 = 10'd791;
a_sign0 = 4'd2; a_sign1 = 4'd2; a_sign2 = 4'd7; a_sign3 = 4'd16;
b_sign0 = 4'd6; b_sign1 = 4'd14; b_sign2 = 4'd1; b_sign3 = 4'd3;
@(posedge clk_i);
a_mant0 = 8'd230; a_mant1 = 8'd96; a_mant2 = 8'd30; a_mant3 = 8'd140;
b_mant0 = 8'd245; b_mant1 = 8'd254; b_mant2 = 8'd226; b_mant3 = 8'd182;
a_exp0 = 10'd227; a_exp1 = 10'd589; a_exp2 = 10'd904; a_exp3 = 10'd288;
b_exp0 = 10'd916; b_exp1 = 10'd141; b_exp2 = 10'd11; b_exp3 = 10'd291;
a_sign0 = 4'd1; a_sign1 = 4'd8; a_sign2 = 4'd8; a_sign3 = 4'd16;
b_sign0 = 4'd12; b_sign1 = 4'd11; b_sign2 = 4'd5; b_sign3 = 4'd4;
@(posedge clk_i);
a_mant0 = 8'd33; a_mant1 = 8'd26; a_mant2 = 8'd243; a_mant3 = 8'd185;
b_mant0 = 8'd50; b_mant1 = 8'd154; b_mant2 = 8'd63; b_mant3 = 8'd120;
a_exp0 = 10'd871; a_exp1 = 10'd442; a_exp2 = 10'd449; a_exp3 = 10'd916;
b_exp0 = 10'd626; b_exp1 = 10'd36; b_exp2 = 10'd994; b_exp3 = 10'd188;
a_sign0 = 4'd5; a_sign1 = 4'd5; a_sign2 = 4'd5; a_sign3 = 4'd12;
b_sign0 = 4'd11; b_sign1 = 4'd9; b_sign2 = 4'd5; b_sign3 = 4'd8;
@(posedge clk_i);
a_mant0 = 8'd102; a_mant1 = 8'd56; a_mant2 = 8'd92; a_mant3 = 8'd47;
b_mant0 = 8'd94; b_mant1 = 8'd142; b_mant2 = 8'd192; b_mant3 = 8'd31;
a_exp0 = 10'd838; a_exp1 = 10'd86; a_exp2 = 10'd418; a_exp3 = 10'd267;
b_exp0 = 10'd780; b_exp1 = 10'd567; b_exp2 = 10'd921; b_exp3 = 10'd231;
a_sign0 = 4'd12; a_sign1 = 4'd6; a_sign2 = 4'd3; a_sign3 = 4'd6;
b_sign0 = 4'd5; b_sign1 = 4'd15; b_sign2 = 4'd9; b_sign3 = 4'd12;
@(posedge clk_i);
shared_exps0 = 8'd146;
shared_exps1 = 8'd118;
a_mant0 = 8'd145; a_mant1 = 8'd89; a_mant2 = 8'd115; a_mant3 = 8'd91;
b_mant0 = 8'd109; b_mant1 = 8'd135; b_mant2 = 8'd56; b_mant3 = 8'd216;
a_exp0 = 10'd728; a_exp1 = 10'd329; a_exp2 = 10'd673; a_exp3 = 10'd298;
b_exp0 = 10'd620; b_exp1 = 10'd777; b_exp2 = 10'd748; b_exp3 = 10'd600;
a_sign0 = 4'd2; a_sign1 = 4'd5; a_sign2 = 4'd3; a_sign3 = 4'd2;
b_sign0 = 4'd2; b_sign1 = 4'd9; b_sign2 = 4'd4; b_sign3 = 4'd8;
@(posedge clk_i);
a_mant0 = 8'd187; a_mant1 = 8'd170; a_mant2 = 8'd127; a_mant3 = 8'd84;
b_mant0 = 8'd108; b_mant1 = 8'd154; b_mant2 = 8'd130; b_mant3 = 8'd161;
a_exp0 = 10'd563; a_exp1 = 10'd508; a_exp2 = 10'd625; a_exp3 = 10'd947;
b_exp0 = 10'd399; b_exp1 = 10'd295; b_exp2 = 10'd10; b_exp3 = 10'd881;
a_sign0 = 4'd12; a_sign1 = 4'd8; a_sign2 = 4'd13; a_sign3 = 4'd10;
b_sign0 = 4'd16; b_sign1 = 4'd0; b_sign2 = 4'd0; b_sign3 = 4'd4;
@(posedge clk_i);
a_mant0 = 8'd10; a_mant1 = 8'd102; a_mant2 = 8'd114; a_mant3 = 8'd43;
b_mant0 = 8'd147; b_mant1 = 8'd34; b_mant2 = 8'd57; b_mant3 = 8'd42;
a_exp0 = 10'd982; a_exp1 = 10'd288; a_exp2 = 10'd865; a_exp3 = 10'd544;
b_exp0 = 10'd653; b_exp1 = 10'd13; b_exp2 = 10'd647; b_exp3 = 10'd348;
a_sign0 = 4'd5; a_sign1 = 4'd7; a_sign2 = 4'd16; a_sign3 = 4'd0;
b_sign0 = 4'd1; b_sign1 = 4'd11; b_sign2 = 4'd8; b_sign3 = 4'd10;
@(posedge clk_i);
a_mant0 = 8'd47; a_mant1 = 8'd95; a_mant2 = 8'd215; a_mant3 = 8'd47;
b_mant0 = 8'd215; b_mant1 = 8'd199; b_mant2 = 8'd160; b_mant3 = 8'd4;
a_exp0 = 10'd737; a_exp1 = 10'd694; a_exp2 = 10'd943; a_exp3 = 10'd279;
b_exp0 = 10'd57; b_exp1 = 10'd811; b_exp2 = 10'd195; b_exp3 = 10'd201;
a_sign0 = 4'd14; a_sign1 = 4'd2; a_sign2 = 4'd11; a_sign3 = 4'd12;
b_sign0 = 4'd14; b_sign1 = 4'd12; b_sign2 = 4'd9; b_sign3 = 4'd14;
@(posedge clk_i);
a_mant0 = 8'd254; a_mant1 = 8'd219; a_mant2 = 8'd171; a_mant3 = 8'd114;
b_mant0 = 8'd103; b_mant1 = 8'd19; b_mant2 = 8'd106; b_mant3 = 8'd103;
a_exp0 = 10'd534; a_exp1 = 10'd557; a_exp2 = 10'd670; a_exp3 = 10'd467;
b_exp0 = 10'd774; b_exp1 = 10'd485; b_exp2 = 10'd462; b_exp3 = 10'd687;
a_sign0 = 4'd13; a_sign1 = 4'd4; a_sign2 = 4'd12; a_sign3 = 4'd7;
b_sign0 = 4'd2; b_sign1 = 4'd14; b_sign2 = 4'd4; b_sign3 = 4'd2;
@(posedge clk_i);
a_mant0 = 8'd249; a_mant1 = 8'd216; a_mant2 = 8'd21; a_mant3 = 8'd193;
b_mant0 = 8'd63; b_mant1 = 8'd121; b_mant2 = 8'd231; b_mant3 = 8'd141;
a_exp0 = 10'd942; a_exp1 = 10'd958; a_exp2 = 10'd76; a_exp3 = 10'd737;
b_exp0 = 10'd460; b_exp1 = 10'd120; b_exp2 = 10'd436; b_exp3 = 10'd600;
a_sign0 = 4'd13; a_sign1 = 4'd1; a_sign2 = 4'd12; a_sign3 = 4'd7;
b_sign0 = 4'd10; b_sign1 = 4'd7; b_sign2 = 4'd10; b_sign3 = 4'd9;
@(posedge clk_i);
a_mant0 = 8'd190; a_mant1 = 8'd135; a_mant2 = 8'd226; a_mant3 = 8'd42;
b_mant0 = 8'd112; b_mant1 = 8'd246; b_mant2 = 8'd81; b_mant3 = 8'd17;
a_exp0 = 10'd691; a_exp1 = 10'd248; a_exp2 = 10'd904; a_exp3 = 10'd853;
b_exp0 = 10'd481; b_exp1 = 10'd177; b_exp2 = 10'd801; b_exp3 = 10'd678;
a_sign0 = 4'd6; a_sign1 = 4'd1; a_sign2 = 4'd3; a_sign3 = 4'd13;
b_sign0 = 4'd1; b_sign1 = 4'd1; b_sign2 = 4'd8; b_sign3 = 4'd5;
@(posedge clk_i);
a_mant0 = 8'd166; a_mant1 = 8'd157; a_mant2 = 8'd112; a_mant3 = 8'd140;
b_mant0 = 8'd22; b_mant1 = 8'd120; b_mant2 = 8'd153; b_mant3 = 8'd27;
a_exp0 = 10'd630; a_exp1 = 10'd998; a_exp2 = 10'd557; a_exp3 = 10'd340;
b_exp0 = 10'd328; b_exp1 = 10'd28; b_exp2 = 10'd755; b_exp3 = 10'd519;
a_sign0 = 4'd3; a_sign1 = 4'd6; a_sign2 = 4'd10; a_sign3 = 4'd1;
b_sign0 = 4'd2; b_sign1 = 4'd2; b_sign2 = 4'd3; b_sign3 = 4'd16;
@(posedge clk_i);
shared_exps0 = 8'd141;
shared_exps1 = 8'd133;
a_mant0 = 8'd52; a_mant1 = 8'd72; a_mant2 = 8'd107; a_mant3 = 8'd241;
b_mant0 = 8'd42; b_mant1 = 8'd26; b_mant2 = 8'd189; b_mant3 = 8'd169;
a_exp0 = 10'd604; a_exp1 = 10'd375; a_exp2 = 10'd218; a_exp3 = 10'd255;
b_exp0 = 10'd981; b_exp1 = 10'd824; b_exp2 = 10'd39; b_exp3 = 10'd43;
a_sign0 = 4'd8; a_sign1 = 4'd13; a_sign2 = 4'd7; a_sign3 = 4'd11;
b_sign0 = 4'd8; b_sign1 = 4'd0; b_sign2 = 4'd4; b_sign3 = 4'd1;
@(posedge clk_i);
a_mant0 = 8'd67; a_mant1 = 8'd145; a_mant2 = 8'd33; a_mant3 = 8'd124;
b_mant0 = 8'd83; b_mant1 = 8'd92; b_mant2 = 8'd114; b_mant3 = 8'd118;
a_exp0 = 10'd76; a_exp1 = 10'd590; a_exp2 = 10'd381; a_exp3 = 10'd654;
b_exp0 = 10'd755; b_exp1 = 10'd939; b_exp2 = 10'd889; b_exp3 = 10'd652;
a_sign0 = 4'd10; a_sign1 = 4'd8; a_sign2 = 4'd2; a_sign3 = 4'd16;
b_sign0 = 4'd13; b_sign1 = 4'd4; b_sign2 = 4'd15; b_sign3 = 4'd4;
@(posedge clk_i);
a_mant0 = 8'd12; a_mant1 = 8'd102; a_mant2 = 8'd174; a_mant3 = 8'd222;
b_mant0 = 8'd8; b_mant1 = 8'd89; b_mant2 = 8'd140; b_mant3 = 8'd122;
a_exp0 = 10'd374; a_exp1 = 10'd197; a_exp2 = 10'd736; a_exp3 = 10'd162;
b_exp0 = 10'd219; b_exp1 = 10'd665; b_exp2 = 10'd164; b_exp3 = 10'd144;
a_sign0 = 4'd8; a_sign1 = 4'd16; a_sign2 = 4'd8; a_sign3 = 4'd3;
b_sign0 = 4'd7; b_sign1 = 4'd11; b_sign2 = 4'd4; b_sign3 = 4'd10;
@(posedge clk_i);
a_mant0 = 8'd163; a_mant1 = 8'd198; a_mant2 = 8'd176; a_mant3 = 8'd50;
b_mant0 = 8'd62; b_mant1 = 8'd113; b_mant2 = 8'd215; b_mant3 = 8'd56;
a_exp0 = 10'd374; a_exp1 = 10'd757; a_exp2 = 10'd673; a_exp3 = 10'd622;
b_exp0 = 10'd75; b_exp1 = 10'd459; b_exp2 = 10'd449; b_exp3 = 10'd617;
a_sign0 = 4'd6; a_sign1 = 4'd10; a_sign2 = 4'd8; a_sign3 = 4'd8;
b_sign0 = 4'd7; b_sign1 = 4'd15; b_sign2 = 4'd10; b_sign3 = 4'd15;
@(posedge clk_i);
a_mant0 = 8'd65; a_mant1 = 8'd99; a_mant2 = 8'd123; a_mant3 = 8'd206;
b_mant0 = 8'd91; b_mant1 = 8'd80; b_mant2 = 8'd234; b_mant3 = 8'd150;
a_exp0 = 10'd406; a_exp1 = 10'd386; a_exp2 = 10'd881; a_exp3 = 10'd512;
b_exp0 = 10'd602; b_exp1 = 10'd903; b_exp2 = 10'd82; b_exp3 = 10'd193;
a_sign0 = 4'd7; a_sign1 = 4'd5; a_sign2 = 4'd4; a_sign3 = 4'd7;
b_sign0 = 4'd9; b_sign1 = 4'd0; b_sign2 = 4'd0; b_sign3 = 4'd9;
@(posedge clk_i);
a_mant0 = 8'd248; a_mant1 = 8'd196; a_mant2 = 8'd250; a_mant3 = 8'd178;
b_mant0 = 8'd138; b_mant1 = 8'd128; b_mant2 = 8'd64; b_mant3 = 8'd31;
a_exp0 = 10'd648; a_exp1 = 10'd546; a_exp2 = 10'd909; a_exp3 = 10'd401;
b_exp0 = 10'd869; b_exp1 = 10'd996; b_exp2 = 10'd420; b_exp3 = 10'd797;
a_sign0 = 4'd8; a_sign1 = 4'd9; a_sign2 = 4'd16; a_sign3 = 4'd3;
b_sign0 = 4'd11; b_sign1 = 4'd10; b_sign2 = 4'd10; b_sign3 = 4'd0;
@(posedge clk_i);
a_mant0 = 8'd55; a_mant1 = 8'd45; a_mant2 = 8'd58; a_mant3 = 8'd215;
b_mant0 = 8'd123; b_mant1 = 8'd244; b_mant2 = 8'd86; b_mant3 = 8'd135;
a_exp0 = 10'd937; a_exp1 = 10'd137; a_exp2 = 10'd344; a_exp3 = 10'd356;
b_exp0 = 10'd156; b_exp1 = 10'd521; b_exp2 = 10'd807; b_exp3 = 10'd40;
a_sign0 = 4'd6; a_sign1 = 4'd7; a_sign2 = 4'd7; a_sign3 = 4'd0;
b_sign0 = 4'd7; b_sign1 = 4'd11; b_sign2 = 4'd9; b_sign3 = 4'd2;
@(posedge clk_i);
a_mant0 = 8'd183; a_mant1 = 8'd98; a_mant2 = 8'd251; a_mant3 = 8'd119;
b_mant0 = 8'd68; b_mant1 = 8'd76; b_mant2 = 8'd49; b_mant3 = 8'd230;
a_exp0 = 10'd821; a_exp1 = 10'd952; a_exp2 = 10'd1015; a_exp3 = 10'd625;
b_exp0 = 10'd897; b_exp1 = 10'd953; b_exp2 = 10'd275; b_exp3 = 10'd966;
a_sign0 = 4'd1; a_sign1 = 4'd0; a_sign2 = 4'd6; a_sign3 = 4'd12;
b_sign0 = 4'd8; b_sign1 = 4'd6; b_sign2 = 4'd16; b_sign3 = 4'd5;
@(posedge clk_i);
shared_exps0 = 8'd171;
shared_exps1 = 8'd125;
rstn = 0;
@(posedge clk_i);
rstn = 1;
a_mant0 = 8'd173; a_mant1 = 8'd182; a_mant2 = 8'd123; a_mant3 = 8'd222;
b_mant0 = 8'd80; b_mant1 = 8'd125; b_mant2 = 8'd113; b_mant3 = 8'd79;
a_exp0 = 10'd722; a_exp1 = 10'd32; a_exp2 = 10'd801; a_exp3 = 10'd867;
b_exp0 = 10'd437; b_exp1 = 10'd299; b_exp2 = 10'd469; b_exp3 = 10'd746;
a_sign0 = 4'd9; a_sign1 = 4'd10; a_sign2 = 4'd4; a_sign3 = 4'd2;
b_sign0 = 4'd10; b_sign1 = 4'd7; b_sign2 = 4'd6; b_sign3 = 4'd4;
@(posedge clk_i);
a_mant0 = 8'd246; a_mant1 = 8'd86; a_mant2 = 8'd217; a_mant3 = 8'd140;
b_mant0 = 8'd205; b_mant1 = 8'd149; b_mant2 = 8'd55; b_mant3 = 8'd186;
a_exp0 = 10'd938; a_exp1 = 10'd592; a_exp2 = 10'd982; a_exp3 = 10'd38;
b_exp0 = 10'd154; b_exp1 = 10'd55; b_exp2 = 10'd738; b_exp3 = 10'd444;
a_sign0 = 4'd16; a_sign1 = 4'd1; a_sign2 = 4'd12; a_sign3 = 4'd14;
b_sign0 = 4'd15; b_sign1 = 4'd12; b_sign2 = 4'd9; b_sign3 = 4'd4;
@(posedge clk_i);
a_mant0 = 8'd23; a_mant1 = 8'd239; a_mant2 = 8'd181; a_mant3 = 8'd203;
b_mant0 = 8'd162; b_mant1 = 8'd24; b_mant2 = 8'd130; b_mant3 = 8'd185;
a_exp0 = 10'd319; a_exp1 = 10'd888; a_exp2 = 10'd410; a_exp3 = 10'd494;
b_exp0 = 10'd529; b_exp1 = 10'd787; b_exp2 = 10'd658; b_exp3 = 10'd765;
a_sign0 = 4'd8; a_sign1 = 4'd1; a_sign2 = 4'd13; a_sign3 = 4'd8;
b_sign0 = 4'd12; b_sign1 = 4'd16; b_sign2 = 4'd11; b_sign3 = 4'd5;
@(posedge clk_i);
a_mant0 = 8'd47; a_mant1 = 8'd182; a_mant2 = 8'd234; a_mant3 = 8'd132;
b_mant0 = 8'd196; b_mant1 = 8'd218; b_mant2 = 8'd242; b_mant3 = 8'd160;
a_exp0 = 10'd71; a_exp1 = 10'd936; a_exp2 = 10'd343; a_exp3 = 10'd536;
b_exp0 = 10'd1006; b_exp1 = 10'd931; b_exp2 = 10'd174; b_exp3 = 10'd791;
a_sign0 = 4'd6; a_sign1 = 4'd5; a_sign2 = 4'd9; a_sign3 = 4'd13;
b_sign0 = 4'd4; b_sign1 = 4'd7; b_sign2 = 4'd11; b_sign3 = 4'd4;
@(posedge clk_i);
a_mant0 = 8'd60; a_mant1 = 8'd190; a_mant2 = 8'd239; a_mant3 = 8'd36;
b_mant0 = 8'd187; b_mant1 = 8'd169; b_mant2 = 8'd235; b_mant3 = 8'd86;
a_exp0 = 10'd8; a_exp1 = 10'd305; a_exp2 = 10'd454; a_exp3 = 10'd973;
b_exp0 = 10'd16; b_exp1 = 10'd32; b_exp2 = 10'd815; b_exp3 = 10'd466;
a_sign0 = 4'd16; a_sign1 = 4'd15; a_sign2 = 4'd6; a_sign3 = 4'd16;
b_sign0 = 4'd4; b_sign1 = 4'd6; b_sign2 = 4'd7; b_sign3 = 4'd13;
@(posedge clk_i);
a_mant0 = 8'd124; a_mant1 = 8'd248; a_mant2 = 8'd220; a_mant3 = 8'd227;
b_mant0 = 8'd36; b_mant1 = 8'd129; b_mant2 = 8'd219; b_mant3 = 8'd163;
a_exp0 = 10'd460; a_exp1 = 10'd697; a_exp2 = 10'd925; a_exp3 = 10'd343;
b_exp0 = 10'd336; b_exp1 = 10'd673; b_exp2 = 10'd534; b_exp3 = 10'd950;
a_sign0 = 4'd13; a_sign1 = 4'd13; a_sign2 = 4'd0; a_sign3 = 4'd4;
b_sign0 = 4'd8; b_sign1 = 4'd15; b_sign2 = 4'd5; b_sign3 = 4'd7;
@(posedge clk_i);
a_mant0 = 8'd22; a_mant1 = 8'd130; a_mant2 = 8'd169; a_mant3 = 8'd232;
b_mant0 = 8'd167; b_mant1 = 8'd182; b_mant2 = 8'd114; b_mant3 = 8'd220;
a_exp0 = 10'd1004; a_exp1 = 10'd688; a_exp2 = 10'd593; a_exp3 = 10'd613;
b_exp0 = 10'd944; b_exp1 = 10'd299; b_exp2 = 10'd111; b_exp3 = 10'd934;
a_sign0 = 4'd9; a_sign1 = 4'd0; a_sign2 = 4'd10; a_sign3 = 4'd8;
b_sign0 = 4'd1; b_sign1 = 4'd10; b_sign2 = 4'd13; b_sign3 = 4'd16;
@(posedge clk_i);
shared_exps0 = 8'd133;
shared_exps1 = 8'd139;
a_mant0 = 8'd251; a_mant1 = 8'd0; a_mant2 = 8'd180; a_mant3 = 8'd89;
b_mant0 = 8'd67; b_mant1 = 8'd95; b_mant2 = 8'd148; b_mant3 = 8'd243;
a_exp0 = 10'd218; a_exp1 = 10'd520; a_exp2 = 10'd955; a_exp3 = 10'd276;
b_exp0 = 10'd256; b_exp1 = 10'd299; b_exp2 = 10'd114; b_exp3 = 10'd962;
a_sign0 = 4'd5; a_sign1 = 4'd0; a_sign2 = 4'd12; a_sign3 = 4'd13;
b_sign0 = 4'd7; b_sign1 = 4'd3; b_sign2 = 4'd5; b_sign3 = 4'd13;
@(posedge clk_i);
a_mant0 = 8'd253; a_mant1 = 8'd184; a_mant2 = 8'd236; a_mant3 = 8'd103;
b_mant0 = 8'd191; b_mant1 = 8'd14; b_mant2 = 8'd117; b_mant3 = 8'd149;
a_exp0 = 10'd224; a_exp1 = 10'd914; a_exp2 = 10'd697; a_exp3 = 10'd122;
b_exp0 = 10'd680; b_exp1 = 10'd29; b_exp2 = 10'd69; b_exp3 = 10'd143;
a_sign0 = 4'd5; a_sign1 = 4'd0; a_sign2 = 4'd6; a_sign3 = 4'd13;
b_sign0 = 4'd5; b_sign1 = 4'd0; b_sign2 = 4'd0; b_sign3 = 4'd1;
@(posedge clk_i);
a_mant0 = 8'd95; a_mant1 = 8'd15; a_mant2 = 8'd82; a_mant3 = 8'd233;
b_mant0 = 8'd196; b_mant1 = 8'd1; b_mant2 = 8'd187; b_mant3 = 8'd251;
a_exp0 = 10'd613; a_exp1 = 10'd244; a_exp2 = 10'd196; a_exp3 = 10'd554;
b_exp0 = 10'd146; b_exp1 = 10'd232; b_exp2 = 10'd363; b_exp3 = 10'd771;
a_sign0 = 4'd6; a_sign1 = 4'd16; a_sign2 = 4'd3; a_sign3 = 4'd11;
b_sign0 = 4'd13; b_sign1 = 4'd14; b_sign2 = 4'd15; b_sign3 = 4'd2;
@(posedge clk_i);
a_mant0 = 8'd42; a_mant1 = 8'd49; a_mant2 = 8'd191; a_mant3 = 8'd33;
b_mant0 = 8'd193; b_mant1 = 8'd138; b_mant2 = 8'd147; b_mant3 = 8'd112;
a_exp0 = 10'd862; a_exp1 = 10'd506; a_exp2 = 10'd733; a_exp3 = 10'd174;
b_exp0 = 10'd409; b_exp1 = 10'd607; b_exp2 = 10'd351; b_exp3 = 10'd627;
a_sign0 = 4'd14; a_sign1 = 4'd4; a_sign2 = 4'd12; a_sign3 = 4'd0;
b_sign0 = 4'd2; b_sign1 = 4'd9; b_sign2 = 4'd7; b_sign3 = 4'd6;
@(posedge clk_i);
a_mant0 = 8'd112; a_mant1 = 8'd221; a_mant2 = 8'd215; a_mant3 = 8'd233;
b_mant0 = 8'd227; b_mant1 = 8'd207; b_mant2 = 8'd83; b_mant3 = 8'd16;
a_exp0 = 10'd208; a_exp1 = 10'd853; a_exp2 = 10'd133; a_exp3 = 10'd868;
b_exp0 = 10'd360; b_exp1 = 10'd645; b_exp2 = 10'd350; b_exp3 = 10'd217;
a_sign0 = 4'd6; a_sign1 = 4'd15; a_sign2 = 4'd16; a_sign3 = 4'd16;
b_sign0 = 4'd15; b_sign1 = 4'd15; b_sign2 = 4'd10; b_sign3 = 4'd6;
@(posedge clk_i);
a_mant0 = 8'd236; a_mant1 = 8'd86; a_mant2 = 8'd141; a_mant3 = 8'd108;
b_mant0 = 8'd150; b_mant1 = 8'd24; b_mant2 = 8'd58; b_mant3 = 8'd169;
a_exp0 = 10'd939; a_exp1 = 10'd379; a_exp2 = 10'd225; a_exp3 = 10'd537;
b_exp0 = 10'd106; b_exp1 = 10'd264; b_exp2 = 10'd11; b_exp3 = 10'd766;
a_sign0 = 4'd3; a_sign1 = 4'd12; a_sign2 = 4'd15; a_sign3 = 4'd11;
b_sign0 = 4'd6; b_sign1 = 4'd1; b_sign2 = 4'd7; b_sign3 = 4'd1;
@(posedge clk_i);
a_mant0 = 8'd190; a_mant1 = 8'd69; a_mant2 = 8'd10; a_mant3 = 8'd69;
b_mant0 = 8'd162; b_mant1 = 8'd109; b_mant2 = 8'd215; b_mant3 = 8'd15;
a_exp0 = 10'd746; a_exp1 = 10'd664; a_exp2 = 10'd17; a_exp3 = 10'd619;
b_exp0 = 10'd338; b_exp1 = 10'd960; b_exp2 = 10'd217; b_exp3 = 10'd790;
a_sign0 = 4'd3; a_sign1 = 4'd12; a_sign2 = 4'd1; a_sign3 = 4'd15;
b_sign0 = 4'd1; b_sign1 = 4'd14; b_sign2 = 4'd7; b_sign3 = 4'd16;
@(posedge clk_i);
a_mant0 = 8'd129; a_mant1 = 8'd93; a_mant2 = 8'd28; a_mant3 = 8'd96;
b_mant0 = 8'd130; b_mant1 = 8'd100; b_mant2 = 8'd114; b_mant3 = 8'd121;
a_exp0 = 10'd69; a_exp1 = 10'd893; a_exp2 = 10'd195; a_exp3 = 10'd16;
b_exp0 = 10'd895; b_exp1 = 10'd1010; b_exp2 = 10'd396; b_exp3 = 10'd747;
a_sign0 = 4'd4; a_sign1 = 4'd5; a_sign2 = 4'd10; a_sign3 = 4'd8;
b_sign0 = 4'd5; b_sign1 = 4'd3; b_sign2 = 4'd12; b_sign3 = 4'd7;
@(posedge clk_i);
shared_exps0 = 8'd134;
shared_exps1 = 8'd127;
a_mant0 = 8'd46; a_mant1 = 8'd240; a_mant2 = 8'd238; a_mant3 = 8'd211;
b_mant0 = 8'd137; b_mant1 = 8'd147; b_mant2 = 8'd134; b_mant3 = 8'd190;
a_exp0 = 10'd884; a_exp1 = 10'd981; a_exp2 = 10'd802; a_exp3 = 10'd886;
b_exp0 = 10'd885; b_exp1 = 10'd700; b_exp2 = 10'd534; b_exp3 = 10'd760;
a_sign0 = 4'd4; a_sign1 = 4'd16; a_sign2 = 4'd6; a_sign3 = 4'd3;
b_sign0 = 4'd10; b_sign1 = 4'd12; b_sign2 = 4'd7; b_sign3 = 4'd10;
@(posedge clk_i);
a_mant0 = 8'd147; a_mant1 = 8'd132; a_mant2 = 8'd96; a_mant3 = 8'd78;
b_mant0 = 8'd118; b_mant1 = 8'd159; b_mant2 = 8'd184; b_mant3 = 8'd4;
a_exp0 = 10'd692; a_exp1 = 10'd126; a_exp2 = 10'd552; a_exp3 = 10'd754;
b_exp0 = 10'd528; b_exp1 = 10'd262; b_exp2 = 10'd902; b_exp3 = 10'd577;
a_sign0 = 4'd15; a_sign1 = 4'd6; a_sign2 = 4'd16; a_sign3 = 4'd4;
b_sign0 = 4'd6; b_sign1 = 4'd1; b_sign2 = 4'd8; b_sign3 = 4'd12;
@(posedge clk_i);
a_mant0 = 8'd160; a_mant1 = 8'd171; a_mant2 = 8'd96; a_mant3 = 8'd188;
b_mant0 = 8'd159; b_mant1 = 8'd204; b_mant2 = 8'd236; b_mant3 = 8'd221;
a_exp0 = 10'd78; a_exp1 = 10'd887; a_exp2 = 10'd29; a_exp3 = 10'd773;
b_exp0 = 10'd258; b_exp1 = 10'd882; b_exp2 = 10'd253; b_exp3 = 10'd512;
a_sign0 = 4'd12; a_sign1 = 4'd0; a_sign2 = 4'd10; a_sign3 = 4'd8;
b_sign0 = 4'd4; b_sign1 = 4'd4; b_sign2 = 4'd5; b_sign3 = 4'd14;
@(posedge clk_i);
a_mant0 = 8'd152; a_mant1 = 8'd187; a_mant2 = 8'd11; a_mant3 = 8'd76;
b_mant0 = 8'd126; b_mant1 = 8'd36; b_mant2 = 8'd203; b_mant3 = 8'd5;
a_exp0 = 10'd264; a_exp1 = 10'd791; a_exp2 = 10'd534; a_exp3 = 10'd929;
b_exp0 = 10'd932; b_exp1 = 10'd520; b_exp2 = 10'd191; b_exp3 = 10'd543;
a_sign0 = 4'd10; a_sign1 = 4'd4; a_sign2 = 4'd5; a_sign3 = 4'd16;
b_sign0 = 4'd16; b_sign1 = 4'd2; b_sign2 = 4'd5; b_sign3 = 4'd1;
@(posedge clk_i);
a_mant0 = 8'd100; a_mant1 = 8'd222; a_mant2 = 8'd24; a_mant3 = 8'd200;
b_mant0 = 8'd53; b_mant1 = 8'd224; b_mant2 = 8'd151; b_mant3 = 8'd191;
a_exp0 = 10'd729; a_exp1 = 10'd170; a_exp2 = 10'd832; a_exp3 = 10'd292;
b_exp0 = 10'd15; b_exp1 = 10'd291; b_exp2 = 10'd60; b_exp3 = 10'd234;
a_sign0 = 4'd9; a_sign1 = 4'd2; a_sign2 = 4'd14; a_sign3 = 4'd1;
b_sign0 = 4'd9; b_sign1 = 4'd6; b_sign2 = 4'd15; b_sign3 = 4'd16;
@(posedge clk_i);
a_mant0 = 8'd213; a_mant1 = 8'd138; a_mant2 = 8'd90; a_mant3 = 8'd189;
b_mant0 = 8'd159; b_mant1 = 8'd214; b_mant2 = 8'd90; b_mant3 = 8'd255;
a_exp0 = 10'd72; a_exp1 = 10'd447; a_exp2 = 10'd518; a_exp3 = 10'd474;
b_exp0 = 10'd361; b_exp1 = 10'd455; b_exp2 = 10'd429; b_exp3 = 10'd524;
a_sign0 = 4'd2; a_sign1 = 4'd16; a_sign2 = 4'd2; a_sign3 = 4'd14;
b_sign0 = 4'd16; b_sign1 = 4'd1; b_sign2 = 4'd13; b_sign3 = 4'd13;
@(posedge clk_i);
a_mant0 = 8'd200; a_mant1 = 8'd156; a_mant2 = 8'd86; a_mant3 = 8'd150;
b_mant0 = 8'd128; b_mant1 = 8'd85; b_mant2 = 8'd50; b_mant3 = 8'd157;
a_exp0 = 10'd261; a_exp1 = 10'd954; a_exp2 = 10'd649; a_exp3 = 10'd690;
b_exp0 = 10'd693; b_exp1 = 10'd735; b_exp2 = 10'd753; b_exp3 = 10'd123;
a_sign0 = 4'd11; a_sign1 = 4'd11; a_sign2 = 4'd12; a_sign3 = 4'd5;
b_sign0 = 4'd12; b_sign1 = 4'd4; b_sign2 = 4'd1; b_sign3 = 4'd5;
@(posedge clk_i);
a_mant0 = 8'd172; a_mant1 = 8'd112; a_mant2 = 8'd141; a_mant3 = 8'd71;
b_mant0 = 8'd144; b_mant1 = 8'd6; b_mant2 = 8'd166; b_mant3 = 8'd142;
a_exp0 = 10'd326; a_exp1 = 10'd122; a_exp2 = 10'd499; a_exp3 = 10'd860;
b_exp0 = 10'd88; b_exp1 = 10'd106; b_exp2 = 10'd556; b_exp3 = 10'd354;
a_sign0 = 4'd4; a_sign1 = 4'd13; a_sign2 = 4'd6; a_sign3 = 4'd11;
b_sign0 = 4'd1; b_sign1 = 4'd4; b_sign2 = 4'd4; b_sign3 = 4'd13;
@(posedge clk_i);
shared_exps0 = 8'd105;
shared_exps1 = 8'd138;
a_mant0 = 8'd113; a_mant1 = 8'd179; a_mant2 = 8'd254; a_mant3 = 8'd93;
b_mant0 = 8'd173; b_mant1 = 8'd206; b_mant2 = 8'd113; b_mant3 = 8'd96;
a_exp0 = 10'd323; a_exp1 = 10'd843; a_exp2 = 10'd306; a_exp3 = 10'd435;
b_exp0 = 10'd736; b_exp1 = 10'd714; b_exp2 = 10'd467; b_exp3 = 10'd263;
a_sign0 = 4'd5; a_sign1 = 4'd7; a_sign2 = 4'd8; a_sign3 = 4'd5;
b_sign0 = 4'd7; b_sign1 = 4'd14; b_sign2 = 4'd8; b_sign3 = 4'd11;
@(posedge clk_i);
a_mant0 = 8'd114; a_mant1 = 8'd172; a_mant2 = 8'd201; a_mant3 = 8'd182;
b_mant0 = 8'd94; b_mant1 = 8'd106; b_mant2 = 8'd184; b_mant3 = 8'd64;
a_exp0 = 10'd979; a_exp1 = 10'd24; a_exp2 = 10'd78; a_exp3 = 10'd539;
b_exp0 = 10'd936; b_exp1 = 10'd61; b_exp2 = 10'd421; b_exp3 = 10'd319;
a_sign0 = 4'd11; a_sign1 = 4'd7; a_sign2 = 4'd16; a_sign3 = 4'd4;
b_sign0 = 4'd14; b_sign1 = 4'd3; b_sign2 = 4'd2; b_sign3 = 4'd10;
@(posedge clk_i);
a_mant0 = 8'd203; a_mant1 = 8'd114; a_mant2 = 8'd127; a_mant3 = 8'd168;
b_mant0 = 8'd71; b_mant1 = 8'd146; b_mant2 = 8'd189; b_mant3 = 8'd61;
a_exp0 = 10'd716; a_exp1 = 10'd490; a_exp2 = 10'd143; a_exp3 = 10'd752;
b_exp0 = 10'd268; b_exp1 = 10'd331; b_exp2 = 10'd463; b_exp3 = 10'd554;
a_sign0 = 4'd1; a_sign1 = 4'd12; a_sign2 = 4'd13; a_sign3 = 4'd15;
b_sign0 = 4'd7; b_sign1 = 4'd2; b_sign2 = 4'd0; b_sign3 = 4'd3;
@(posedge clk_i);
a_mant0 = 8'd191; a_mant1 = 8'd140; a_mant2 = 8'd111; a_mant3 = 8'd72;
b_mant0 = 8'd214; b_mant1 = 8'd44; b_mant2 = 8'd87; b_mant3 = 8'd53;
a_exp0 = 10'd429; a_exp1 = 10'd726; a_exp2 = 10'd144; a_exp3 = 10'd188;
b_exp0 = 10'd749; b_exp1 = 10'd885; b_exp2 = 10'd128; b_exp3 = 10'd116;
a_sign0 = 4'd14; a_sign1 = 4'd15; a_sign2 = 4'd12; a_sign3 = 4'd9;
b_sign0 = 4'd3; b_sign1 = 4'd11; b_sign2 = 4'd9; b_sign3 = 4'd3;
@(posedge clk_i);
a_mant0 = 8'd87; a_mant1 = 8'd17; a_mant2 = 8'd8; a_mant3 = 8'd133;
b_mant0 = 8'd118; b_mant1 = 8'd83; b_mant2 = 8'd141; b_mant3 = 8'd243;
a_exp0 = 10'd836; a_exp1 = 10'd328; a_exp2 = 10'd902; a_exp3 = 10'd162;
b_exp0 = 10'd456; b_exp1 = 10'd242; b_exp2 = 10'd330; b_exp3 = 10'd114;
a_sign0 = 4'd5; a_sign1 = 4'd12; a_sign2 = 4'd3; a_sign3 = 4'd6;
b_sign0 = 4'd2; b_sign1 = 4'd4; b_sign2 = 4'd15; b_sign3 = 4'd0;
@(posedge clk_i);
a_mant0 = 8'd224; a_mant1 = 8'd95; a_mant2 = 8'd177; a_mant3 = 8'd31;
b_mant0 = 8'd206; b_mant1 = 8'd106; b_mant2 = 8'd197; b_mant3 = 8'd72;
a_exp0 = 10'd148; a_exp1 = 10'd233; a_exp2 = 10'd964; a_exp3 = 10'd881;
b_exp0 = 10'd852; b_exp1 = 10'd570; b_exp2 = 10'd491; b_exp3 = 10'd583;
a_sign0 = 4'd14; a_sign1 = 4'd0; a_sign2 = 4'd1; a_sign3 = 4'd7;
b_sign0 = 4'd7; b_sign1 = 4'd16; b_sign2 = 4'd4; b_sign3 = 4'd1;
@(posedge clk_i);
a_mant0 = 8'd78; a_mant1 = 8'd83; a_mant2 = 8'd131; a_mant3 = 8'd193;
b_mant0 = 8'd103; b_mant1 = 8'd172; b_mant2 = 8'd40; b_mant3 = 8'd156;
a_exp0 = 10'd1014; a_exp1 = 10'd333; a_exp2 = 10'd974; a_exp3 = 10'd0;
b_exp0 = 10'd168; b_exp1 = 10'd300; b_exp2 = 10'd675; b_exp3 = 10'd470;
a_sign0 = 4'd8; a_sign1 = 4'd13; a_sign2 = 4'd14; a_sign3 = 4'd10;
b_sign0 = 4'd11; b_sign1 = 4'd0; b_sign2 = 4'd5; b_sign3 = 4'd16;
@(posedge clk_i);
a_mant0 = 8'd53; a_mant1 = 8'd229; a_mant2 = 8'd110; a_mant3 = 8'd111;
b_mant0 = 8'd103; b_mant1 = 8'd214; b_mant2 = 8'd142; b_mant3 = 8'd126;
a_exp0 = 10'd33; a_exp1 = 10'd884; a_exp2 = 10'd922; a_exp3 = 10'd711;
b_exp0 = 10'd393; b_exp1 = 10'd153; b_exp2 = 10'd852; b_exp3 = 10'd402;
a_sign0 = 4'd13; a_sign1 = 4'd16; a_sign2 = 4'd11; a_sign3 = 4'd3;
b_sign0 = 4'd5; b_sign1 = 4'd10; b_sign2 = 4'd16; b_sign3 = 4'd6;
@(posedge clk_i);
shared_exps0 = 8'd145;
shared_exps1 = 8'd103;
rstn = 0;
@(posedge clk_i);
rstn = 1;
a_mant0 = 8'd161; a_mant1 = 8'd140; a_mant2 = 8'd151; a_mant3 = 8'd176;
b_mant0 = 8'd161; b_mant1 = 8'd194; b_mant2 = 8'd29; b_mant3 = 8'd200;
a_exp0 = 10'd352; a_exp1 = 10'd439; a_exp2 = 10'd97; a_exp3 = 10'd364;
b_exp0 = 10'd466; b_exp1 = 10'd22; b_exp2 = 10'd388; b_exp3 = 10'd749;
a_sign0 = 4'd14; a_sign1 = 4'd6; a_sign2 = 4'd13; a_sign3 = 4'd10;
b_sign0 = 4'd16; b_sign1 = 4'd8; b_sign2 = 4'd9; b_sign3 = 4'd0;
@(posedge clk_i);
a_mant0 = 8'd28; a_mant1 = 8'd80; a_mant2 = 8'd93; a_mant3 = 8'd34;
b_mant0 = 8'd102; b_mant1 = 8'd97; b_mant2 = 8'd176; b_mant3 = 8'd248;
a_exp0 = 10'd605; a_exp1 = 10'd170; a_exp2 = 10'd919; a_exp3 = 10'd528;
b_exp0 = 10'd574; b_exp1 = 10'd273; b_exp2 = 10'd692; b_exp3 = 10'd625;
a_sign0 = 4'd3; a_sign1 = 4'd8; a_sign2 = 4'd9; a_sign3 = 4'd4;
b_sign0 = 4'd6; b_sign1 = 4'd0; b_sign2 = 4'd15; b_sign3 = 4'd13;
@(posedge clk_i);
a_mant0 = 8'd66; a_mant1 = 8'd26; a_mant2 = 8'd181; a_mant3 = 8'd39;
b_mant0 = 8'd219; b_mant1 = 8'd85; b_mant2 = 8'd246; b_mant3 = 8'd221;
a_exp0 = 10'd138; a_exp1 = 10'd80; a_exp2 = 10'd506; a_exp3 = 10'd197;
b_exp0 = 10'd848; b_exp1 = 10'd504; b_exp2 = 10'd865; b_exp3 = 10'd326;
a_sign0 = 4'd11; a_sign1 = 4'd6; a_sign2 = 4'd5; a_sign3 = 4'd11;
b_sign0 = 4'd9; b_sign1 = 4'd10; b_sign2 = 4'd3; b_sign3 = 4'd6;
@(posedge clk_i);
a_mant0 = 8'd240; a_mant1 = 8'd224; a_mant2 = 8'd246; a_mant3 = 8'd68;
b_mant0 = 8'd95; b_mant1 = 8'd43; b_mant2 = 8'd8; b_mant3 = 8'd38;
a_exp0 = 10'd626; a_exp1 = 10'd669; a_exp2 = 10'd42; a_exp3 = 10'd872;
b_exp0 = 10'd823; b_exp1 = 10'd927; b_exp2 = 10'd1012; b_exp3 = 10'd21;
a_sign0 = 4'd14; a_sign1 = 4'd1; a_sign2 = 4'd8; a_sign3 = 4'd5;
b_sign0 = 4'd2; b_sign1 = 4'd15; b_sign2 = 4'd11; b_sign3 = 4'd4;
@(posedge clk_i);
a_mant0 = 8'd117; a_mant1 = 8'd234; a_mant2 = 8'd36; a_mant3 = 8'd135;
b_mant0 = 8'd209; b_mant1 = 8'd108; b_mant2 = 8'd53; b_mant3 = 8'd161;
a_exp0 = 10'd200; a_exp1 = 10'd899; a_exp2 = 10'd254; a_exp3 = 10'd894;
b_exp0 = 10'd576; b_exp1 = 10'd469; b_exp2 = 10'd864; b_exp3 = 10'd550;
a_sign0 = 4'd13; a_sign1 = 4'd6; a_sign2 = 4'd8; a_sign3 = 4'd10;
b_sign0 = 4'd13; b_sign1 = 4'd16; b_sign2 = 4'd11; b_sign3 = 4'd11;
@(posedge clk_i);
a_mant0 = 8'd123; a_mant1 = 8'd249; a_mant2 = 8'd250; a_mant3 = 8'd165;
b_mant0 = 8'd82; b_mant1 = 8'd95; b_mant2 = 8'd142; b_mant3 = 8'd245;
a_exp0 = 10'd804; a_exp1 = 10'd651; a_exp2 = 10'd878; a_exp3 = 10'd225;
b_exp0 = 10'd819; b_exp1 = 10'd837; b_exp2 = 10'd577; b_exp3 = 10'd840;
a_sign0 = 4'd8; a_sign1 = 4'd10; a_sign2 = 4'd2; a_sign3 = 4'd16;
b_sign0 = 4'd0; b_sign1 = 4'd15; b_sign2 = 4'd2; b_sign3 = 4'd8;
@(posedge clk_i);
a_mant0 = 8'd22; a_mant1 = 8'd114; a_mant2 = 8'd212; a_mant3 = 8'd148;
b_mant0 = 8'd221; b_mant1 = 8'd176; b_mant2 = 8'd115; b_mant3 = 8'd21;
a_exp0 = 10'd704; a_exp1 = 10'd793; a_exp2 = 10'd363; a_exp3 = 10'd686;
b_exp0 = 10'd27; b_exp1 = 10'd181; b_exp2 = 10'd868; b_exp3 = 10'd534;
a_sign0 = 4'd0; a_sign1 = 4'd4; a_sign2 = 4'd16; a_sign3 = 4'd5;
b_sign0 = 4'd2; b_sign1 = 4'd16; b_sign2 = 4'd13; b_sign3 = 4'd16;
@(posedge clk_i);
shared_exps0 = 8'd153;
shared_exps1 = 8'd147;
a_mant0 = 8'd27; a_mant1 = 8'd24; a_mant2 = 8'd143; a_mant3 = 8'd224;
b_mant0 = 8'd83; b_mant1 = 8'd100; b_mant2 = 8'd34; b_mant3 = 8'd50;
a_exp0 = 10'd968; a_exp1 = 10'd548; a_exp2 = 10'd2; a_exp3 = 10'd305;
b_exp0 = 10'd230; b_exp1 = 10'd727; b_exp2 = 10'd847; b_exp3 = 10'd216;
a_sign0 = 4'd0; a_sign1 = 4'd16; a_sign2 = 4'd5; a_sign3 = 4'd13;
b_sign0 = 4'd15; b_sign1 = 4'd13; b_sign2 = 4'd15; b_sign3 = 4'd10;
@(posedge clk_i);
a_mant0 = 8'd159; a_mant1 = 8'd92; a_mant2 = 8'd112; a_mant3 = 8'd189;
b_mant0 = 8'd164; b_mant1 = 8'd107; b_mant2 = 8'd50; b_mant3 = 8'd179;
a_exp0 = 10'd711; a_exp1 = 10'd781; a_exp2 = 10'd212; a_exp3 = 10'd860;
b_exp0 = 10'd445; b_exp1 = 10'd991; b_exp2 = 10'd925; b_exp3 = 10'd749;
a_sign0 = 4'd7; a_sign1 = 4'd13; a_sign2 = 4'd10; a_sign3 = 4'd15;
b_sign0 = 4'd0; b_sign1 = 4'd2; b_sign2 = 4'd2; b_sign3 = 4'd12;
@(posedge clk_i);
a_mant0 = 8'd198; a_mant1 = 8'd65; a_mant2 = 8'd127; a_mant3 = 8'd183;
b_mant0 = 8'd102; b_mant1 = 8'd155; b_mant2 = 8'd153; b_mant3 = 8'd107;
a_exp0 = 10'd243; a_exp1 = 10'd167; a_exp2 = 10'd760; a_exp3 = 10'd34;
b_exp0 = 10'd375; b_exp1 = 10'd152; b_exp2 = 10'd839; b_exp3 = 10'd184;
a_sign0 = 4'd14; a_sign1 = 4'd2; a_sign2 = 4'd9; a_sign3 = 4'd7;
b_sign0 = 4'd6; b_sign1 = 4'd14; b_sign2 = 4'd16; b_sign3 = 4'd11;
@(posedge clk_i);
a_mant0 = 8'd230; a_mant1 = 8'd220; a_mant2 = 8'd215; a_mant3 = 8'd108;
b_mant0 = 8'd135; b_mant1 = 8'd42; b_mant2 = 8'd218; b_mant3 = 8'd15;
a_exp0 = 10'd467; a_exp1 = 10'd203; a_exp2 = 10'd809; a_exp3 = 10'd210;
b_exp0 = 10'd190; b_exp1 = 10'd688; b_exp2 = 10'd66; b_exp3 = 10'd523;
a_sign0 = 4'd10; a_sign1 = 4'd15; a_sign2 = 4'd8; a_sign3 = 4'd4;
b_sign0 = 4'd10; b_sign1 = 4'd5; b_sign2 = 4'd15; b_sign3 = 4'd1;
@(posedge clk_i);
a_mant0 = 8'd70; a_mant1 = 8'd216; a_mant2 = 8'd52; a_mant3 = 8'd102;
b_mant0 = 8'd98; b_mant1 = 8'd171; b_mant2 = 8'd149; b_mant3 = 8'd236;
a_exp0 = 10'd38; a_exp1 = 10'd75; a_exp2 = 10'd309; a_exp3 = 10'd194;
b_exp0 = 10'd897; b_exp1 = 10'd412; b_exp2 = 10'd399; b_exp3 = 10'd63;
a_sign0 = 4'd1; a_sign1 = 4'd12; a_sign2 = 4'd4; a_sign3 = 4'd9;
b_sign0 = 4'd5; b_sign1 = 4'd0; b_sign2 = 4'd14; b_sign3 = 4'd14;
@(posedge clk_i);
a_mant0 = 8'd251; a_mant1 = 8'd242; a_mant2 = 8'd120; a_mant3 = 8'd237;
b_mant0 = 8'd228; b_mant1 = 8'd62; b_mant2 = 8'd160; b_mant3 = 8'd64;
a_exp0 = 10'd453; a_exp1 = 10'd466; a_exp2 = 10'd968; a_exp3 = 10'd631;
b_exp0 = 10'd666; b_exp1 = 10'd213; b_exp2 = 10'd46; b_exp3 = 10'd119;
a_sign0 = 4'd4; a_sign1 = 4'd12; a_sign2 = 4'd6; a_sign3 = 4'd2;
b_sign0 = 4'd8; b_sign1 = 4'd3; b_sign2 = 4'd11; b_sign3 = 4'd3;
@(posedge clk_i);
a_mant0 = 8'd108; a_mant1 = 8'd246; a_mant2 = 8'd35; a_mant3 = 8'd143;
b_mant0 = 8'd209; b_mant1 = 8'd30; b_mant2 = 8'd41; b_mant3 = 8'd74;
a_exp0 = 10'd306; a_exp1 = 10'd36; a_exp2 = 10'd784; a_exp3 = 10'd116;
b_exp0 = 10'd334; b_exp1 = 10'd250; b_exp2 = 10'd932; b_exp3 = 10'd30;
a_sign0 = 4'd11; a_sign1 = 4'd5; a_sign2 = 4'd14; a_sign3 = 4'd3;
b_sign0 = 4'd13; b_sign1 = 4'd2; b_sign2 = 4'd6; b_sign3 = 4'd6;
@(posedge clk_i);
a_mant0 = 8'd249; a_mant1 = 8'd130; a_mant2 = 8'd144; a_mant3 = 8'd243;
b_mant0 = 8'd177; b_mant1 = 8'd59; b_mant2 = 8'd239; b_mant3 = 8'd175;
a_exp0 = 10'd148; a_exp1 = 10'd363; a_exp2 = 10'd590; a_exp3 = 10'd840;
b_exp0 = 10'd518; b_exp1 = 10'd999; b_exp2 = 10'd323; b_exp3 = 10'd197;
a_sign0 = 4'd13; a_sign1 = 4'd6; a_sign2 = 4'd16; a_sign3 = 4'd16;
b_sign0 = 4'd9; b_sign1 = 4'd3; b_sign2 = 4'd1; b_sign3 = 4'd6;
@(posedge clk_i);
shared_exps0 = 8'd137;
shared_exps1 = 8'd136;
a_mant0 = 8'd219; a_mant1 = 8'd206; a_mant2 = 8'd64; a_mant3 = 8'd15;
b_mant0 = 8'd0; b_mant1 = 8'd231; b_mant2 = 8'd55; b_mant3 = 8'd44;
a_exp0 = 10'd5; a_exp1 = 10'd908; a_exp2 = 10'd853; a_exp3 = 10'd59;
b_exp0 = 10'd290; b_exp1 = 10'd945; b_exp2 = 10'd755; b_exp3 = 10'd956;
a_sign0 = 4'd3; a_sign1 = 4'd1; a_sign2 = 4'd3; a_sign3 = 4'd8;
b_sign0 = 4'd1; b_sign1 = 4'd4; b_sign2 = 4'd7; b_sign3 = 4'd7;
@(posedge clk_i);
a_mant0 = 8'd201; a_mant1 = 8'd144; a_mant2 = 8'd230; a_mant3 = 8'd157;
b_mant0 = 8'd254; b_mant1 = 8'd173; b_mant2 = 8'd251; b_mant3 = 8'd248;
a_exp0 = 10'd158; a_exp1 = 10'd142; a_exp2 = 10'd197; a_exp3 = 10'd501;
b_exp0 = 10'd587; b_exp1 = 10'd447; b_exp2 = 10'd505; b_exp3 = 10'd542;
a_sign0 = 4'd2; a_sign1 = 4'd5; a_sign2 = 4'd2; a_sign3 = 4'd16;
b_sign0 = 4'd16; b_sign1 = 4'd15; b_sign2 = 4'd5; b_sign3 = 4'd10;
@(posedge clk_i);
a_mant0 = 8'd207; a_mant1 = 8'd223; a_mant2 = 8'd194; a_mant3 = 8'd196;
b_mant0 = 8'd16; b_mant1 = 8'd192; b_mant2 = 8'd199; b_mant3 = 8'd195;
a_exp0 = 10'd492; a_exp1 = 10'd791; a_exp2 = 10'd704; a_exp3 = 10'd929;
b_exp0 = 10'd1019; b_exp1 = 10'd553; b_exp2 = 10'd776; b_exp3 = 10'd888;
a_sign0 = 4'd16; a_sign1 = 4'd7; a_sign2 = 4'd12; a_sign3 = 4'd7;
b_sign0 = 4'd8; b_sign1 = 4'd10; b_sign2 = 4'd2; b_sign3 = 4'd6;
@(posedge clk_i);
a_mant0 = 8'd21; a_mant1 = 8'd26; a_mant2 = 8'd237; a_mant3 = 8'd91;
b_mant0 = 8'd24; b_mant1 = 8'd60; b_mant2 = 8'd74; b_mant3 = 8'd117;
a_exp0 = 10'd263; a_exp1 = 10'd593; a_exp2 = 10'd129; a_exp3 = 10'd384;
b_exp0 = 10'd1016; b_exp1 = 10'd636; b_exp2 = 10'd799; b_exp3 = 10'd731;
a_sign0 = 4'd12; a_sign1 = 4'd7; a_sign2 = 4'd15; a_sign3 = 4'd10;
b_sign0 = 4'd8; b_sign1 = 4'd14; b_sign2 = 4'd6; b_sign3 = 4'd7;
@(posedge clk_i);
a_mant0 = 8'd0; a_mant1 = 8'd47; a_mant2 = 8'd11; a_mant3 = 8'd106;
b_mant0 = 8'd212; b_mant1 = 8'd21; b_mant2 = 8'd50; b_mant3 = 8'd195;
a_exp0 = 10'd144; a_exp1 = 10'd592; a_exp2 = 10'd666; a_exp3 = 10'd611;
b_exp0 = 10'd66; b_exp1 = 10'd803; b_exp2 = 10'd850; b_exp3 = 10'd430;
a_sign0 = 4'd8; a_sign1 = 4'd2; a_sign2 = 4'd7; a_sign3 = 4'd10;
b_sign0 = 4'd13; b_sign1 = 4'd15; b_sign2 = 4'd10; b_sign3 = 4'd0;
@(posedge clk_i);
a_mant0 = 8'd8; a_mant1 = 8'd150; a_mant2 = 8'd74; a_mant3 = 8'd180;
b_mant0 = 8'd222; b_mant1 = 8'd98; b_mant2 = 8'd33; b_mant3 = 8'd229;
a_exp0 = 10'd759; a_exp1 = 10'd596; a_exp2 = 10'd434; a_exp3 = 10'd674;
b_exp0 = 10'd529; b_exp1 = 10'd569; b_exp2 = 10'd381; b_exp3 = 10'd188;
a_sign0 = 4'd16; a_sign1 = 4'd13; a_sign2 = 4'd3; a_sign3 = 4'd15;
b_sign0 = 4'd2; b_sign1 = 4'd7; b_sign2 = 4'd13; b_sign3 = 4'd5;
@(posedge clk_i);
a_mant0 = 8'd207; a_mant1 = 8'd29; a_mant2 = 8'd120; a_mant3 = 8'd97;
b_mant0 = 8'd70; b_mant1 = 8'd12; b_mant2 = 8'd134; b_mant3 = 8'd31;
a_exp0 = 10'd586; a_exp1 = 10'd646; a_exp2 = 10'd621; a_exp3 = 10'd586;
b_exp0 = 10'd439; b_exp1 = 10'd614; b_exp2 = 10'd564; b_exp3 = 10'd222;
a_sign0 = 4'd0; a_sign1 = 4'd12; a_sign2 = 4'd10; a_sign3 = 4'd5;
b_sign0 = 4'd6; b_sign1 = 4'd8; b_sign2 = 4'd2; b_sign3 = 4'd1;
@(posedge clk_i);
a_mant0 = 8'd78; a_mant1 = 8'd121; a_mant2 = 8'd17; a_mant3 = 8'd75;
b_mant0 = 8'd219; b_mant1 = 8'd178; b_mant2 = 8'd236; b_mant3 = 8'd231;
a_exp0 = 10'd915; a_exp1 = 10'd888; a_exp2 = 10'd677; a_exp3 = 10'd811;
b_exp0 = 10'd149; b_exp1 = 10'd560; b_exp2 = 10'd710; b_exp3 = 10'd380;
a_sign0 = 4'd7; a_sign1 = 4'd13; a_sign2 = 4'd2; a_sign3 = 4'd5;
b_sign0 = 4'd7; b_sign1 = 4'd5; b_sign2 = 4'd8; b_sign3 = 4'd13;
@(posedge clk_i);
shared_exps0 = 8'd134;
shared_exps1 = 8'd137;
a_mant0 = 8'd82; a_mant1 = 8'd86; a_mant2 = 8'd200; a_mant3 = 8'd190;
b_mant0 = 8'd41; b_mant1 = 8'd168; b_mant2 = 8'd204; b_mant3 = 8'd188;
a_exp0 = 10'd443; a_exp1 = 10'd929; a_exp2 = 10'd236; a_exp3 = 10'd175;
b_exp0 = 10'd714; b_exp1 = 10'd945; b_exp2 = 10'd0; b_exp3 = 10'd599;
a_sign0 = 4'd2; a_sign1 = 4'd5; a_sign2 = 4'd14; a_sign3 = 4'd10;
b_sign0 = 4'd7; b_sign1 = 4'd6; b_sign2 = 4'd3; b_sign3 = 4'd7;
@(posedge clk_i);
a_mant0 = 8'd65; a_mant1 = 8'd213; a_mant2 = 8'd2; a_mant3 = 8'd154;
b_mant0 = 8'd135; b_mant1 = 8'd56; b_mant2 = 8'd173; b_mant3 = 8'd54;
a_exp0 = 10'd94; a_exp1 = 10'd309; a_exp2 = 10'd541; a_exp3 = 10'd934;
b_exp0 = 10'd839; b_exp1 = 10'd639; b_exp2 = 10'd808; b_exp3 = 10'd625;
a_sign0 = 4'd7; a_sign1 = 4'd12; a_sign2 = 4'd7; a_sign3 = 4'd3;
b_sign0 = 4'd14; b_sign1 = 4'd9; b_sign2 = 4'd14; b_sign3 = 4'd13;
@(posedge clk_i);
a_mant0 = 8'd231; a_mant1 = 8'd72; a_mant2 = 8'd159; a_mant3 = 8'd126;
b_mant0 = 8'd10; b_mant1 = 8'd99; b_mant2 = 8'd148; b_mant3 = 8'd213;
a_exp0 = 10'd947; a_exp1 = 10'd905; a_exp2 = 10'd623; a_exp3 = 10'd484;
b_exp0 = 10'd748; b_exp1 = 10'd631; b_exp2 = 10'd660; b_exp3 = 10'd939;
a_sign0 = 4'd6; a_sign1 = 4'd4; a_sign2 = 4'd13; a_sign3 = 4'd3;
b_sign0 = 4'd9; b_sign1 = 4'd8; b_sign2 = 4'd14; b_sign3 = 4'd2;
@(posedge clk_i);
a_mant0 = 8'd229; a_mant1 = 8'd7; a_mant2 = 8'd31; a_mant3 = 8'd88;
b_mant0 = 8'd84; b_mant1 = 8'd128; b_mant2 = 8'd151; b_mant3 = 8'd135;
a_exp0 = 10'd541; a_exp1 = 10'd131; a_exp2 = 10'd185; a_exp3 = 10'd555;
b_exp0 = 10'd436; b_exp1 = 10'd209; b_exp2 = 10'd110; b_exp3 = 10'd518;
a_sign0 = 4'd8; a_sign1 = 4'd1; a_sign2 = 4'd7; a_sign3 = 4'd6;
b_sign0 = 4'd8; b_sign1 = 4'd4; b_sign2 = 4'd3; b_sign3 = 4'd13;
@(posedge clk_i);
a_mant0 = 8'd96; a_mant1 = 8'd233; a_mant2 = 8'd195; a_mant3 = 8'd196;
b_mant0 = 8'd89; b_mant1 = 8'd92; b_mant2 = 8'd77; b_mant3 = 8'd250;
a_exp0 = 10'd317; a_exp1 = 10'd179; a_exp2 = 10'd462; a_exp3 = 10'd998;
b_exp0 = 10'd626; b_exp1 = 10'd252; b_exp2 = 10'd184; b_exp3 = 10'd794;
a_sign0 = 4'd14; a_sign1 = 4'd14; a_sign2 = 4'd1; a_sign3 = 4'd14;
b_sign0 = 4'd6; b_sign1 = 4'd7; b_sign2 = 4'd8; b_sign3 = 4'd16;
@(posedge clk_i);
a_mant0 = 8'd27; a_mant1 = 8'd231; a_mant2 = 8'd252; a_mant3 = 8'd27;
b_mant0 = 8'd75; b_mant1 = 8'd137; b_mant2 = 8'd80; b_mant3 = 8'd69;
a_exp0 = 10'd743; a_exp1 = 10'd818; a_exp2 = 10'd514; a_exp3 = 10'd334;
b_exp0 = 10'd194; b_exp1 = 10'd872; b_exp2 = 10'd708; b_exp3 = 10'd390;
a_sign0 = 4'd15; a_sign1 = 4'd2; a_sign2 = 4'd12; a_sign3 = 4'd7;
b_sign0 = 4'd10; b_sign1 = 4'd5; b_sign2 = 4'd3; b_sign3 = 4'd0;
@(posedge clk_i);
a_mant0 = 8'd177; a_mant1 = 8'd153; a_mant2 = 8'd163; a_mant3 = 8'd78;
b_mant0 = 8'd224; b_mant1 = 8'd17; b_mant2 = 8'd120; b_mant3 = 8'd101;
a_exp0 = 10'd945; a_exp1 = 10'd753; a_exp2 = 10'd646; a_exp3 = 10'd313;
b_exp0 = 10'd460; b_exp1 = 10'd714; b_exp2 = 10'd910; b_exp3 = 10'd645;
a_sign0 = 4'd2; a_sign1 = 4'd1; a_sign2 = 4'd10; a_sign3 = 4'd8;
b_sign0 = 4'd5; b_sign1 = 4'd15; b_sign2 = 4'd10; b_sign3 = 4'd6;
@(posedge clk_i);
a_mant0 = 8'd117; a_mant1 = 8'd210; a_mant2 = 8'd49; a_mant3 = 8'd45;
b_mant0 = 8'd119; b_mant1 = 8'd171; b_mant2 = 8'd27; b_mant3 = 8'd255;
a_exp0 = 10'd946; a_exp1 = 10'd560; a_exp2 = 10'd474; a_exp3 = 10'd790;
b_exp0 = 10'd354; b_exp1 = 10'd940; b_exp2 = 10'd44; b_exp3 = 10'd593;
a_sign0 = 4'd1; a_sign1 = 4'd4; a_sign2 = 4'd11; a_sign3 = 4'd16;
b_sign0 = 4'd15; b_sign1 = 4'd9; b_sign2 = 4'd14; b_sign3 = 4'd11;
@(posedge clk_i);
shared_exps0 = 8'd118;
shared_exps1 = 8'd96;
rstn = 0;
@(posedge clk_i);
rstn = 1;
a_mant0 = 8'd73; a_mant1 = 8'd171; a_mant2 = 8'd85; a_mant3 = 8'd162;
b_mant0 = 8'd203; b_mant1 = 8'd226; b_mant2 = 8'd231; b_mant3 = 8'd13;
a_exp0 = 10'd988; a_exp1 = 10'd787; a_exp2 = 10'd770; a_exp3 = 10'd58;
b_exp0 = 10'd453; b_exp1 = 10'd80; b_exp2 = 10'd727; b_exp3 = 10'd1019;
a_sign0 = 4'd2; a_sign1 = 4'd16; a_sign2 = 4'd5; a_sign3 = 4'd11;
b_sign0 = 4'd12; b_sign1 = 4'd7; b_sign2 = 4'd7; b_sign3 = 4'd0;
@(posedge clk_i);
a_mant0 = 8'd97; a_mant1 = 8'd86; a_mant2 = 8'd163; a_mant3 = 8'd253;
b_mant0 = 8'd93; b_mant1 = 8'd244; b_mant2 = 8'd70; b_mant3 = 8'd247;
a_exp0 = 10'd740; a_exp1 = 10'd75; a_exp2 = 10'd752; a_exp3 = 10'd840;
b_exp0 = 10'd941; b_exp1 = 10'd802; b_exp2 = 10'd785; b_exp3 = 10'd915;
a_sign0 = 4'd10; a_sign1 = 4'd3; a_sign2 = 4'd13; a_sign3 = 4'd4;
b_sign0 = 4'd16; b_sign1 = 4'd10; b_sign2 = 4'd13; b_sign3 = 4'd10;
@(posedge clk_i);
a_mant0 = 8'd213; a_mant1 = 8'd180; a_mant2 = 8'd224; a_mant3 = 8'd84;
b_mant0 = 8'd132; b_mant1 = 8'd135; b_mant2 = 8'd173; b_mant3 = 8'd209;
a_exp0 = 10'd449; a_exp1 = 10'd901; a_exp2 = 10'd957; a_exp3 = 10'd586;
b_exp0 = 10'd572; b_exp1 = 10'd551; b_exp2 = 10'd662; b_exp3 = 10'd1017;
a_sign0 = 4'd14; a_sign1 = 4'd3; a_sign2 = 4'd10; a_sign3 = 4'd1;
b_sign0 = 4'd9; b_sign1 = 4'd15; b_sign2 = 4'd1; b_sign3 = 4'd9;
@(posedge clk_i);
a_mant0 = 8'd244; a_mant1 = 8'd68; a_mant2 = 8'd16; a_mant3 = 8'd166;
b_mant0 = 8'd96; b_mant1 = 8'd100; b_mant2 = 8'd57; b_mant3 = 8'd136;
a_exp0 = 10'd848; a_exp1 = 10'd1021; a_exp2 = 10'd1006; a_exp3 = 10'd883;
b_exp0 = 10'd582; b_exp1 = 10'd64; b_exp2 = 10'd879; b_exp3 = 10'd713;
a_sign0 = 4'd0; a_sign1 = 4'd7; a_sign2 = 4'd0; a_sign3 = 4'd2;
b_sign0 = 4'd14; b_sign1 = 4'd13; b_sign2 = 4'd2; b_sign3 = 4'd14;
@(posedge clk_i);
a_mant0 = 8'd229; a_mant1 = 8'd216; a_mant2 = 8'd249; a_mant3 = 8'd219;
b_mant0 = 8'd46; b_mant1 = 8'd2; b_mant2 = 8'd161; b_mant3 = 8'd120;
a_exp0 = 10'd790; a_exp1 = 10'd732; a_exp2 = 10'd587; a_exp3 = 10'd350;
b_exp0 = 10'd837; b_exp1 = 10'd609; b_exp2 = 10'd424; b_exp3 = 10'd730;
a_sign0 = 4'd9; a_sign1 = 4'd6; a_sign2 = 4'd1; a_sign3 = 4'd8;
b_sign0 = 4'd11; b_sign1 = 4'd6; b_sign2 = 4'd9; b_sign3 = 4'd11;
@(posedge clk_i);
a_mant0 = 8'd78; a_mant1 = 8'd118; a_mant2 = 8'd18; a_mant3 = 8'd232;
b_mant0 = 8'd127; b_mant1 = 8'd110; b_mant2 = 8'd219; b_mant3 = 8'd139;
a_exp0 = 10'd759; a_exp1 = 10'd714; a_exp2 = 10'd378; a_exp3 = 10'd991;
b_exp0 = 10'd767; b_exp1 = 10'd105; b_exp2 = 10'd6; b_exp3 = 10'd866;
a_sign0 = 4'd7; a_sign1 = 4'd11; a_sign2 = 4'd12; a_sign3 = 4'd11;
b_sign0 = 4'd16; b_sign1 = 4'd13; b_sign2 = 4'd5; b_sign3 = 4'd4;
@(posedge clk_i);
a_mant0 = 8'd148; a_mant1 = 8'd202; a_mant2 = 8'd128; a_mant3 = 8'd106;
b_mant0 = 8'd69; b_mant1 = 8'd230; b_mant2 = 8'd180; b_mant3 = 8'd217;
a_exp0 = 10'd384; a_exp1 = 10'd813; a_exp2 = 10'd119; a_exp3 = 10'd131;
b_exp0 = 10'd308; b_exp1 = 10'd736; b_exp2 = 10'd129; b_exp3 = 10'd514;
a_sign0 = 4'd12; a_sign1 = 4'd2; a_sign2 = 4'd5; a_sign3 = 4'd7;
b_sign0 = 4'd10; b_sign1 = 4'd3; b_sign2 = 4'd6; b_sign3 = 4'd10;
@(posedge clk_i);
shared_exps0 = 8'd125;
shared_exps1 = 8'd124;
a_mant0 = 8'd156; a_mant1 = 8'd10; a_mant2 = 8'd239; a_mant3 = 8'd173;
b_mant0 = 8'd199; b_mant1 = 8'd72; b_mant2 = 8'd208; b_mant3 = 8'd230;
a_exp0 = 10'd337; a_exp1 = 10'd42; a_exp2 = 10'd776; a_exp3 = 10'd722;
b_exp0 = 10'd271; b_exp1 = 10'd865; b_exp2 = 10'd280; b_exp3 = 10'd933;
a_sign0 = 4'd10; a_sign1 = 4'd3; a_sign2 = 4'd12; a_sign3 = 4'd9;
b_sign0 = 4'd3; b_sign1 = 4'd16; b_sign2 = 4'd4; b_sign3 = 4'd9;
@(posedge clk_i);
a_mant0 = 8'd234; a_mant1 = 8'd146; a_mant2 = 8'd117; a_mant3 = 8'd235;
b_mant0 = 8'd16; b_mant1 = 8'd41; b_mant2 = 8'd178; b_mant3 = 8'd128;
a_exp0 = 10'd472; a_exp1 = 10'd99; a_exp2 = 10'd1011; a_exp3 = 10'd377;
b_exp0 = 10'd612; b_exp1 = 10'd199; b_exp2 = 10'd635; b_exp3 = 10'd745;
a_sign0 = 4'd14; a_sign1 = 4'd2; a_sign2 = 4'd0; a_sign3 = 4'd15;
b_sign0 = 4'd9; b_sign1 = 4'd3; b_sign2 = 4'd11; b_sign3 = 4'd5;
@(posedge clk_i);
a_mant0 = 8'd237; a_mant1 = 8'd226; a_mant2 = 8'd78; a_mant3 = 8'd37;
b_mant0 = 8'd11; b_mant1 = 8'd182; b_mant2 = 8'd204; b_mant3 = 8'd63;
a_exp0 = 10'd706; a_exp1 = 10'd121; a_exp2 = 10'd5; a_exp3 = 10'd559;
b_exp0 = 10'd435; b_exp1 = 10'd792; b_exp2 = 10'd425; b_exp3 = 10'd596;
a_sign0 = 4'd13; a_sign1 = 4'd15; a_sign2 = 4'd9; a_sign3 = 4'd14;
b_sign0 = 4'd3; b_sign1 = 4'd0; b_sign2 = 4'd9; b_sign3 = 4'd15;
@(posedge clk_i);
a_mant0 = 8'd225; a_mant1 = 8'd92; a_mant2 = 8'd121; a_mant3 = 8'd214;
b_mant0 = 8'd17; b_mant1 = 8'd158; b_mant2 = 8'd154; b_mant3 = 8'd221;
a_exp0 = 10'd583; a_exp1 = 10'd784; a_exp2 = 10'd669; a_exp3 = 10'd306;
b_exp0 = 10'd427; b_exp1 = 10'd552; b_exp2 = 10'd711; b_exp3 = 10'd461;
a_sign0 = 4'd16; a_sign1 = 4'd9; a_sign2 = 4'd6; a_sign3 = 4'd11;
b_sign0 = 4'd11; b_sign1 = 4'd4; b_sign2 = 4'd2; b_sign3 = 4'd15;
@(posedge clk_i);
a_mant0 = 8'd14; a_mant1 = 8'd102; a_mant2 = 8'd118; a_mant3 = 8'd136;
b_mant0 = 8'd160; b_mant1 = 8'd72; b_mant2 = 8'd7; b_mant3 = 8'd211;
a_exp0 = 10'd555; a_exp1 = 10'd32; a_exp2 = 10'd978; a_exp3 = 10'd892;
b_exp0 = 10'd374; b_exp1 = 10'd681; b_exp2 = 10'd63; b_exp3 = 10'd17;
a_sign0 = 4'd16; a_sign1 = 4'd9; a_sign2 = 4'd1; a_sign3 = 4'd15;
b_sign0 = 4'd1; b_sign1 = 4'd16; b_sign2 = 4'd0; b_sign3 = 4'd16;
@(posedge clk_i);
a_mant0 = 8'd238; a_mant1 = 8'd232; a_mant2 = 8'd55; a_mant3 = 8'd82;
b_mant0 = 8'd246; b_mant1 = 8'd105; b_mant2 = 8'd241; b_mant3 = 8'd3;
a_exp0 = 10'd140; a_exp1 = 10'd378; a_exp2 = 10'd963; a_exp3 = 10'd190;
b_exp0 = 10'd148; b_exp1 = 10'd226; b_exp2 = 10'd584; b_exp3 = 10'd648;
a_sign0 = 4'd0; a_sign1 = 4'd13; a_sign2 = 4'd8; a_sign3 = 4'd3;
b_sign0 = 4'd0; b_sign1 = 4'd2; b_sign2 = 4'd12; b_sign3 = 4'd2;
@(posedge clk_i);
a_mant0 = 8'd139; a_mant1 = 8'd46; a_mant2 = 8'd90; a_mant3 = 8'd46;
b_mant0 = 8'd104; b_mant1 = 8'd101; b_mant2 = 8'd24; b_mant3 = 8'd172;
a_exp0 = 10'd598; a_exp1 = 10'd430; a_exp2 = 10'd864; a_exp3 = 10'd678;
b_exp0 = 10'd1008; b_exp1 = 10'd939; b_exp2 = 10'd135; b_exp3 = 10'd362;
a_sign0 = 4'd0; a_sign1 = 4'd0; a_sign2 = 4'd15; a_sign3 = 4'd5;
b_sign0 = 4'd4; b_sign1 = 4'd1; b_sign2 = 4'd13; b_sign3 = 4'd5;
@(posedge clk_i);
a_mant0 = 8'd113; a_mant1 = 8'd117; a_mant2 = 8'd8; a_mant3 = 8'd22;
b_mant0 = 8'd25; b_mant1 = 8'd227; b_mant2 = 8'd19; b_mant3 = 8'd100;
a_exp0 = 10'd708; a_exp1 = 10'd556; a_exp2 = 10'd493; a_exp3 = 10'd680;
b_exp0 = 10'd167; b_exp1 = 10'd338; b_exp2 = 10'd145; b_exp3 = 10'd238;
a_sign0 = 4'd3; a_sign1 = 4'd13; a_sign2 = 4'd9; a_sign3 = 4'd3;
b_sign0 = 4'd9; b_sign1 = 4'd5; b_sign2 = 4'd2; b_sign3 = 4'd12;
@(posedge clk_i);
shared_exps0 = 8'd139;
shared_exps1 = 8'd143;
a_mant0 = 8'd83; a_mant1 = 8'd76; a_mant2 = 8'd23; a_mant3 = 8'd12;
b_mant0 = 8'd107; b_mant1 = 8'd84; b_mant2 = 8'd220; b_mant3 = 8'd168;
a_exp0 = 10'd577; a_exp1 = 10'd500; a_exp2 = 10'd307; a_exp3 = 10'd920;
b_exp0 = 10'd442; b_exp1 = 10'd693; b_exp2 = 10'd741; b_exp3 = 10'd861;
a_sign0 = 4'd8; a_sign1 = 4'd2; a_sign2 = 4'd11; a_sign3 = 4'd0;
b_sign0 = 4'd14; b_sign1 = 4'd4; b_sign2 = 4'd5; b_sign3 = 4'd11;
@(posedge clk_i);
a_mant0 = 8'd167; a_mant1 = 8'd23; a_mant2 = 8'd68; a_mant3 = 8'd182;
b_mant0 = 8'd171; b_mant1 = 8'd138; b_mant2 = 8'd244; b_mant3 = 8'd139;
a_exp0 = 10'd8; a_exp1 = 10'd522; a_exp2 = 10'd549; a_exp3 = 10'd883;
b_exp0 = 10'd455; b_exp1 = 10'd501; b_exp2 = 10'd263; b_exp3 = 10'd713;
a_sign0 = 4'd9; a_sign1 = 4'd6; a_sign2 = 4'd11; a_sign3 = 4'd14;
b_sign0 = 4'd5; b_sign1 = 4'd8; b_sign2 = 4'd15; b_sign3 = 4'd10;
@(posedge clk_i);
a_mant0 = 8'd9; a_mant1 = 8'd149; a_mant2 = 8'd95; a_mant3 = 8'd40;
b_mant0 = 8'd161; b_mant1 = 8'd220; b_mant2 = 8'd198; b_mant3 = 8'd30;
a_exp0 = 10'd926; a_exp1 = 10'd285; a_exp2 = 10'd79; a_exp3 = 10'd303;
b_exp0 = 10'd823; b_exp1 = 10'd816; b_exp2 = 10'd1011; b_exp3 = 10'd155;
a_sign0 = 4'd13; a_sign1 = 4'd9; a_sign2 = 4'd7; a_sign3 = 4'd11;
b_sign0 = 4'd3; b_sign1 = 4'd12; b_sign2 = 4'd14; b_sign3 = 4'd3;
@(posedge clk_i);
a_mant0 = 8'd104; a_mant1 = 8'd204; a_mant2 = 8'd229; a_mant3 = 8'd24;
b_mant0 = 8'd216; b_mant1 = 8'd148; b_mant2 = 8'd210; b_mant3 = 8'd235;
a_exp0 = 10'd386; a_exp1 = 10'd100; a_exp2 = 10'd930; a_exp3 = 10'd596;
b_exp0 = 10'd294; b_exp1 = 10'd126; b_exp2 = 10'd578; b_exp3 = 10'd937;
a_sign0 = 4'd9; a_sign1 = 4'd4; a_sign2 = 4'd11; a_sign3 = 4'd5;
b_sign0 = 4'd15; b_sign1 = 4'd12; b_sign2 = 4'd11; b_sign3 = 4'd5;
@(posedge clk_i);
a_mant0 = 8'd224; a_mant1 = 8'd46; a_mant2 = 8'd15; a_mant3 = 8'd23;
b_mant0 = 8'd252; b_mant1 = 8'd11; b_mant2 = 8'd187; b_mant3 = 8'd171;
a_exp0 = 10'd707; a_exp1 = 10'd127; a_exp2 = 10'd158; a_exp3 = 10'd602;
b_exp0 = 10'd198; b_exp1 = 10'd552; b_exp2 = 10'd550; b_exp3 = 10'd511;
a_sign0 = 4'd11; a_sign1 = 4'd1; a_sign2 = 4'd16; a_sign3 = 4'd2;
b_sign0 = 4'd5; b_sign1 = 4'd7; b_sign2 = 4'd2; b_sign3 = 4'd13;
@(posedge clk_i);
a_mant0 = 8'd183; a_mant1 = 8'd239; a_mant2 = 8'd65; a_mant3 = 8'd56;
b_mant0 = 8'd23; b_mant1 = 8'd215; b_mant2 = 8'd56; b_mant3 = 8'd37;
a_exp0 = 10'd705; a_exp1 = 10'd986; a_exp2 = 10'd713; a_exp3 = 10'd228;
b_exp0 = 10'd372; b_exp1 = 10'd986; b_exp2 = 10'd868; b_exp3 = 10'd254;
a_sign0 = 4'd5; a_sign1 = 4'd9; a_sign2 = 4'd3; a_sign3 = 4'd4;
b_sign0 = 4'd3; b_sign1 = 4'd8; b_sign2 = 4'd10; b_sign3 = 4'd5;
@(posedge clk_i);
a_mant0 = 8'd143; a_mant1 = 8'd34; a_mant2 = 8'd126; a_mant3 = 8'd108;
b_mant0 = 8'd235; b_mant1 = 8'd139; b_mant2 = 8'd118; b_mant3 = 8'd49;
a_exp0 = 10'd244; a_exp1 = 10'd18; a_exp2 = 10'd335; a_exp3 = 10'd3;
b_exp0 = 10'd834; b_exp1 = 10'd751; b_exp2 = 10'd963; b_exp3 = 10'd378;
a_sign0 = 4'd13; a_sign1 = 4'd7; a_sign2 = 4'd14; a_sign3 = 4'd13;
b_sign0 = 4'd15; b_sign1 = 4'd4; b_sign2 = 4'd14; b_sign3 = 4'd2;
@(posedge clk_i);
a_mant0 = 8'd144; a_mant1 = 8'd166; a_mant2 = 8'd152; a_mant3 = 8'd56;
b_mant0 = 8'd130; b_mant1 = 8'd84; b_mant2 = 8'd3; b_mant3 = 8'd42;
a_exp0 = 10'd174; a_exp1 = 10'd536; a_exp2 = 10'd281; a_exp3 = 10'd340;
b_exp0 = 10'd904; b_exp1 = 10'd541; b_exp2 = 10'd832; b_exp3 = 10'd323;
a_sign0 = 4'd16; a_sign1 = 4'd2; a_sign2 = 4'd1; a_sign3 = 4'd8;
b_sign0 = 4'd13; b_sign1 = 4'd12; b_sign2 = 4'd9; b_sign3 = 4'd8;
@(posedge clk_i);
shared_exps0 = 8'd128;
shared_exps1 = 8'd130;
a_mant0 = 8'd190; a_mant1 = 8'd220; a_mant2 = 8'd209; a_mant3 = 8'd145;
b_mant0 = 8'd11; b_mant1 = 8'd208; b_mant2 = 8'd86; b_mant3 = 8'd249;
a_exp0 = 10'd472; a_exp1 = 10'd832; a_exp2 = 10'd693; a_exp3 = 10'd30;
b_exp0 = 10'd434; b_exp1 = 10'd940; b_exp2 = 10'd354; b_exp3 = 10'd174;
a_sign0 = 4'd9; a_sign1 = 4'd0; a_sign2 = 4'd9; a_sign3 = 4'd4;
b_sign0 = 4'd12; b_sign1 = 4'd6; b_sign2 = 4'd15; b_sign3 = 4'd10;
@(posedge clk_i);
a_mant0 = 8'd160; a_mant1 = 8'd227; a_mant2 = 8'd231; a_mant3 = 8'd230;
b_mant0 = 8'd110; b_mant1 = 8'd127; b_mant2 = 8'd8; b_mant3 = 8'd171;
a_exp0 = 10'd799; a_exp1 = 10'd64; a_exp2 = 10'd8; a_exp3 = 10'd200;
b_exp0 = 10'd808; b_exp1 = 10'd637; b_exp2 = 10'd960; b_exp3 = 10'd152;
a_sign0 = 4'd10; a_sign1 = 4'd2; a_sign2 = 4'd9; a_sign3 = 4'd4;
b_sign0 = 4'd5; b_sign1 = 4'd3; b_sign2 = 4'd5; b_sign3 = 4'd11;
@(posedge clk_i);
a_mant0 = 8'd144; a_mant1 = 8'd165; a_mant2 = 8'd17; a_mant3 = 8'd11;
b_mant0 = 8'd170; b_mant1 = 8'd129; b_mant2 = 8'd98; b_mant3 = 8'd123;
a_exp0 = 10'd202; a_exp1 = 10'd617; a_exp2 = 10'd914; a_exp3 = 10'd805;
b_exp0 = 10'd979; b_exp1 = 10'd855; b_exp2 = 10'd798; b_exp3 = 10'd756;
a_sign0 = 4'd0; a_sign1 = 4'd7; a_sign2 = 4'd14; a_sign3 = 4'd15;
b_sign0 = 4'd9; b_sign1 = 4'd6; b_sign2 = 4'd1; b_sign3 = 4'd3;
@(posedge clk_i);
a_mant0 = 8'd83; a_mant1 = 8'd18; a_mant2 = 8'd1; a_mant3 = 8'd207;
b_mant0 = 8'd232; b_mant1 = 8'd204; b_mant2 = 8'd75; b_mant3 = 8'd230;
a_exp0 = 10'd639; a_exp1 = 10'd373; a_exp2 = 10'd156; a_exp3 = 10'd712;
b_exp0 = 10'd624; b_exp1 = 10'd939; b_exp2 = 10'd706; b_exp3 = 10'd810;
a_sign0 = 4'd4; a_sign1 = 4'd2; a_sign2 = 4'd11; a_sign3 = 4'd0;
b_sign0 = 4'd5; b_sign1 = 4'd16; b_sign2 = 4'd9; b_sign3 = 4'd14;
@(posedge clk_i);
a_mant0 = 8'd177; a_mant1 = 8'd108; a_mant2 = 8'd228; a_mant3 = 8'd214;
b_mant0 = 8'd212; b_mant1 = 8'd174; b_mant2 = 8'd9; b_mant3 = 8'd161;
a_exp0 = 10'd155; a_exp1 = 10'd831; a_exp2 = 10'd511; a_exp3 = 10'd568;
b_exp0 = 10'd956; b_exp1 = 10'd320; b_exp2 = 10'd1007; b_exp3 = 10'd546;
a_sign0 = 4'd3; a_sign1 = 4'd1; a_sign2 = 4'd15; a_sign3 = 4'd0;
b_sign0 = 4'd1; b_sign1 = 4'd0; b_sign2 = 4'd8; b_sign3 = 4'd3;
@(posedge clk_i);
a_mant0 = 8'd104; a_mant1 = 8'd44; a_mant2 = 8'd169; a_mant3 = 8'd44;
b_mant0 = 8'd70; b_mant1 = 8'd114; b_mant2 = 8'd73; b_mant3 = 8'd244;
a_exp0 = 10'd705; a_exp1 = 10'd694; a_exp2 = 10'd563; a_exp3 = 10'd423;
b_exp0 = 10'd698; b_exp1 = 10'd356; b_exp2 = 10'd590; b_exp3 = 10'd55;
a_sign0 = 4'd6; a_sign1 = 4'd14; a_sign2 = 4'd10; a_sign3 = 4'd12;
b_sign0 = 4'd16; b_sign1 = 4'd15; b_sign2 = 4'd3; b_sign3 = 4'd7;
@(posedge clk_i);
a_mant0 = 8'd80; a_mant1 = 8'd88; a_mant2 = 8'd172; a_mant3 = 8'd49;
b_mant0 = 8'd105; b_mant1 = 8'd9; b_mant2 = 8'd106; b_mant3 = 8'd94;
a_exp0 = 10'd513; a_exp1 = 10'd310; a_exp2 = 10'd125; a_exp3 = 10'd461;
b_exp0 = 10'd435; b_exp1 = 10'd721; b_exp2 = 10'd390; b_exp3 = 10'd715;
a_sign0 = 4'd15; a_sign1 = 4'd13; a_sign2 = 4'd12; a_sign3 = 4'd7;
b_sign0 = 4'd14; b_sign1 = 4'd10; b_sign2 = 4'd9; b_sign3 = 4'd3;
@(posedge clk_i);
a_mant0 = 8'd2; a_mant1 = 8'd46; a_mant2 = 8'd241; a_mant3 = 8'd119;
b_mant0 = 8'd236; b_mant1 = 8'd58; b_mant2 = 8'd31; b_mant3 = 8'd7;
a_exp0 = 10'd70; a_exp1 = 10'd668; a_exp2 = 10'd487; a_exp3 = 10'd306;
b_exp0 = 10'd86; b_exp1 = 10'd753; b_exp2 = 10'd570; b_exp3 = 10'd157;
a_sign0 = 4'd7; a_sign1 = 4'd14; a_sign2 = 4'd15; a_sign3 = 4'd0;
b_sign0 = 4'd14; b_sign1 = 4'd7; b_sign2 = 4'd4; b_sign3 = 4'd5;
@(posedge clk_i);
shared_exps0 = 8'd100;
shared_exps1 = 8'd138;
rstn = 0;
@(posedge clk_i);
rstn = 1;
a_mant0 = 8'd30; a_mant1 = 8'd242; a_mant2 = 8'd24; a_mant3 = 8'd224;
b_mant0 = 8'd97; b_mant1 = 8'd221; b_mant2 = 8'd133; b_mant3 = 8'd188;
a_exp0 = 10'd52; a_exp1 = 10'd207; a_exp2 = 10'd133; a_exp3 = 10'd392;
b_exp0 = 10'd542; b_exp1 = 10'd468; b_exp2 = 10'd1008; b_exp3 = 10'd51;
a_sign0 = 4'd4; a_sign1 = 4'd12; a_sign2 = 4'd11; a_sign3 = 4'd11;
b_sign0 = 4'd0; b_sign1 = 4'd2; b_sign2 = 4'd5; b_sign3 = 4'd13;
@(posedge clk_i);
a_mant0 = 8'd235; a_mant1 = 8'd243; a_mant2 = 8'd113; a_mant3 = 8'd206;
b_mant0 = 8'd29; b_mant1 = 8'd130; b_mant2 = 8'd24; b_mant3 = 8'd153;
a_exp0 = 10'd608; a_exp1 = 10'd833; a_exp2 = 10'd314; a_exp3 = 10'd562;
b_exp0 = 10'd1004; b_exp1 = 10'd74; b_exp2 = 10'd9; b_exp3 = 10'd692;
a_sign0 = 4'd8; a_sign1 = 4'd11; a_sign2 = 4'd16; a_sign3 = 4'd16;
b_sign0 = 4'd15; b_sign1 = 4'd14; b_sign2 = 4'd2; b_sign3 = 4'd4;
@(posedge clk_i);
a_mant0 = 8'd207; a_mant1 = 8'd99; a_mant2 = 8'd131; a_mant3 = 8'd234;
b_mant0 = 8'd224; b_mant1 = 8'd241; b_mant2 = 8'd187; b_mant3 = 8'd153;
a_exp0 = 10'd859; a_exp1 = 10'd534; a_exp2 = 10'd942; a_exp3 = 10'd171;
b_exp0 = 10'd15; b_exp1 = 10'd270; b_exp2 = 10'd609; b_exp3 = 10'd510;
a_sign0 = 4'd12; a_sign1 = 4'd2; a_sign2 = 4'd8; a_sign3 = 4'd8;
b_sign0 = 4'd8; b_sign1 = 4'd3; b_sign2 = 4'd8; b_sign3 = 4'd11;
@(posedge clk_i);
a_mant0 = 8'd199; a_mant1 = 8'd175; a_mant2 = 8'd176; a_mant3 = 8'd126;
b_mant0 = 8'd87; b_mant1 = 8'd204; b_mant2 = 8'd27; b_mant3 = 8'd202;
a_exp0 = 10'd915; a_exp1 = 10'd551; a_exp2 = 10'd616; a_exp3 = 10'd382;
b_exp0 = 10'd897; b_exp1 = 10'd273; b_exp2 = 10'd773; b_exp3 = 10'd549;
a_sign0 = 4'd12; a_sign1 = 4'd11; a_sign2 = 4'd5; a_sign3 = 4'd6;
b_sign0 = 4'd6; b_sign1 = 4'd1; b_sign2 = 4'd8; b_sign3 = 4'd14;
@(posedge clk_i);
a_mant0 = 8'd169; a_mant1 = 8'd87; a_mant2 = 8'd149; a_mant3 = 8'd58;
b_mant0 = 8'd91; b_mant1 = 8'd18; b_mant2 = 8'd250; b_mant3 = 8'd179;
a_exp0 = 10'd986; a_exp1 = 10'd886; a_exp2 = 10'd483; a_exp3 = 10'd968;
b_exp0 = 10'd480; b_exp1 = 10'd370; b_exp2 = 10'd645; b_exp3 = 10'd687;
a_sign0 = 4'd14; a_sign1 = 4'd8; a_sign2 = 4'd8; a_sign3 = 4'd3;
b_sign0 = 4'd6; b_sign1 = 4'd3; b_sign2 = 4'd2; b_sign3 = 4'd1;
@(posedge clk_i);
a_mant0 = 8'd190; a_mant1 = 8'd32; a_mant2 = 8'd159; a_mant3 = 8'd88;
b_mant0 = 8'd136; b_mant1 = 8'd220; b_mant2 = 8'd40; b_mant3 = 8'd36;
a_exp0 = 10'd600; a_exp1 = 10'd893; a_exp2 = 10'd284; a_exp3 = 10'd849;
b_exp0 = 10'd42; b_exp1 = 10'd850; b_exp2 = 10'd599; b_exp3 = 10'd942;
a_sign0 = 4'd1; a_sign1 = 4'd9; a_sign2 = 4'd12; a_sign3 = 4'd8;
b_sign0 = 4'd12; b_sign1 = 4'd10; b_sign2 = 4'd16; b_sign3 = 4'd13;
@(posedge clk_i);
a_mant0 = 8'd255; a_mant1 = 8'd135; a_mant2 = 8'd111; a_mant3 = 8'd98;
b_mant0 = 8'd20; b_mant1 = 8'd94; b_mant2 = 8'd38; b_mant3 = 8'd229;
a_exp0 = 10'd831; a_exp1 = 10'd838; a_exp2 = 10'd779; a_exp3 = 10'd850;
b_exp0 = 10'd42; b_exp1 = 10'd549; b_exp2 = 10'd142; b_exp3 = 10'd684;
a_sign0 = 4'd8; a_sign1 = 4'd13; a_sign2 = 4'd1; a_sign3 = 4'd4;
b_sign0 = 4'd16; b_sign1 = 4'd9; b_sign2 = 4'd9; b_sign3 = 4'd4;
@(posedge clk_i);
shared_exps0 = 8'd109;
shared_exps1 = 8'd148;
a_mant0 = 8'd8; a_mant1 = 8'd218; a_mant2 = 8'd174; a_mant3 = 8'd203;
b_mant0 = 8'd146; b_mant1 = 8'd105; b_mant2 = 8'd191; b_mant3 = 8'd158;
a_exp0 = 10'd660; a_exp1 = 10'd749; a_exp2 = 10'd883; a_exp3 = 10'd393;
b_exp0 = 10'd452; b_exp1 = 10'd674; b_exp2 = 10'd272; b_exp3 = 10'd801;
a_sign0 = 4'd9; a_sign1 = 4'd12; a_sign2 = 4'd7; a_sign3 = 4'd11;
b_sign0 = 4'd10; b_sign1 = 4'd15; b_sign2 = 4'd11; b_sign3 = 4'd0;
@(posedge clk_i);
a_mant0 = 8'd120; a_mant1 = 8'd204; a_mant2 = 8'd161; a_mant3 = 8'd206;
b_mant0 = 8'd237; b_mant1 = 8'd116; b_mant2 = 8'd87; b_mant3 = 8'd94;
a_exp0 = 10'd102; a_exp1 = 10'd745; a_exp2 = 10'd937; a_exp3 = 10'd141;
b_exp0 = 10'd92; b_exp1 = 10'd531; b_exp2 = 10'd500; b_exp3 = 10'd315;
a_sign0 = 4'd16; a_sign1 = 4'd13; a_sign2 = 4'd5; a_sign3 = 4'd9;
b_sign0 = 4'd10; b_sign1 = 4'd4; b_sign2 = 4'd1; b_sign3 = 4'd16;
@(posedge clk_i);
a_mant0 = 8'd80; a_mant1 = 8'd64; a_mant2 = 8'd246; a_mant3 = 8'd43;
b_mant0 = 8'd191; b_mant1 = 8'd35; b_mant2 = 8'd141; b_mant3 = 8'd12;
a_exp0 = 10'd671; a_exp1 = 10'd55; a_exp2 = 10'd804; a_exp3 = 10'd887;
b_exp0 = 10'd537; b_exp1 = 10'd795; b_exp2 = 10'd350; b_exp3 = 10'd86;
a_sign0 = 4'd1; a_sign1 = 4'd15; a_sign2 = 4'd14; a_sign3 = 4'd3;
b_sign0 = 4'd2; b_sign1 = 4'd2; b_sign2 = 4'd2; b_sign3 = 4'd0;
@(posedge clk_i);
a_mant0 = 8'd92; a_mant1 = 8'd68; a_mant2 = 8'd76; a_mant3 = 8'd48;
b_mant0 = 8'd212; b_mant1 = 8'd44; b_mant2 = 8'd121; b_mant3 = 8'd202;
a_exp0 = 10'd517; a_exp1 = 10'd712; a_exp2 = 10'd4; a_exp3 = 10'd741;
b_exp0 = 10'd576; b_exp1 = 10'd505; b_exp2 = 10'd1; b_exp3 = 10'd984;
a_sign0 = 4'd3; a_sign1 = 4'd10; a_sign2 = 4'd16; a_sign3 = 4'd9;
b_sign0 = 4'd1; b_sign1 = 4'd4; b_sign2 = 4'd16; b_sign3 = 4'd5;
@(posedge clk_i);
a_mant0 = 8'd23; a_mant1 = 8'd211; a_mant2 = 8'd173; a_mant3 = 8'd109;
b_mant0 = 8'd111; b_mant1 = 8'd236; b_mant2 = 8'd201; b_mant3 = 8'd211;
a_exp0 = 10'd585; a_exp1 = 10'd800; a_exp2 = 10'd183; a_exp3 = 10'd516;
b_exp0 = 10'd925; b_exp1 = 10'd903; b_exp2 = 10'd556; b_exp3 = 10'd319;
a_sign0 = 4'd2; a_sign1 = 4'd3; a_sign2 = 4'd9; a_sign3 = 4'd1;
b_sign0 = 4'd1; b_sign1 = 4'd16; b_sign2 = 4'd13; b_sign3 = 4'd10;
@(posedge clk_i);
a_mant0 = 8'd59; a_mant1 = 8'd233; a_mant2 = 8'd35; a_mant3 = 8'd44;
b_mant0 = 8'd176; b_mant1 = 8'd227; b_mant2 = 8'd250; b_mant3 = 8'd174;
a_exp0 = 10'd652; a_exp1 = 10'd20; a_exp2 = 10'd56; a_exp3 = 10'd211;
b_exp0 = 10'd822; b_exp1 = 10'd691; b_exp2 = 10'd500; b_exp3 = 10'd508;
a_sign0 = 4'd14; a_sign1 = 4'd8; a_sign2 = 4'd13; a_sign3 = 4'd3;
b_sign0 = 4'd12; b_sign1 = 4'd7; b_sign2 = 4'd15; b_sign3 = 4'd3;
@(posedge clk_i);
a_mant0 = 8'd185; a_mant1 = 8'd140; a_mant2 = 8'd29; a_mant3 = 8'd245;
b_mant0 = 8'd222; b_mant1 = 8'd236; b_mant2 = 8'd139; b_mant3 = 8'd168;
a_exp0 = 10'd417; a_exp1 = 10'd400; a_exp2 = 10'd411; a_exp3 = 10'd965;
b_exp0 = 10'd523; b_exp1 = 10'd919; b_exp2 = 10'd777; b_exp3 = 10'd570;
a_sign0 = 4'd12; a_sign1 = 4'd16; a_sign2 = 4'd16; a_sign3 = 4'd15;
b_sign0 = 4'd10; b_sign1 = 4'd4; b_sign2 = 4'd5; b_sign3 = 4'd6;
@(posedge clk_i);
a_mant0 = 8'd186; a_mant1 = 8'd51; a_mant2 = 8'd165; a_mant3 = 8'd63;
b_mant0 = 8'd128; b_mant1 = 8'd72; b_mant2 = 8'd115; b_mant3 = 8'd108;
a_exp0 = 10'd734; a_exp1 = 10'd944; a_exp2 = 10'd525; a_exp3 = 10'd84;
b_exp0 = 10'd1009; b_exp1 = 10'd26; b_exp2 = 10'd703; b_exp3 = 10'd260;
a_sign0 = 4'd16; a_sign1 = 4'd7; a_sign2 = 4'd16; a_sign3 = 4'd9;
b_sign0 = 4'd4; b_sign1 = 4'd16; b_sign2 = 4'd15; b_sign3 = 4'd7;
@(posedge clk_i);
shared_exps0 = 8'd117;
shared_exps1 = 8'd126;
a_mant0 = 8'd253; a_mant1 = 8'd158; a_mant2 = 8'd231; a_mant3 = 8'd151;
b_mant0 = 8'd240; b_mant1 = 8'd79; b_mant2 = 8'd93; b_mant3 = 8'd210;
a_exp0 = 10'd444; a_exp1 = 10'd59; a_exp2 = 10'd27; a_exp3 = 10'd7;
b_exp0 = 10'd197; b_exp1 = 10'd318; b_exp2 = 10'd351; b_exp3 = 10'd350;
a_sign0 = 4'd8; a_sign1 = 4'd3; a_sign2 = 4'd14; a_sign3 = 4'd10;
b_sign0 = 4'd2; b_sign1 = 4'd3; b_sign2 = 4'd12; b_sign3 = 4'd10;
@(posedge clk_i);
a_mant0 = 8'd136; a_mant1 = 8'd99; a_mant2 = 8'd26; a_mant3 = 8'd19;
b_mant0 = 8'd231; b_mant1 = 8'd63; b_mant2 = 8'd59; b_mant3 = 8'd232;
a_exp0 = 10'd982; a_exp1 = 10'd1021; a_exp2 = 10'd676; a_exp3 = 10'd729;
b_exp0 = 10'd445; b_exp1 = 10'd705; b_exp2 = 10'd520; b_exp3 = 10'd463;
a_sign0 = 4'd13; a_sign1 = 4'd11; a_sign2 = 4'd14; a_sign3 = 4'd8;
b_sign0 = 4'd1; b_sign1 = 4'd6; b_sign2 = 4'd7; b_sign3 = 4'd10;
@(posedge clk_i);
a_mant0 = 8'd90; a_mant1 = 8'd172; a_mant2 = 8'd15; a_mant3 = 8'd48;
b_mant0 = 8'd229; b_mant1 = 8'd35; b_mant2 = 8'd243; b_mant3 = 8'd2;
a_exp0 = 10'd945; a_exp1 = 10'd682; a_exp2 = 10'd920; a_exp3 = 10'd583;
b_exp0 = 10'd383; b_exp1 = 10'd201; b_exp2 = 10'd515; b_exp3 = 10'd208;
a_sign0 = 4'd14; a_sign1 = 4'd0; a_sign2 = 4'd9; a_sign3 = 4'd13;
b_sign0 = 4'd13; b_sign1 = 4'd6; b_sign2 = 4'd4; b_sign3 = 4'd10;
@(posedge clk_i);
a_mant0 = 8'd12; a_mant1 = 8'd235; a_mant2 = 8'd148; a_mant3 = 8'd194;
b_mant0 = 8'd104; b_mant1 = 8'd136; b_mant2 = 8'd34; b_mant3 = 8'd14;
a_exp0 = 10'd648; a_exp1 = 10'd62; a_exp2 = 10'd252; a_exp3 = 10'd791;
b_exp0 = 10'd286; b_exp1 = 10'd615; b_exp2 = 10'd880; b_exp3 = 10'd888;
a_sign0 = 4'd1; a_sign1 = 4'd0; a_sign2 = 4'd16; a_sign3 = 4'd5;
b_sign0 = 4'd5; b_sign1 = 4'd0; b_sign2 = 4'd9; b_sign3 = 4'd15;
@(posedge clk_i);
a_mant0 = 8'd84; a_mant1 = 8'd91; a_mant2 = 8'd167; a_mant3 = 8'd140;
b_mant0 = 8'd140; b_mant1 = 8'd216; b_mant2 = 8'd115; b_mant3 = 8'd32;
a_exp0 = 10'd381; a_exp1 = 10'd150; a_exp2 = 10'd531; a_exp3 = 10'd0;
b_exp0 = 10'd348; b_exp1 = 10'd955; b_exp2 = 10'd37; b_exp3 = 10'd744;
a_sign0 = 4'd12; a_sign1 = 4'd14; a_sign2 = 4'd8; a_sign3 = 4'd3;
b_sign0 = 4'd16; b_sign1 = 4'd3; b_sign2 = 4'd9; b_sign3 = 4'd11;
@(posedge clk_i);
a_mant0 = 8'd57; a_mant1 = 8'd117; a_mant2 = 8'd57; a_mant3 = 8'd58;
b_mant0 = 8'd68; b_mant1 = 8'd206; b_mant2 = 8'd246; b_mant3 = 8'd98;
a_exp0 = 10'd105; a_exp1 = 10'd10; a_exp2 = 10'd762; a_exp3 = 10'd1010;
b_exp0 = 10'd878; b_exp1 = 10'd916; b_exp2 = 10'd128; b_exp3 = 10'd551;
a_sign0 = 4'd16; a_sign1 = 4'd16; a_sign2 = 4'd9; a_sign3 = 4'd16;
b_sign0 = 4'd12; b_sign1 = 4'd14; b_sign2 = 4'd11; b_sign3 = 4'd6;
@(posedge clk_i);
a_mant0 = 8'd63; a_mant1 = 8'd140; a_mant2 = 8'd193; a_mant3 = 8'd18;
b_mant0 = 8'd33; b_mant1 = 8'd209; b_mant2 = 8'd229; b_mant3 = 8'd201;
a_exp0 = 10'd52; a_exp1 = 10'd810; a_exp2 = 10'd5; a_exp3 = 10'd916;
b_exp0 = 10'd731; b_exp1 = 10'd780; b_exp2 = 10'd284; b_exp3 = 10'd827;
a_sign0 = 4'd0; a_sign1 = 4'd10; a_sign2 = 4'd4; a_sign3 = 4'd11;
b_sign0 = 4'd12; b_sign1 = 4'd2; b_sign2 = 4'd5; b_sign3 = 4'd14;
@(posedge clk_i);
a_mant0 = 8'd99; a_mant1 = 8'd81; a_mant2 = 8'd98; a_mant3 = 8'd65;
b_mant0 = 8'd248; b_mant1 = 8'd200; b_mant2 = 8'd249; b_mant3 = 8'd64;
a_exp0 = 10'd524; a_exp1 = 10'd413; a_exp2 = 10'd632; a_exp3 = 10'd967;
b_exp0 = 10'd390; b_exp1 = 10'd611; b_exp2 = 10'd751; b_exp3 = 10'd80;
a_sign0 = 4'd8; a_sign1 = 4'd4; a_sign2 = 4'd13; a_sign3 = 4'd2;
b_sign0 = 4'd12; b_sign1 = 4'd7; b_sign2 = 4'd10; b_sign3 = 4'd6;
@(posedge clk_i);
shared_exps0 = 8'd122;
shared_exps1 = 8'd114;
a_mant0 = 8'd203; a_mant1 = 8'd100; a_mant2 = 8'd247; a_mant3 = 8'd151;
b_mant0 = 8'd152; b_mant1 = 8'd183; b_mant2 = 8'd237; b_mant3 = 8'd155;
a_exp0 = 10'd465; a_exp1 = 10'd928; a_exp2 = 10'd644; a_exp3 = 10'd370;
b_exp0 = 10'd886; b_exp1 = 10'd609; b_exp2 = 10'd848; b_exp3 = 10'd6;
a_sign0 = 4'd16; a_sign1 = 4'd0; a_sign2 = 4'd10; a_sign3 = 4'd7;
b_sign0 = 4'd6; b_sign1 = 4'd15; b_sign2 = 4'd2; b_sign3 = 4'd6;
@(posedge clk_i);
a_mant0 = 8'd152; a_mant1 = 8'd177; a_mant2 = 8'd216; a_mant3 = 8'd104;
b_mant0 = 8'd167; b_mant1 = 8'd113; b_mant2 = 8'd147; b_mant3 = 8'd68;
a_exp0 = 10'd1013; a_exp1 = 10'd906; a_exp2 = 10'd912; a_exp3 = 10'd452;
b_exp0 = 10'd1016; b_exp1 = 10'd840; b_exp2 = 10'd266; b_exp3 = 10'd989;
a_sign0 = 4'd9; a_sign1 = 4'd12; a_sign2 = 4'd11; a_sign3 = 4'd1;
b_sign0 = 4'd12; b_sign1 = 4'd6; b_sign2 = 4'd2; b_sign3 = 4'd12;
@(posedge clk_i);
a_mant0 = 8'd53; a_mant1 = 8'd127; a_mant2 = 8'd218; a_mant3 = 8'd84;
b_mant0 = 8'd122; b_mant1 = 8'd216; b_mant2 = 8'd166; b_mant3 = 8'd248;
a_exp0 = 10'd720; a_exp1 = 10'd28; a_exp2 = 10'd186; a_exp3 = 10'd448;
b_exp0 = 10'd621; b_exp1 = 10'd630; b_exp2 = 10'd828; b_exp3 = 10'd983;
a_sign0 = 4'd8; a_sign1 = 4'd0; a_sign2 = 4'd0; a_sign3 = 4'd7;
b_sign0 = 4'd2; b_sign1 = 4'd8; b_sign2 = 4'd15; b_sign3 = 4'd5;
@(posedge clk_i);
a_mant0 = 8'd127; a_mant1 = 8'd7; a_mant2 = 8'd72; a_mant3 = 8'd62;
b_mant0 = 8'd246; b_mant1 = 8'd196; b_mant2 = 8'd181; b_mant3 = 8'd15;
a_exp0 = 10'd443; a_exp1 = 10'd84; a_exp2 = 10'd1004; a_exp3 = 10'd984;
b_exp0 = 10'd897; b_exp1 = 10'd305; b_exp2 = 10'd316; b_exp3 = 10'd862;
a_sign0 = 4'd10; a_sign1 = 4'd10; a_sign2 = 4'd12; a_sign3 = 4'd9;
b_sign0 = 4'd2; b_sign1 = 4'd2; b_sign2 = 4'd10; b_sign3 = 4'd7;
@(posedge clk_i);
a_mant0 = 8'd197; a_mant1 = 8'd139; a_mant2 = 8'd111; a_mant3 = 8'd101;
b_mant0 = 8'd235; b_mant1 = 8'd114; b_mant2 = 8'd12; b_mant3 = 8'd100;
a_exp0 = 10'd600; a_exp1 = 10'd170; a_exp2 = 10'd662; a_exp3 = 10'd593;
b_exp0 = 10'd617; b_exp1 = 10'd630; b_exp2 = 10'd449; b_exp3 = 10'd319;
a_sign0 = 4'd9; a_sign1 = 4'd3; a_sign2 = 4'd13; a_sign3 = 4'd10;
b_sign0 = 4'd2; b_sign1 = 4'd15; b_sign2 = 4'd15; b_sign3 = 4'd1;
@(posedge clk_i);
a_mant0 = 8'd204; a_mant1 = 8'd65; a_mant2 = 8'd238; a_mant3 = 8'd176;
b_mant0 = 8'd254; b_mant1 = 8'd233; b_mant2 = 8'd243; b_mant3 = 8'd84;
a_exp0 = 10'd829; a_exp1 = 10'd544; a_exp2 = 10'd751; a_exp3 = 10'd493;
b_exp0 = 10'd7; b_exp1 = 10'd29; b_exp2 = 10'd460; b_exp3 = 10'd459;
a_sign0 = 4'd8; a_sign1 = 4'd8; a_sign2 = 4'd7; a_sign3 = 4'd13;
b_sign0 = 4'd14; b_sign1 = 4'd3; b_sign2 = 4'd6; b_sign3 = 4'd9;
@(posedge clk_i);
a_mant0 = 8'd248; a_mant1 = 8'd183; a_mant2 = 8'd205; a_mant3 = 8'd239;
b_mant0 = 8'd37; b_mant1 = 8'd87; b_mant2 = 8'd126; b_mant3 = 8'd192;
a_exp0 = 10'd876; a_exp1 = 10'd133; a_exp2 = 10'd949; a_exp3 = 10'd170;
b_exp0 = 10'd332; b_exp1 = 10'd150; b_exp2 = 10'd553; b_exp3 = 10'd325;
a_sign0 = 4'd16; a_sign1 = 4'd14; a_sign2 = 4'd10; a_sign3 = 4'd13;
b_sign0 = 4'd12; b_sign1 = 4'd5; b_sign2 = 4'd13; b_sign3 = 4'd3;
@(posedge clk_i);
a_mant0 = 8'd223; a_mant1 = 8'd80; a_mant2 = 8'd223; a_mant3 = 8'd26;
b_mant0 = 8'd148; b_mant1 = 8'd65; b_mant2 = 8'd231; b_mant3 = 8'd155;
a_exp0 = 10'd489; a_exp1 = 10'd864; a_exp2 = 10'd97; a_exp3 = 10'd757;
b_exp0 = 10'd144; b_exp1 = 10'd633; b_exp2 = 10'd486; b_exp3 = 10'd685;
a_sign0 = 4'd12; a_sign1 = 4'd8; a_sign2 = 4'd3; a_sign3 = 4'd7;
b_sign0 = 4'd1; b_sign1 = 4'd6; b_sign2 = 4'd13; b_sign3 = 4'd14;
@(posedge clk_i);
shared_exps0 = 8'd136;
shared_exps1 = 8'd133;
rstn = 0;
@(posedge clk_i);
rstn = 1;
a_mant0 = 8'd210; a_mant1 = 8'd182; a_mant2 = 8'd82; a_mant3 = 8'd60;
b_mant0 = 8'd207; b_mant1 = 8'd55; b_mant2 = 8'd37; b_mant3 = 8'd5;
a_exp0 = 10'd105; a_exp1 = 10'd527; a_exp2 = 10'd910; a_exp3 = 10'd584;
b_exp0 = 10'd534; b_exp1 = 10'd390; b_exp2 = 10'd899; b_exp3 = 10'd616;
a_sign0 = 4'd13; a_sign1 = 4'd12; a_sign2 = 4'd3; a_sign3 = 4'd16;
b_sign0 = 4'd14; b_sign1 = 4'd9; b_sign2 = 4'd13; b_sign3 = 4'd2;
@(posedge clk_i);
a_mant0 = 8'd195; a_mant1 = 8'd67; a_mant2 = 8'd40; a_mant3 = 8'd199;
b_mant0 = 8'd35; b_mant1 = 8'd50; b_mant2 = 8'd70; b_mant3 = 8'd180;
a_exp0 = 10'd228; a_exp1 = 10'd238; a_exp2 = 10'd228; a_exp3 = 10'd193;
b_exp0 = 10'd515; b_exp1 = 10'd193; b_exp2 = 10'd172; b_exp3 = 10'd319;
a_sign0 = 4'd8; a_sign1 = 4'd16; a_sign2 = 4'd0; a_sign3 = 4'd8;
b_sign0 = 4'd9; b_sign1 = 4'd5; b_sign2 = 4'd12; b_sign3 = 4'd8;
@(posedge clk_i);
a_mant0 = 8'd27; a_mant1 = 8'd223; a_mant2 = 8'd96; a_mant3 = 8'd213;
b_mant0 = 8'd50; b_mant1 = 8'd70; b_mant2 = 8'd110; b_mant3 = 8'd168;
a_exp0 = 10'd35; a_exp1 = 10'd465; a_exp2 = 10'd870; a_exp3 = 10'd608;
b_exp0 = 10'd259; b_exp1 = 10'd474; b_exp2 = 10'd235; b_exp3 = 10'd880;
a_sign0 = 4'd9; a_sign1 = 4'd1; a_sign2 = 4'd14; a_sign3 = 4'd8;
b_sign0 = 4'd3; b_sign1 = 4'd6; b_sign2 = 4'd0; b_sign3 = 4'd12;
@(posedge clk_i);
a_mant0 = 8'd123; a_mant1 = 8'd194; a_mant2 = 8'd126; a_mant3 = 8'd234;
b_mant0 = 8'd166; b_mant1 = 8'd130; b_mant2 = 8'd49; b_mant3 = 8'd231;
a_exp0 = 10'd162; a_exp1 = 10'd342; a_exp2 = 10'd493; a_exp3 = 10'd502;
b_exp0 = 10'd532; b_exp1 = 10'd983; b_exp2 = 10'd373; b_exp3 = 10'd632;
a_sign0 = 4'd16; a_sign1 = 4'd2; a_sign2 = 4'd8; a_sign3 = 4'd9;
b_sign0 = 4'd1; b_sign1 = 4'd7; b_sign2 = 4'd8; b_sign3 = 4'd12;
@(posedge clk_i);
a_mant0 = 8'd64; a_mant1 = 8'd37; a_mant2 = 8'd118; a_mant3 = 8'd68;
b_mant0 = 8'd236; b_mant1 = 8'd210; b_mant2 = 8'd147; b_mant3 = 8'd191;
a_exp0 = 10'd426; a_exp1 = 10'd180; a_exp2 = 10'd409; a_exp3 = 10'd729;
b_exp0 = 10'd672; b_exp1 = 10'd241; b_exp2 = 10'd72; b_exp3 = 10'd10;
a_sign0 = 4'd14; a_sign1 = 4'd2; a_sign2 = 4'd2; a_sign3 = 4'd16;
b_sign0 = 4'd1; b_sign1 = 4'd2; b_sign2 = 4'd10; b_sign3 = 4'd7;
@(posedge clk_i);
a_mant0 = 8'd230; a_mant1 = 8'd188; a_mant2 = 8'd40; a_mant3 = 8'd146;
b_mant0 = 8'd107; b_mant1 = 8'd162; b_mant2 = 8'd121; b_mant3 = 8'd19;
a_exp0 = 10'd796; a_exp1 = 10'd128; a_exp2 = 10'd716; a_exp3 = 10'd174;
b_exp0 = 10'd380; b_exp1 = 10'd297; b_exp2 = 10'd305; b_exp3 = 10'd821;
a_sign0 = 4'd15; a_sign1 = 4'd14; a_sign2 = 4'd11; a_sign3 = 4'd7;
b_sign0 = 4'd0; b_sign1 = 4'd6; b_sign2 = 4'd2; b_sign3 = 4'd6;
@(posedge clk_i);
a_mant0 = 8'd110; a_mant1 = 8'd51; a_mant2 = 8'd216; a_mant3 = 8'd125;
b_mant0 = 8'd226; b_mant1 = 8'd110; b_mant2 = 8'd25; b_mant3 = 8'd4;
a_exp0 = 10'd115; a_exp1 = 10'd735; a_exp2 = 10'd197; a_exp3 = 10'd839;
b_exp0 = 10'd583; b_exp1 = 10'd757; b_exp2 = 10'd638; b_exp3 = 10'd621;
a_sign0 = 4'd16; a_sign1 = 4'd6; a_sign2 = 4'd6; a_sign3 = 4'd12;
b_sign0 = 4'd0; b_sign1 = 4'd0; b_sign2 = 4'd14; b_sign3 = 4'd1;
@(posedge clk_i);
shared_exps0 = 8'd116;
shared_exps1 = 8'd129;
a_mant0 = 8'd84; a_mant1 = 8'd122; a_mant2 = 8'd56; a_mant3 = 8'd157;
b_mant0 = 8'd207; b_mant1 = 8'd226; b_mant2 = 8'd146; b_mant3 = 8'd116;
a_exp0 = 10'd54; a_exp1 = 10'd166; a_exp2 = 10'd564; a_exp3 = 10'd137;
b_exp0 = 10'd111; b_exp1 = 10'd631; b_exp2 = 10'd279; b_exp3 = 10'd756;
a_sign0 = 4'd3; a_sign1 = 4'd5; a_sign2 = 4'd10; a_sign3 = 4'd8;
b_sign0 = 4'd5; b_sign1 = 4'd16; b_sign2 = 4'd3; b_sign3 = 4'd7;
@(posedge clk_i);
a_mant0 = 8'd101; a_mant1 = 8'd214; a_mant2 = 8'd133; a_mant3 = 8'd113;
b_mant0 = 8'd169; b_mant1 = 8'd170; b_mant2 = 8'd24; b_mant3 = 8'd100;
a_exp0 = 10'd314; a_exp1 = 10'd622; a_exp2 = 10'd500; a_exp3 = 10'd608;
b_exp0 = 10'd739; b_exp1 = 10'd1009; b_exp2 = 10'd613; b_exp3 = 10'd603;
a_sign0 = 4'd0; a_sign1 = 4'd3; a_sign2 = 4'd8; a_sign3 = 4'd2;
b_sign0 = 4'd11; b_sign1 = 4'd7; b_sign2 = 4'd1; b_sign3 = 4'd9;
@(posedge clk_i);
a_mant0 = 8'd19; a_mant1 = 8'd43; a_mant2 = 8'd204; a_mant3 = 8'd237;
b_mant0 = 8'd83; b_mant1 = 8'd58; b_mant2 = 8'd91; b_mant3 = 8'd149;
a_exp0 = 10'd315; a_exp1 = 10'd809; a_exp2 = 10'd872; a_exp3 = 10'd958;
b_exp0 = 10'd710; b_exp1 = 10'd575; b_exp2 = 10'd826; b_exp3 = 10'd639;
a_sign0 = 4'd6; a_sign1 = 4'd15; a_sign2 = 4'd8; a_sign3 = 4'd0;
b_sign0 = 4'd7; b_sign1 = 4'd8; b_sign2 = 4'd5; b_sign3 = 4'd13;
@(posedge clk_i);
a_mant0 = 8'd194; a_mant1 = 8'd251; a_mant2 = 8'd115; a_mant3 = 8'd173;
b_mant0 = 8'd235; b_mant1 = 8'd234; b_mant2 = 8'd234; b_mant3 = 8'd92;
a_exp0 = 10'd320; a_exp1 = 10'd428; a_exp2 = 10'd484; a_exp3 = 10'd672;
b_exp0 = 10'd251; b_exp1 = 10'd401; b_exp2 = 10'd771; b_exp3 = 10'd883;
a_sign0 = 4'd15; a_sign1 = 4'd2; a_sign2 = 4'd1; a_sign3 = 4'd14;
b_sign0 = 4'd9; b_sign1 = 4'd11; b_sign2 = 4'd16; b_sign3 = 4'd0;
@(posedge clk_i);
a_mant0 = 8'd169; a_mant1 = 8'd103; a_mant2 = 8'd77; a_mant3 = 8'd121;
b_mant0 = 8'd183; b_mant1 = 8'd166; b_mant2 = 8'd132; b_mant3 = 8'd179;
a_exp0 = 10'd829; a_exp1 = 10'd610; a_exp2 = 10'd427; a_exp3 = 10'd650;
b_exp0 = 10'd929; b_exp1 = 10'd243; b_exp2 = 10'd319; b_exp3 = 10'd71;
a_sign0 = 4'd12; a_sign1 = 4'd13; a_sign2 = 4'd11; a_sign3 = 4'd8;
b_sign0 = 4'd11; b_sign1 = 4'd16; b_sign2 = 4'd7; b_sign3 = 4'd3;
@(posedge clk_i);
a_mant0 = 8'd104; a_mant1 = 8'd158; a_mant2 = 8'd64; a_mant3 = 8'd111;
b_mant0 = 8'd61; b_mant1 = 8'd190; b_mant2 = 8'd95; b_mant3 = 8'd148;
a_exp0 = 10'd191; a_exp1 = 10'd961; a_exp2 = 10'd198; a_exp3 = 10'd463;
b_exp0 = 10'd462; b_exp1 = 10'd850; b_exp2 = 10'd769; b_exp3 = 10'd883;
a_sign0 = 4'd16; a_sign1 = 4'd7; a_sign2 = 4'd4; a_sign3 = 4'd0;
b_sign0 = 4'd8; b_sign1 = 4'd2; b_sign2 = 4'd8; b_sign3 = 4'd10;
@(posedge clk_i);
a_mant0 = 8'd112; a_mant1 = 8'd139; a_mant2 = 8'd223; a_mant3 = 8'd240;
b_mant0 = 8'd37; b_mant1 = 8'd37; b_mant2 = 8'd227; b_mant3 = 8'd170;
a_exp0 = 10'd810; a_exp1 = 10'd368; a_exp2 = 10'd604; a_exp3 = 10'd366;
b_exp0 = 10'd3; b_exp1 = 10'd344; b_exp2 = 10'd415; b_exp3 = 10'd200;
a_sign0 = 4'd6; a_sign1 = 4'd1; a_sign2 = 4'd16; a_sign3 = 4'd8;
b_sign0 = 4'd12; b_sign1 = 4'd4; b_sign2 = 4'd4; b_sign3 = 4'd6;
@(posedge clk_i);
a_mant0 = 8'd152; a_mant1 = 8'd221; a_mant2 = 8'd28; a_mant3 = 8'd54;
b_mant0 = 8'd121; b_mant1 = 8'd40; b_mant2 = 8'd60; b_mant3 = 8'd248;
a_exp0 = 10'd761; a_exp1 = 10'd516; a_exp2 = 10'd288; a_exp3 = 10'd957;
b_exp0 = 10'd648; b_exp1 = 10'd216; b_exp2 = 10'd76; b_exp3 = 10'd678;
a_sign0 = 4'd5; a_sign1 = 4'd1; a_sign2 = 4'd7; a_sign3 = 4'd4;
b_sign0 = 4'd10; b_sign1 = 4'd12; b_sign2 = 4'd14; b_sign3 = 4'd6;
@(posedge clk_i);
shared_exps0 = 8'd130;
shared_exps1 = 8'd112;
a_mant0 = 8'd139; a_mant1 = 8'd4; a_mant2 = 8'd160; a_mant3 = 8'd221;
b_mant0 = 8'd145; b_mant1 = 8'd164; b_mant2 = 8'd55; b_mant3 = 8'd45;
a_exp0 = 10'd217; a_exp1 = 10'd443; a_exp2 = 10'd753; a_exp3 = 10'd134;
b_exp0 = 10'd143; b_exp1 = 10'd973; b_exp2 = 10'd754; b_exp3 = 10'd263;
a_sign0 = 4'd12; a_sign1 = 4'd3; a_sign2 = 4'd1; a_sign3 = 4'd10;
b_sign0 = 4'd11; b_sign1 = 4'd11; b_sign2 = 4'd10; b_sign3 = 4'd3;
@(posedge clk_i);
a_mant0 = 8'd69; a_mant1 = 8'd13; a_mant2 = 8'd217; a_mant3 = 8'd27;
b_mant0 = 8'd207; b_mant1 = 8'd253; b_mant2 = 8'd41; b_mant3 = 8'd253;
a_exp0 = 10'd877; a_exp1 = 10'd857; a_exp2 = 10'd365; a_exp3 = 10'd724;
b_exp0 = 10'd85; b_exp1 = 10'd505; b_exp2 = 10'd312; b_exp3 = 10'd733;
a_sign0 = 4'd8; a_sign1 = 4'd15; a_sign2 = 4'd15; a_sign3 = 4'd2;
b_sign0 = 4'd7; b_sign1 = 4'd15; b_sign2 = 4'd16; b_sign3 = 4'd7;
@(posedge clk_i);
a_mant0 = 8'd49; a_mant1 = 8'd133; a_mant2 = 8'd182; a_mant3 = 8'd134;
b_mant0 = 8'd230; b_mant1 = 8'd116; b_mant2 = 8'd35; b_mant3 = 8'd30;
a_exp0 = 10'd51; a_exp1 = 10'd385; a_exp2 = 10'd38; a_exp3 = 10'd171;
b_exp0 = 10'd360; b_exp1 = 10'd86; b_exp2 = 10'd251; b_exp3 = 10'd14;
a_sign0 = 4'd7; a_sign1 = 4'd8; a_sign2 = 4'd15; a_sign3 = 4'd10;
b_sign0 = 4'd6; b_sign1 = 4'd10; b_sign2 = 4'd10; b_sign3 = 4'd2;
@(posedge clk_i);
a_mant0 = 8'd183; a_mant1 = 8'd174; a_mant2 = 8'd211; a_mant3 = 8'd27;
b_mant0 = 8'd141; b_mant1 = 8'd96; b_mant2 = 8'd223; b_mant3 = 8'd109;
a_exp0 = 10'd584; a_exp1 = 10'd133; a_exp2 = 10'd334; a_exp3 = 10'd117;
b_exp0 = 10'd115; b_exp1 = 10'd281; b_exp2 = 10'd561; b_exp3 = 10'd352;
a_sign0 = 4'd13; a_sign1 = 4'd8; a_sign2 = 4'd3; a_sign3 = 4'd4;
b_sign0 = 4'd2; b_sign1 = 4'd4; b_sign2 = 4'd11; b_sign3 = 4'd10;
@(posedge clk_i);
a_mant0 = 8'd126; a_mant1 = 8'd120; a_mant2 = 8'd200; a_mant3 = 8'd30;
b_mant0 = 8'd54; b_mant1 = 8'd213; b_mant2 = 8'd127; b_mant3 = 8'd68;
a_exp0 = 10'd837; a_exp1 = 10'd457; a_exp2 = 10'd867; a_exp3 = 10'd746;
b_exp0 = 10'd272; b_exp1 = 10'd709; b_exp2 = 10'd329; b_exp3 = 10'd203;
a_sign0 = 4'd14; a_sign1 = 4'd4; a_sign2 = 4'd1; a_sign3 = 4'd3;
b_sign0 = 4'd4; b_sign1 = 4'd5; b_sign2 = 4'd0; b_sign3 = 4'd1;
@(posedge clk_i);
a_mant0 = 8'd124; a_mant1 = 8'd20; a_mant2 = 8'd21; a_mant3 = 8'd207;
b_mant0 = 8'd26; b_mant1 = 8'd133; b_mant2 = 8'd43; b_mant3 = 8'd223;
a_exp0 = 10'd357; a_exp1 = 10'd254; a_exp2 = 10'd358; a_exp3 = 10'd423;
b_exp0 = 10'd744; b_exp1 = 10'd961; b_exp2 = 10'd177; b_exp3 = 10'd663;
a_sign0 = 4'd6; a_sign1 = 4'd10; a_sign2 = 4'd7; a_sign3 = 4'd5;
b_sign0 = 4'd12; b_sign1 = 4'd6; b_sign2 = 4'd7; b_sign3 = 4'd12;
@(posedge clk_i);
a_mant0 = 8'd64; a_mant1 = 8'd98; a_mant2 = 8'd91; a_mant3 = 8'd30;
b_mant0 = 8'd177; b_mant1 = 8'd56; b_mant2 = 8'd63; b_mant3 = 8'd169;
a_exp0 = 10'd310; a_exp1 = 10'd852; a_exp2 = 10'd605; a_exp3 = 10'd290;
b_exp0 = 10'd234; b_exp1 = 10'd529; b_exp2 = 10'd38; b_exp3 = 10'd628;
a_sign0 = 4'd5; a_sign1 = 4'd4; a_sign2 = 4'd13; a_sign3 = 4'd15;
b_sign0 = 4'd0; b_sign1 = 4'd13; b_sign2 = 4'd7; b_sign3 = 4'd0;
@(posedge clk_i);
a_mant0 = 8'd5; a_mant1 = 8'd248; a_mant2 = 8'd180; a_mant3 = 8'd22;
b_mant0 = 8'd42; b_mant1 = 8'd231; b_mant2 = 8'd74; b_mant3 = 8'd77;
a_exp0 = 10'd321; a_exp1 = 10'd67; a_exp2 = 10'd633; a_exp3 = 10'd120;
b_exp0 = 10'd302; b_exp1 = 10'd52; b_exp2 = 10'd40; b_exp3 = 10'd211;
a_sign0 = 4'd16; a_sign1 = 4'd14; a_sign2 = 4'd1; a_sign3 = 4'd15;
b_sign0 = 4'd16; b_sign1 = 4'd5; b_sign2 = 4'd7; b_sign3 = 4'd13;
@(posedge clk_i);
shared_exps0 = 8'd137;
shared_exps1 = 8'd110;
a_mant0 = 8'd161; a_mant1 = 8'd208; a_mant2 = 8'd37; a_mant3 = 8'd160;
b_mant0 = 8'd207; b_mant1 = 8'd213; b_mant2 = 8'd119; b_mant3 = 8'd211;
a_exp0 = 10'd174; a_exp1 = 10'd420; a_exp2 = 10'd282; a_exp3 = 10'd975;
b_exp0 = 10'd942; b_exp1 = 10'd916; b_exp2 = 10'd551; b_exp3 = 10'd529;
a_sign0 = 4'd9; a_sign1 = 4'd12; a_sign2 = 4'd2; a_sign3 = 4'd5;
b_sign0 = 4'd5; b_sign1 = 4'd15; b_sign2 = 4'd2; b_sign3 = 4'd0;
@(posedge clk_i);
a_mant0 = 8'd75; a_mant1 = 8'd155; a_mant2 = 8'd208; a_mant3 = 8'd81;
b_mant0 = 8'd34; b_mant1 = 8'd50; b_mant2 = 8'd30; b_mant3 = 8'd229;
a_exp0 = 10'd206; a_exp1 = 10'd692; a_exp2 = 10'd322; a_exp3 = 10'd636;
b_exp0 = 10'd91; b_exp1 = 10'd903; b_exp2 = 10'd127; b_exp3 = 10'd854;
a_sign0 = 4'd0; a_sign1 = 4'd4; a_sign2 = 4'd15; a_sign3 = 4'd1;
b_sign0 = 4'd16; b_sign1 = 4'd5; b_sign2 = 4'd11; b_sign3 = 4'd2;
@(posedge clk_i);
a_mant0 = 8'd244; a_mant1 = 8'd208; a_mant2 = 8'd15; a_mant3 = 8'd208;
b_mant0 = 8'd244; b_mant1 = 8'd208; b_mant2 = 8'd186; b_mant3 = 8'd112;
a_exp0 = 10'd263; a_exp1 = 10'd999; a_exp2 = 10'd12; a_exp3 = 10'd749;
b_exp0 = 10'd47; b_exp1 = 10'd212; b_exp2 = 10'd171; b_exp3 = 10'd478;
a_sign0 = 4'd9; a_sign1 = 4'd8; a_sign2 = 4'd12; a_sign3 = 4'd11;
b_sign0 = 4'd16; b_sign1 = 4'd16; b_sign2 = 4'd6; b_sign3 = 4'd12;
@(posedge clk_i);
a_mant0 = 8'd231; a_mant1 = 8'd235; a_mant2 = 8'd0; a_mant3 = 8'd131;
b_mant0 = 8'd157; b_mant1 = 8'd47; b_mant2 = 8'd255; b_mant3 = 8'd134;
a_exp0 = 10'd396; a_exp1 = 10'd787; a_exp2 = 10'd876; a_exp3 = 10'd542;
b_exp0 = 10'd1009; b_exp1 = 10'd979; b_exp2 = 10'd375; b_exp3 = 10'd703;
a_sign0 = 4'd9; a_sign1 = 4'd11; a_sign2 = 4'd15; a_sign3 = 4'd16;
b_sign0 = 4'd15; b_sign1 = 4'd14; b_sign2 = 4'd16; b_sign3 = 4'd6;
@(posedge clk_i);
a_mant0 = 8'd120; a_mant1 = 8'd118; a_mant2 = 8'd195; a_mant3 = 8'd14;
b_mant0 = 8'd147; b_mant1 = 8'd58; b_mant2 = 8'd153; b_mant3 = 8'd176;
a_exp0 = 10'd932; a_exp1 = 10'd304; a_exp2 = 10'd312; a_exp3 = 10'd852;
b_exp0 = 10'd949; b_exp1 = 10'd149; b_exp2 = 10'd448; b_exp3 = 10'd115;
a_sign0 = 4'd8; a_sign1 = 4'd4; a_sign2 = 4'd3; a_sign3 = 4'd6;
b_sign0 = 4'd9; b_sign1 = 4'd13; b_sign2 = 4'd11; b_sign3 = 4'd9;
@(posedge clk_i);
a_mant0 = 8'd187; a_mant1 = 8'd46; a_mant2 = 8'd197; a_mant3 = 8'd24;
b_mant0 = 8'd247; b_mant1 = 8'd51; b_mant2 = 8'd37; b_mant3 = 8'd97;
a_exp0 = 10'd320; a_exp1 = 10'd809; a_exp2 = 10'd537; a_exp3 = 10'd723;
b_exp0 = 10'd795; b_exp1 = 10'd212; b_exp2 = 10'd203; b_exp3 = 10'd511;
a_sign0 = 4'd1; a_sign1 = 4'd0; a_sign2 = 4'd0; a_sign3 = 4'd1;
b_sign0 = 4'd6; b_sign1 = 4'd15; b_sign2 = 4'd4; b_sign3 = 4'd5;
@(posedge clk_i);
a_mant0 = 8'd74; a_mant1 = 8'd115; a_mant2 = 8'd34; a_mant3 = 8'd13;
b_mant0 = 8'd245; b_mant1 = 8'd77; b_mant2 = 8'd133; b_mant3 = 8'd202;
a_exp0 = 10'd908; a_exp1 = 10'd227; a_exp2 = 10'd517; a_exp3 = 10'd358;
b_exp0 = 10'd364; b_exp1 = 10'd544; b_exp2 = 10'd938; b_exp3 = 10'd944;
a_sign0 = 4'd4; a_sign1 = 4'd5; a_sign2 = 4'd11; a_sign3 = 4'd2;
b_sign0 = 4'd6; b_sign1 = 4'd6; b_sign2 = 4'd2; b_sign3 = 4'd5;
@(posedge clk_i);
a_mant0 = 8'd128; a_mant1 = 8'd175; a_mant2 = 8'd135; a_mant3 = 8'd129;
b_mant0 = 8'd228; b_mant1 = 8'd143; b_mant2 = 8'd176; b_mant3 = 8'd165;
a_exp0 = 10'd800; a_exp1 = 10'd951; a_exp2 = 10'd771; a_exp3 = 10'd240;
b_exp0 = 10'd844; b_exp1 = 10'd845; b_exp2 = 10'd755; b_exp3 = 10'd1014;
a_sign0 = 4'd0; a_sign1 = 4'd7; a_sign2 = 4'd5; a_sign3 = 4'd11;
b_sign0 = 4'd15; b_sign1 = 4'd4; b_sign2 = 4'd15; b_sign3 = 4'd3;
@(posedge clk_i);
shared_exps0 = 8'd119;
shared_exps1 = 8'd139;
rstn = 0;
@(posedge clk_i);
rstn = 1;
a_mant0 = 8'd82; a_mant1 = 8'd120; a_mant2 = 8'd127; a_mant3 = 8'd71;
b_mant0 = 8'd155; b_mant1 = 8'd57; b_mant2 = 8'd44; b_mant3 = 8'd31;
a_exp0 = 10'd779; a_exp1 = 10'd632; a_exp2 = 10'd453; a_exp3 = 10'd534;
b_exp0 = 10'd327; b_exp1 = 10'd496; b_exp2 = 10'd559; b_exp3 = 10'd143;
a_sign0 = 4'd0; a_sign1 = 4'd16; a_sign2 = 4'd15; a_sign3 = 4'd9;
b_sign0 = 4'd4; b_sign1 = 4'd15; b_sign2 = 4'd8; b_sign3 = 4'd0;
@(posedge clk_i);
a_mant0 = 8'd65; a_mant1 = 8'd234; a_mant2 = 8'd231; a_mant3 = 8'd84;
b_mant0 = 8'd57; b_mant1 = 8'd128; b_mant2 = 8'd20; b_mant3 = 8'd30;
a_exp0 = 10'd716; a_exp1 = 10'd296; a_exp2 = 10'd844; a_exp3 = 10'd856;
b_exp0 = 10'd925; b_exp1 = 10'd358; b_exp2 = 10'd1007; b_exp3 = 10'd180;
a_sign0 = 4'd1; a_sign1 = 4'd13; a_sign2 = 4'd16; a_sign3 = 4'd12;
b_sign0 = 4'd10; b_sign1 = 4'd0; b_sign2 = 4'd1; b_sign3 = 4'd14;
@(posedge clk_i);
a_mant0 = 8'd228; a_mant1 = 8'd41; a_mant2 = 8'd239; a_mant3 = 8'd98;
b_mant0 = 8'd128; b_mant1 = 8'd124; b_mant2 = 8'd221; b_mant3 = 8'd101;
a_exp0 = 10'd1006; a_exp1 = 10'd575; a_exp2 = 10'd341; a_exp3 = 10'd530;
b_exp0 = 10'd50; b_exp1 = 10'd923; b_exp2 = 10'd799; b_exp3 = 10'd202;
a_sign0 = 4'd12; a_sign1 = 4'd9; a_sign2 = 4'd13; a_sign3 = 4'd12;
b_sign0 = 4'd13; b_sign1 = 4'd9; b_sign2 = 4'd5; b_sign3 = 4'd9;
@(posedge clk_i);
a_mant0 = 8'd130; a_mant1 = 8'd86; a_mant2 = 8'd223; a_mant3 = 8'd177;
b_mant0 = 8'd196; b_mant1 = 8'd183; b_mant2 = 8'd200; b_mant3 = 8'd80;
a_exp0 = 10'd35; a_exp1 = 10'd236; a_exp2 = 10'd666; a_exp3 = 10'd545;
b_exp0 = 10'd456; b_exp1 = 10'd926; b_exp2 = 10'd916; b_exp3 = 10'd483;
a_sign0 = 4'd14; a_sign1 = 4'd3; a_sign2 = 4'd14; a_sign3 = 4'd9;
b_sign0 = 4'd1; b_sign1 = 4'd12; b_sign2 = 4'd0; b_sign3 = 4'd15;
@(posedge clk_i);
a_mant0 = 8'd138; a_mant1 = 8'd71; a_mant2 = 8'd21; a_mant3 = 8'd218;
b_mant0 = 8'd237; b_mant1 = 8'd94; b_mant2 = 8'd185; b_mant3 = 8'd142;
a_exp0 = 10'd64; a_exp1 = 10'd525; a_exp2 = 10'd244; a_exp3 = 10'd408;
b_exp0 = 10'd298; b_exp1 = 10'd734; b_exp2 = 10'd157; b_exp3 = 10'd236;
a_sign0 = 4'd9; a_sign1 = 4'd4; a_sign2 = 4'd3; a_sign3 = 4'd9;
b_sign0 = 4'd11; b_sign1 = 4'd1; b_sign2 = 4'd9; b_sign3 = 4'd2;
@(posedge clk_i);
a_mant0 = 8'd178; a_mant1 = 8'd40; a_mant2 = 8'd73; a_mant3 = 8'd226;
b_mant0 = 8'd29; b_mant1 = 8'd154; b_mant2 = 8'd50; b_mant3 = 8'd47;
a_exp0 = 10'd334; a_exp1 = 10'd772; a_exp2 = 10'd250; a_exp3 = 10'd212;
b_exp0 = 10'd564; b_exp1 = 10'd864; b_exp2 = 10'd222; b_exp3 = 10'd844;
a_sign0 = 4'd9; a_sign1 = 4'd14; a_sign2 = 4'd0; a_sign3 = 4'd16;
b_sign0 = 4'd4; b_sign1 = 4'd6; b_sign2 = 4'd5; b_sign3 = 4'd12;
@(posedge clk_i);
a_mant0 = 8'd76; a_mant1 = 8'd177; a_mant2 = 8'd228; a_mant3 = 8'd253;
b_mant0 = 8'd174; b_mant1 = 8'd73; b_mant2 = 8'd85; b_mant3 = 8'd1;
a_exp0 = 10'd164; a_exp1 = 10'd131; a_exp2 = 10'd701; a_exp3 = 10'd187;
b_exp0 = 10'd782; b_exp1 = 10'd990; b_exp2 = 10'd581; b_exp3 = 10'd760;
a_sign0 = 4'd13; a_sign1 = 4'd16; a_sign2 = 4'd3; a_sign3 = 4'd10;
b_sign0 = 4'd7; b_sign1 = 4'd10; b_sign2 = 4'd0; b_sign3 = 4'd3;
@(posedge clk_i);
shared_exps0 = 8'd124;
shared_exps1 = 8'd124;
a_mant0 = 8'd126; a_mant1 = 8'd103; a_mant2 = 8'd145; a_mant3 = 8'd66;
b_mant0 = 8'd113; b_mant1 = 8'd26; b_mant2 = 8'd34; b_mant3 = 8'd44;
a_exp0 = 10'd842; a_exp1 = 10'd810; a_exp2 = 10'd645; a_exp3 = 10'd53;
b_exp0 = 10'd154; b_exp1 = 10'd322; b_exp2 = 10'd641; b_exp3 = 10'd211;
a_sign0 = 4'd7; a_sign1 = 4'd14; a_sign2 = 4'd1; a_sign3 = 4'd2;
b_sign0 = 4'd1; b_sign1 = 4'd14; b_sign2 = 4'd12; b_sign3 = 4'd1;
@(posedge clk_i);
a_mant0 = 8'd33; a_mant1 = 8'd218; a_mant2 = 8'd198; a_mant3 = 8'd78;
b_mant0 = 8'd6; b_mant1 = 8'd37; b_mant2 = 8'd146; b_mant3 = 8'd21;
a_exp0 = 10'd535; a_exp1 = 10'd680; a_exp2 = 10'd741; a_exp3 = 10'd131;
b_exp0 = 10'd579; b_exp1 = 10'd977; b_exp2 = 10'd520; b_exp3 = 10'd959;
a_sign0 = 4'd11; a_sign1 = 4'd5; a_sign2 = 4'd1; a_sign3 = 4'd11;
b_sign0 = 4'd3; b_sign1 = 4'd6; b_sign2 = 4'd10; b_sign3 = 4'd4;
@(posedge clk_i);
a_mant0 = 8'd226; a_mant1 = 8'd45; a_mant2 = 8'd83; a_mant3 = 8'd194;
b_mant0 = 8'd80; b_mant1 = 8'd76; b_mant2 = 8'd0; b_mant3 = 8'd218;
a_exp0 = 10'd127; a_exp1 = 10'd837; a_exp2 = 10'd676; a_exp3 = 10'd333;
b_exp0 = 10'd792; b_exp1 = 10'd477; b_exp2 = 10'd377; b_exp3 = 10'd919;
a_sign0 = 4'd15; a_sign1 = 4'd8; a_sign2 = 4'd11; a_sign3 = 4'd9;
b_sign0 = 4'd15; b_sign1 = 4'd0; b_sign2 = 4'd15; b_sign3 = 4'd2;
@(posedge clk_i);
a_mant0 = 8'd104; a_mant1 = 8'd41; a_mant2 = 8'd178; a_mant3 = 8'd68;
b_mant0 = 8'd225; b_mant1 = 8'd5; b_mant2 = 8'd60; b_mant3 = 8'd94;
a_exp0 = 10'd319; a_exp1 = 10'd270; a_exp2 = 10'd917; a_exp3 = 10'd109;
b_exp0 = 10'd699; b_exp1 = 10'd625; b_exp2 = 10'd1003; b_exp3 = 10'd703;
a_sign0 = 4'd12; a_sign1 = 4'd7; a_sign2 = 4'd8; a_sign3 = 4'd0;
b_sign0 = 4'd15; b_sign1 = 4'd16; b_sign2 = 4'd7; b_sign3 = 4'd1;
@(posedge clk_i);
a_mant0 = 8'd86; a_mant1 = 8'd83; a_mant2 = 8'd63; a_mant3 = 8'd52;
b_mant0 = 8'd12; b_mant1 = 8'd104; b_mant2 = 8'd102; b_mant3 = 8'd34;
a_exp0 = 10'd82; a_exp1 = 10'd331; a_exp2 = 10'd576; a_exp3 = 10'd639;
b_exp0 = 10'd34; b_exp1 = 10'd903; b_exp2 = 10'd222; b_exp3 = 10'd67;
a_sign0 = 4'd14; a_sign1 = 4'd4; a_sign2 = 4'd0; a_sign3 = 4'd12;
b_sign0 = 4'd2; b_sign1 = 4'd13; b_sign2 = 4'd12; b_sign3 = 4'd3;
@(posedge clk_i);
a_mant0 = 8'd111; a_mant1 = 8'd5; a_mant2 = 8'd172; a_mant3 = 8'd114;
b_mant0 = 8'd48; b_mant1 = 8'd218; b_mant2 = 8'd127; b_mant3 = 8'd69;
a_exp0 = 10'd973; a_exp1 = 10'd131; a_exp2 = 10'd68; a_exp3 = 10'd358;
b_exp0 = 10'd805; b_exp1 = 10'd608; b_exp2 = 10'd159; b_exp3 = 10'd608;
a_sign0 = 4'd14; a_sign1 = 4'd12; a_sign2 = 4'd0; a_sign3 = 4'd14;
b_sign0 = 4'd13; b_sign1 = 4'd1; b_sign2 = 4'd12; b_sign3 = 4'd3;
@(posedge clk_i);
a_mant0 = 8'd242; a_mant1 = 8'd30; a_mant2 = 8'd104; a_mant3 = 8'd24;
b_mant0 = 8'd193; b_mant1 = 8'd101; b_mant2 = 8'd89; b_mant3 = 8'd221;
a_exp0 = 10'd824; a_exp1 = 10'd165; a_exp2 = 10'd373; a_exp3 = 10'd923;
b_exp0 = 10'd624; b_exp1 = 10'd101; b_exp2 = 10'd237; b_exp3 = 10'd902;
a_sign0 = 4'd2; a_sign1 = 4'd6; a_sign2 = 4'd11; a_sign3 = 4'd0;
b_sign0 = 4'd6; b_sign1 = 4'd2; b_sign2 = 4'd2; b_sign3 = 4'd15;
@(posedge clk_i);
a_mant0 = 8'd159; a_mant1 = 8'd50; a_mant2 = 8'd121; a_mant3 = 8'd153;
b_mant0 = 8'd202; b_mant1 = 8'd95; b_mant2 = 8'd3; b_mant3 = 8'd81;
a_exp0 = 10'd88; a_exp1 = 10'd634; a_exp2 = 10'd910; a_exp3 = 10'd260;
b_exp0 = 10'd123; b_exp1 = 10'd980; b_exp2 = 10'd904; b_exp3 = 10'd46;
a_sign0 = 4'd1; a_sign1 = 4'd13; a_sign2 = 4'd8; a_sign3 = 4'd6;
b_sign0 = 4'd16; b_sign1 = 4'd15; b_sign2 = 4'd1; b_sign3 = 4'd9;
@(posedge clk_i);
shared_exps0 = 8'd139;
shared_exps1 = 8'd99;
a_mant0 = 8'd112; a_mant1 = 8'd198; a_mant2 = 8'd218; a_mant3 = 8'd252;
b_mant0 = 8'd109; b_mant1 = 8'd7; b_mant2 = 8'd194; b_mant3 = 8'd206;
a_exp0 = 10'd735; a_exp1 = 10'd834; a_exp2 = 10'd717; a_exp3 = 10'd186;
b_exp0 = 10'd693; b_exp1 = 10'd804; b_exp2 = 10'd113; b_exp3 = 10'd528;
a_sign0 = 4'd2; a_sign1 = 4'd5; a_sign2 = 4'd8; a_sign3 = 4'd14;
b_sign0 = 4'd16; b_sign1 = 4'd2; b_sign2 = 4'd3; b_sign3 = 4'd13;
@(posedge clk_i);
a_mant0 = 8'd208; a_mant1 = 8'd36; a_mant2 = 8'd54; a_mant3 = 8'd185;
b_mant0 = 8'd251; b_mant1 = 8'd6; b_mant2 = 8'd67; b_mant3 = 8'd44;
a_exp0 = 10'd331; a_exp1 = 10'd600; a_exp2 = 10'd19; a_exp3 = 10'd598;
b_exp0 = 10'd875; b_exp1 = 10'd457; b_exp2 = 10'd162; b_exp3 = 10'd399;
a_sign0 = 4'd5; a_sign1 = 4'd4; a_sign2 = 4'd11; a_sign3 = 4'd6;
b_sign0 = 4'd4; b_sign1 = 4'd16; b_sign2 = 4'd7; b_sign3 = 4'd6;
@(posedge clk_i);
a_mant0 = 8'd170; a_mant1 = 8'd104; a_mant2 = 8'd152; a_mant3 = 8'd31;
b_mant0 = 8'd116; b_mant1 = 8'd101; b_mant2 = 8'd233; b_mant3 = 8'd138;
a_exp0 = 10'd897; a_exp1 = 10'd860; a_exp2 = 10'd758; a_exp3 = 10'd361;
b_exp0 = 10'd818; b_exp1 = 10'd930; b_exp2 = 10'd86; b_exp3 = 10'd417;
a_sign0 = 4'd3; a_sign1 = 4'd14; a_sign2 = 4'd14; a_sign3 = 4'd12;
b_sign0 = 4'd3; b_sign1 = 4'd9; b_sign2 = 4'd12; b_sign3 = 4'd14;
@(posedge clk_i);
a_mant0 = 8'd212; a_mant1 = 8'd236; a_mant2 = 8'd203; a_mant3 = 8'd236;
b_mant0 = 8'd112; b_mant1 = 8'd88; b_mant2 = 8'd159; b_mant3 = 8'd148;
a_exp0 = 10'd431; a_exp1 = 10'd670; a_exp2 = 10'd899; a_exp3 = 10'd48;
b_exp0 = 10'd259; b_exp1 = 10'd337; b_exp2 = 10'd22; b_exp3 = 10'd101;
a_sign0 = 4'd4; a_sign1 = 4'd1; a_sign2 = 4'd10; a_sign3 = 4'd8;
b_sign0 = 4'd15; b_sign1 = 4'd9; b_sign2 = 4'd7; b_sign3 = 4'd13;
@(posedge clk_i);
a_mant0 = 8'd102; a_mant1 = 8'd27; a_mant2 = 8'd23; a_mant3 = 8'd239;
b_mant0 = 8'd250; b_mant1 = 8'd206; b_mant2 = 8'd249; b_mant3 = 8'd4;
a_exp0 = 10'd575; a_exp1 = 10'd605; a_exp2 = 10'd745; a_exp3 = 10'd403;
b_exp0 = 10'd820; b_exp1 = 10'd276; b_exp2 = 10'd268; b_exp3 = 10'd91;
a_sign0 = 4'd14; a_sign1 = 4'd4; a_sign2 = 4'd9; a_sign3 = 4'd1;
b_sign0 = 4'd7; b_sign1 = 4'd6; b_sign2 = 4'd11; b_sign3 = 4'd3;
@(posedge clk_i);
a_mant0 = 8'd85; a_mant1 = 8'd53; a_mant2 = 8'd202; a_mant3 = 8'd131;
b_mant0 = 8'd204; b_mant1 = 8'd204; b_mant2 = 8'd250; b_mant3 = 8'd216;
a_exp0 = 10'd483; a_exp1 = 10'd925; a_exp2 = 10'd419; a_exp3 = 10'd910;
b_exp0 = 10'd711; b_exp1 = 10'd783; b_exp2 = 10'd645; b_exp3 = 10'd216;
a_sign0 = 4'd3; a_sign1 = 4'd7; a_sign2 = 4'd2; a_sign3 = 4'd9;
b_sign0 = 4'd8; b_sign1 = 4'd16; b_sign2 = 4'd13; b_sign3 = 4'd6;
@(posedge clk_i);
a_mant0 = 8'd27; a_mant1 = 8'd67; a_mant2 = 8'd253; a_mant3 = 8'd113;
b_mant0 = 8'd62; b_mant1 = 8'd154; b_mant2 = 8'd187; b_mant3 = 8'd254;
a_exp0 = 10'd71; a_exp1 = 10'd270; a_exp2 = 10'd374; a_exp3 = 10'd719;
b_exp0 = 10'd681; b_exp1 = 10'd972; b_exp2 = 10'd772; b_exp3 = 10'd1023;
a_sign0 = 4'd12; a_sign1 = 4'd5; a_sign2 = 4'd0; a_sign3 = 4'd14;
b_sign0 = 4'd15; b_sign1 = 4'd5; b_sign2 = 4'd11; b_sign3 = 4'd13;
@(posedge clk_i);
a_mant0 = 8'd79; a_mant1 = 8'd213; a_mant2 = 8'd187; a_mant3 = 8'd253;
b_mant0 = 8'd63; b_mant1 = 8'd160; b_mant2 = 8'd207; b_mant3 = 8'd225;
a_exp0 = 10'd642; a_exp1 = 10'd686; a_exp2 = 10'd695; a_exp3 = 10'd748;
b_exp0 = 10'd28; b_exp1 = 10'd23; b_exp2 = 10'd411; b_exp3 = 10'd863;
a_sign0 = 4'd5; a_sign1 = 4'd13; a_sign2 = 4'd11; a_sign3 = 4'd11;
b_sign0 = 4'd4; b_sign1 = 4'd10; b_sign2 = 4'd15; b_sign3 = 4'd5;
@(posedge clk_i);
shared_exps0 = 8'd119;
shared_exps1 = 8'd142;
a_mant0 = 8'd119; a_mant1 = 8'd103; a_mant2 = 8'd72; a_mant3 = 8'd37;
b_mant0 = 8'd136; b_mant1 = 8'd140; b_mant2 = 8'd121; b_mant3 = 8'd137;
a_exp0 = 10'd654; a_exp1 = 10'd165; a_exp2 = 10'd198; a_exp3 = 10'd927;
b_exp0 = 10'd764; b_exp1 = 10'd420; b_exp2 = 10'd940; b_exp3 = 10'd296;
a_sign0 = 4'd5; a_sign1 = 4'd9; a_sign2 = 4'd10; a_sign3 = 4'd0;
b_sign0 = 4'd9; b_sign1 = 4'd15; b_sign2 = 4'd9; b_sign3 = 4'd5;
@(posedge clk_i);
a_mant0 = 8'd217; a_mant1 = 8'd85; a_mant2 = 8'd9; a_mant3 = 8'd115;
b_mant0 = 8'd109; b_mant1 = 8'd94; b_mant2 = 8'd57; b_mant3 = 8'd117;
a_exp0 = 10'd344; a_exp1 = 10'd651; a_exp2 = 10'd364; a_exp3 = 10'd846;
b_exp0 = 10'd677; b_exp1 = 10'd556; b_exp2 = 10'd377; b_exp3 = 10'd320;
a_sign0 = 4'd8; a_sign1 = 4'd8; a_sign2 = 4'd8; a_sign3 = 4'd1;
b_sign0 = 4'd9; b_sign1 = 4'd4; b_sign2 = 4'd14; b_sign3 = 4'd7;
@(posedge clk_i);
a_mant0 = 8'd90; a_mant1 = 8'd36; a_mant2 = 8'd242; a_mant3 = 8'd148;
b_mant0 = 8'd140; b_mant1 = 8'd162; b_mant2 = 8'd62; b_mant3 = 8'd211;
a_exp0 = 10'd392; a_exp1 = 10'd400; a_exp2 = 10'd653; a_exp3 = 10'd206;
b_exp0 = 10'd200; b_exp1 = 10'd579; b_exp2 = 10'd95; b_exp3 = 10'd411;
a_sign0 = 4'd16; a_sign1 = 4'd3; a_sign2 = 4'd6; a_sign3 = 4'd4;
b_sign0 = 4'd0; b_sign1 = 4'd0; b_sign2 = 4'd15; b_sign3 = 4'd14;
@(posedge clk_i);
a_mant0 = 8'd90; a_mant1 = 8'd202; a_mant2 = 8'd65; a_mant3 = 8'd209;
b_mant0 = 8'd78; b_mant1 = 8'd195; b_mant2 = 8'd18; b_mant3 = 8'd29;
a_exp0 = 10'd637; a_exp1 = 10'd348; a_exp2 = 10'd616; a_exp3 = 10'd550;
b_exp0 = 10'd903; b_exp1 = 10'd898; b_exp2 = 10'd281; b_exp3 = 10'd204;
a_sign0 = 4'd14; a_sign1 = 4'd5; a_sign2 = 4'd1; a_sign3 = 4'd1;
b_sign0 = 4'd4; b_sign1 = 4'd1; b_sign2 = 4'd11; b_sign3 = 4'd8;
@(posedge clk_i);
a_mant0 = 8'd122; a_mant1 = 8'd51; a_mant2 = 8'd239; a_mant3 = 8'd44;
b_mant0 = 8'd0; b_mant1 = 8'd47; b_mant2 = 8'd68; b_mant3 = 8'd130;
a_exp0 = 10'd481; a_exp1 = 10'd670; a_exp2 = 10'd886; a_exp3 = 10'd248;
b_exp0 = 10'd39; b_exp1 = 10'd490; b_exp2 = 10'd99; b_exp3 = 10'd497;
a_sign0 = 4'd14; a_sign1 = 4'd14; a_sign2 = 4'd7; a_sign3 = 4'd4;
b_sign0 = 4'd3; b_sign1 = 4'd1; b_sign2 = 4'd9; b_sign3 = 4'd10;
@(posedge clk_i);
a_mant0 = 8'd63; a_mant1 = 8'd101; a_mant2 = 8'd207; a_mant3 = 8'd148;
b_mant0 = 8'd190; b_mant1 = 8'd199; b_mant2 = 8'd1; b_mant3 = 8'd165;
a_exp0 = 10'd801; a_exp1 = 10'd32; a_exp2 = 10'd1005; a_exp3 = 10'd570;
b_exp0 = 10'd794; b_exp1 = 10'd612; b_exp2 = 10'd917; b_exp3 = 10'd764;
a_sign0 = 4'd0; a_sign1 = 4'd9; a_sign2 = 4'd16; a_sign3 = 4'd8;
b_sign0 = 4'd12; b_sign1 = 4'd14; b_sign2 = 4'd2; b_sign3 = 4'd6;
@(posedge clk_i);
a_mant0 = 8'd210; a_mant1 = 8'd227; a_mant2 = 8'd169; a_mant3 = 8'd106;
b_mant0 = 8'd172; b_mant1 = 8'd3; b_mant2 = 8'd137; b_mant3 = 8'd5;
a_exp0 = 10'd880; a_exp1 = 10'd719; a_exp2 = 10'd947; a_exp3 = 10'd1000;
b_exp0 = 10'd101; b_exp1 = 10'd984; b_exp2 = 10'd83; b_exp3 = 10'd845;
a_sign0 = 4'd13; a_sign1 = 4'd0; a_sign2 = 4'd8; a_sign3 = 4'd5;
b_sign0 = 4'd15; b_sign1 = 4'd12; b_sign2 = 4'd13; b_sign3 = 4'd9;
@(posedge clk_i);
a_mant0 = 8'd160; a_mant1 = 8'd239; a_mant2 = 8'd246; a_mant3 = 8'd145;
b_mant0 = 8'd137; b_mant1 = 8'd99; b_mant2 = 8'd1; b_mant3 = 8'd195;
a_exp0 = 10'd737; a_exp1 = 10'd1010; a_exp2 = 10'd78; a_exp3 = 10'd744;
b_exp0 = 10'd845; b_exp1 = 10'd129; b_exp2 = 10'd148; b_exp3 = 10'd313;
a_sign0 = 4'd10; a_sign1 = 4'd1; a_sign2 = 4'd0; a_sign3 = 4'd14;
b_sign0 = 4'd6; b_sign1 = 4'd14; b_sign2 = 4'd8; b_sign3 = 4'd15;
@(posedge clk_i);
shared_exps0 = 8'd129;
shared_exps1 = 8'd106;
rstn = 0;
@(posedge clk_i);
rstn = 1;
a_mant0 = 8'd98; a_mant1 = 8'd115; a_mant2 = 8'd234; a_mant3 = 8'd27;
b_mant0 = 8'd168; b_mant1 = 8'd73; b_mant2 = 8'd134; b_mant3 = 8'd19;
a_exp0 = 10'd61; a_exp1 = 10'd507; a_exp2 = 10'd665; a_exp3 = 10'd418;
b_exp0 = 10'd96; b_exp1 = 10'd338; b_exp2 = 10'd501; b_exp3 = 10'd662;
a_sign0 = 4'd9; a_sign1 = 4'd15; a_sign2 = 4'd15; a_sign3 = 4'd16;
b_sign0 = 4'd10; b_sign1 = 4'd9; b_sign2 = 4'd8; b_sign3 = 4'd0;
@(posedge clk_i);
a_mant0 = 8'd179; a_mant1 = 8'd62; a_mant2 = 8'd38; a_mant3 = 8'd157;
b_mant0 = 8'd187; b_mant1 = 8'd219; b_mant2 = 8'd126; b_mant3 = 8'd82;
a_exp0 = 10'd234; a_exp1 = 10'd950; a_exp2 = 10'd848; a_exp3 = 10'd169;
b_exp0 = 10'd258; b_exp1 = 10'd644; b_exp2 = 10'd356; b_exp3 = 10'd817;
a_sign0 = 4'd0; a_sign1 = 4'd16; a_sign2 = 4'd12; a_sign3 = 4'd9;
b_sign0 = 4'd10; b_sign1 = 4'd6; b_sign2 = 4'd8; b_sign3 = 4'd9;
@(posedge clk_i);
a_mant0 = 8'd164; a_mant1 = 8'd135; a_mant2 = 8'd214; a_mant3 = 8'd115;
b_mant0 = 8'd228; b_mant1 = 8'd201; b_mant2 = 8'd175; b_mant3 = 8'd69;
a_exp0 = 10'd387; a_exp1 = 10'd708; a_exp2 = 10'd105; a_exp3 = 10'd779;
b_exp0 = 10'd415; b_exp1 = 10'd651; b_exp2 = 10'd182; b_exp3 = 10'd747;
a_sign0 = 4'd8; a_sign1 = 4'd6; a_sign2 = 4'd14; a_sign3 = 4'd9;
b_sign0 = 4'd6; b_sign1 = 4'd11; b_sign2 = 4'd9; b_sign3 = 4'd0;
@(posedge clk_i);
a_mant0 = 8'd158; a_mant1 = 8'd85; a_mant2 = 8'd48; a_mant3 = 8'd154;
b_mant0 = 8'd184; b_mant1 = 8'd114; b_mant2 = 8'd48; b_mant3 = 8'd190;
a_exp0 = 10'd18; a_exp1 = 10'd641; a_exp2 = 10'd913; a_exp3 = 10'd318;
b_exp0 = 10'd389; b_exp1 = 10'd515; b_exp2 = 10'd395; b_exp3 = 10'd156;
a_sign0 = 4'd10; a_sign1 = 4'd16; a_sign2 = 4'd15; a_sign3 = 4'd3;
b_sign0 = 4'd0; b_sign1 = 4'd3; b_sign2 = 4'd11; b_sign3 = 4'd10;
@(posedge clk_i);
a_mant0 = 8'd137; a_mant1 = 8'd154; a_mant2 = 8'd132; a_mant3 = 8'd155;
b_mant0 = 8'd18; b_mant1 = 8'd244; b_mant2 = 8'd193; b_mant3 = 8'd83;
a_exp0 = 10'd734; a_exp1 = 10'd533; a_exp2 = 10'd677; a_exp3 = 10'd505;
b_exp0 = 10'd560; b_exp1 = 10'd708; b_exp2 = 10'd82; b_exp3 = 10'd708;
a_sign0 = 4'd13; a_sign1 = 4'd11; a_sign2 = 4'd13; a_sign3 = 4'd8;
b_sign0 = 4'd15; b_sign1 = 4'd0; b_sign2 = 4'd13; b_sign3 = 4'd5;
@(posedge clk_i);
a_mant0 = 8'd23; a_mant1 = 8'd230; a_mant2 = 8'd27; a_mant3 = 8'd232;
b_mant0 = 8'd126; b_mant1 = 8'd7; b_mant2 = 8'd100; b_mant3 = 8'd186;
a_exp0 = 10'd813; a_exp1 = 10'd251; a_exp2 = 10'd152; a_exp3 = 10'd124;
b_exp0 = 10'd968; b_exp1 = 10'd684; b_exp2 = 10'd766; b_exp3 = 10'd371;
a_sign0 = 4'd9; a_sign1 = 4'd5; a_sign2 = 4'd3; a_sign3 = 4'd15;
b_sign0 = 4'd2; b_sign1 = 4'd14; b_sign2 = 4'd11; b_sign3 = 4'd5;
@(posedge clk_i);
a_mant0 = 8'd249; a_mant1 = 8'd184; a_mant2 = 8'd92; a_mant3 = 8'd43;
b_mant0 = 8'd213; b_mant1 = 8'd24; b_mant2 = 8'd30; b_mant3 = 8'd27;
a_exp0 = 10'd410; a_exp1 = 10'd559; a_exp2 = 10'd951; a_exp3 = 10'd933;
b_exp0 = 10'd880; b_exp1 = 10'd173; b_exp2 = 10'd240; b_exp3 = 10'd955;
a_sign0 = 4'd3; a_sign1 = 4'd6; a_sign2 = 4'd9; a_sign3 = 4'd3;
b_sign0 = 4'd16; b_sign1 = 4'd14; b_sign2 = 4'd2; b_sign3 = 4'd0;
@(posedge clk_i);
shared_exps0 = 8'd155;
shared_exps1 = 8'd120;
a_mant0 = 8'd189; a_mant1 = 8'd239; a_mant2 = 8'd145; a_mant3 = 8'd51;
b_mant0 = 8'd26; b_mant1 = 8'd172; b_mant2 = 8'd171; b_mant3 = 8'd110;
a_exp0 = 10'd838; a_exp1 = 10'd998; a_exp2 = 10'd610; a_exp3 = 10'd922;
b_exp0 = 10'd491; b_exp1 = 10'd138; b_exp2 = 10'd651; b_exp3 = 10'd649;
a_sign0 = 4'd11; a_sign1 = 4'd4; a_sign2 = 4'd4; a_sign3 = 4'd8;
b_sign0 = 4'd12; b_sign1 = 4'd0; b_sign2 = 4'd3; b_sign3 = 4'd1;
@(posedge clk_i);
a_mant0 = 8'd231; a_mant1 = 8'd217; a_mant2 = 8'd43; a_mant3 = 8'd41;
b_mant0 = 8'd50; b_mant1 = 8'd72; b_mant2 = 8'd98; b_mant3 = 8'd121;
a_exp0 = 10'd467; a_exp1 = 10'd643; a_exp2 = 10'd587; a_exp3 = 10'd551;
b_exp0 = 10'd948; b_exp1 = 10'd660; b_exp2 = 10'd597; b_exp3 = 10'd193;
a_sign0 = 4'd9; a_sign1 = 4'd2; a_sign2 = 4'd1; a_sign3 = 4'd13;
b_sign0 = 4'd15; b_sign1 = 4'd3; b_sign2 = 4'd7; b_sign3 = 4'd7;
@(posedge clk_i);
a_mant0 = 8'd135; a_mant1 = 8'd130; a_mant2 = 8'd101; a_mant3 = 8'd123;
b_mant0 = 8'd222; b_mant1 = 8'd138; b_mant2 = 8'd216; b_mant3 = 8'd34;
a_exp0 = 10'd47; a_exp1 = 10'd28; a_exp2 = 10'd766; a_exp3 = 10'd592;
b_exp0 = 10'd496; b_exp1 = 10'd524; b_exp2 = 10'd517; b_exp3 = 10'd786;
a_sign0 = 4'd15; a_sign1 = 4'd3; a_sign2 = 4'd5; a_sign3 = 4'd9;
b_sign0 = 4'd12; b_sign1 = 4'd16; b_sign2 = 4'd12; b_sign3 = 4'd2;
@(posedge clk_i);
a_mant0 = 8'd220; a_mant1 = 8'd186; a_mant2 = 8'd150; a_mant3 = 8'd165;
b_mant0 = 8'd19; b_mant1 = 8'd252; b_mant2 = 8'd54; b_mant3 = 8'd60;
a_exp0 = 10'd508; a_exp1 = 10'd985; a_exp2 = 10'd49; a_exp3 = 10'd724;
b_exp0 = 10'd597; b_exp1 = 10'd174; b_exp2 = 10'd12; b_exp3 = 10'd746;
a_sign0 = 4'd0; a_sign1 = 4'd12; a_sign2 = 4'd1; a_sign3 = 4'd11;
b_sign0 = 4'd14; b_sign1 = 4'd5; b_sign2 = 4'd10; b_sign3 = 4'd11;
@(posedge clk_i);
a_mant0 = 8'd236; a_mant1 = 8'd2; a_mant2 = 8'd164; a_mant3 = 8'd184;
b_mant0 = 8'd99; b_mant1 = 8'd110; b_mant2 = 8'd33; b_mant3 = 8'd53;
a_exp0 = 10'd737; a_exp1 = 10'd181; a_exp2 = 10'd281; a_exp3 = 10'd915;
b_exp0 = 10'd176; b_exp1 = 10'd489; b_exp2 = 10'd280; b_exp3 = 10'd372;
a_sign0 = 4'd16; a_sign1 = 4'd3; a_sign2 = 4'd6; a_sign3 = 4'd16;
b_sign0 = 4'd14; b_sign1 = 4'd9; b_sign2 = 4'd3; b_sign3 = 4'd5;
@(posedge clk_i);
a_mant0 = 8'd105; a_mant1 = 8'd12; a_mant2 = 8'd22; a_mant3 = 8'd113;
b_mant0 = 8'd152; b_mant1 = 8'd173; b_mant2 = 8'd30; b_mant3 = 8'd19;
a_exp0 = 10'd236; a_exp1 = 10'd838; a_exp2 = 10'd227; a_exp3 = 10'd710;
b_exp0 = 10'd879; b_exp1 = 10'd888; b_exp2 = 10'd552; b_exp3 = 10'd180;
a_sign0 = 4'd6; a_sign1 = 4'd16; a_sign2 = 4'd8; a_sign3 = 4'd0;
b_sign0 = 4'd9; b_sign1 = 4'd12; b_sign2 = 4'd0; b_sign3 = 4'd8;
@(posedge clk_i);
a_mant0 = 8'd3; a_mant1 = 8'd150; a_mant2 = 8'd239; a_mant3 = 8'd162;
b_mant0 = 8'd104; b_mant1 = 8'd116; b_mant2 = 8'd123; b_mant3 = 8'd133;
a_exp0 = 10'd309; a_exp1 = 10'd731; a_exp2 = 10'd490; a_exp3 = 10'd509;
b_exp0 = 10'd326; b_exp1 = 10'd34; b_exp2 = 10'd777; b_exp3 = 10'd568;
a_sign0 = 4'd7; a_sign1 = 4'd13; a_sign2 = 4'd1; a_sign3 = 4'd13;
b_sign0 = 4'd16; b_sign1 = 4'd4; b_sign2 = 4'd9; b_sign3 = 4'd12;
@(posedge clk_i);
a_mant0 = 8'd56; a_mant1 = 8'd63; a_mant2 = 8'd54; a_mant3 = 8'd178;
b_mant0 = 8'd243; b_mant1 = 8'd72; b_mant2 = 8'd223; b_mant3 = 8'd238;
a_exp0 = 10'd441; a_exp1 = 10'd567; a_exp2 = 10'd833; a_exp3 = 10'd848;
b_exp0 = 10'd841; b_exp1 = 10'd584; b_exp2 = 10'd540; b_exp3 = 10'd1003;
a_sign0 = 4'd8; a_sign1 = 4'd14; a_sign2 = 4'd2; a_sign3 = 4'd12;
b_sign0 = 4'd3; b_sign1 = 4'd0; b_sign2 = 4'd15; b_sign3 = 4'd9;
@(posedge clk_i);
shared_exps0 = 8'd126;
shared_exps1 = 8'd124;
a_mant0 = 8'd156; a_mant1 = 8'd67; a_mant2 = 8'd115; a_mant3 = 8'd111;
b_mant0 = 8'd228; b_mant1 = 8'd198; b_mant2 = 8'd111; b_mant3 = 8'd135;
a_exp0 = 10'd391; a_exp1 = 10'd665; a_exp2 = 10'd614; a_exp3 = 10'd973;
b_exp0 = 10'd816; b_exp1 = 10'd340; b_exp2 = 10'd685; b_exp3 = 10'd410;
a_sign0 = 4'd13; a_sign1 = 4'd9; a_sign2 = 4'd9; a_sign3 = 4'd13;
b_sign0 = 4'd13; b_sign1 = 4'd3; b_sign2 = 4'd11; b_sign3 = 4'd5;
@(posedge clk_i);
a_mant0 = 8'd202; a_mant1 = 8'd192; a_mant2 = 8'd3; a_mant3 = 8'd239;
b_mant0 = 8'd176; b_mant1 = 8'd154; b_mant2 = 8'd138; b_mant3 = 8'd136;
a_exp0 = 10'd485; a_exp1 = 10'd527; a_exp2 = 10'd872; a_exp3 = 10'd437;
b_exp0 = 10'd371; b_exp1 = 10'd580; b_exp2 = 10'd709; b_exp3 = 10'd748;
a_sign0 = 4'd8; a_sign1 = 4'd7; a_sign2 = 4'd14; a_sign3 = 4'd10;
b_sign0 = 4'd14; b_sign1 = 4'd3; b_sign2 = 4'd2; b_sign3 = 4'd14;
@(posedge clk_i);
a_mant0 = 8'd27; a_mant1 = 8'd86; a_mant2 = 8'd105; a_mant3 = 8'd83;
b_mant0 = 8'd53; b_mant1 = 8'd108; b_mant2 = 8'd46; b_mant3 = 8'd199;
a_exp0 = 10'd170; a_exp1 = 10'd864; a_exp2 = 10'd423; a_exp3 = 10'd773;
b_exp0 = 10'd435; b_exp1 = 10'd863; b_exp2 = 10'd77; b_exp3 = 10'd742;
a_sign0 = 4'd3; a_sign1 = 4'd15; a_sign2 = 4'd10; a_sign3 = 4'd1;
b_sign0 = 4'd15; b_sign1 = 4'd16; b_sign2 = 4'd15; b_sign3 = 4'd0;
@(posedge clk_i);
a_mant0 = 8'd121; a_mant1 = 8'd34; a_mant2 = 8'd194; a_mant3 = 8'd211;
b_mant0 = 8'd145; b_mant1 = 8'd83; b_mant2 = 8'd66; b_mant3 = 8'd230;
a_exp0 = 10'd477; a_exp1 = 10'd911; a_exp2 = 10'd387; a_exp3 = 10'd151;
b_exp0 = 10'd116; b_exp1 = 10'd140; b_exp2 = 10'd1006; b_exp3 = 10'd818;
a_sign0 = 4'd5; a_sign1 = 4'd0; a_sign2 = 4'd13; a_sign3 = 4'd13;
b_sign0 = 4'd5; b_sign1 = 4'd3; b_sign2 = 4'd9; b_sign3 = 4'd11;
@(posedge clk_i);
a_mant0 = 8'd115; a_mant1 = 8'd233; a_mant2 = 8'd55; a_mant3 = 8'd194;
b_mant0 = 8'd52; b_mant1 = 8'd85; b_mant2 = 8'd235; b_mant3 = 8'd133;
a_exp0 = 10'd116; a_exp1 = 10'd476; a_exp2 = 10'd339; a_exp3 = 10'd260;
b_exp0 = 10'd768; b_exp1 = 10'd71; b_exp2 = 10'd180; b_exp3 = 10'd305;
a_sign0 = 4'd0; a_sign1 = 4'd3; a_sign2 = 4'd11; a_sign3 = 4'd7;
b_sign0 = 4'd8; b_sign1 = 4'd7; b_sign2 = 4'd2; b_sign3 = 4'd3;
@(posedge clk_i);
a_mant0 = 8'd131; a_mant1 = 8'd2; a_mant2 = 8'd236; a_mant3 = 8'd3;
b_mant0 = 8'd197; b_mant1 = 8'd164; b_mant2 = 8'd169; b_mant3 = 8'd79;
a_exp0 = 10'd727; a_exp1 = 10'd756; a_exp2 = 10'd750; a_exp3 = 10'd792;
b_exp0 = 10'd826; b_exp1 = 10'd728; b_exp2 = 10'd136; b_exp3 = 10'd936;
a_sign0 = 4'd3; a_sign1 = 4'd2; a_sign2 = 4'd7; a_sign3 = 4'd12;
b_sign0 = 4'd8; b_sign1 = 4'd3; b_sign2 = 4'd9; b_sign3 = 4'd9;
@(posedge clk_i);
a_mant0 = 8'd12; a_mant1 = 8'd182; a_mant2 = 8'd44; a_mant3 = 8'd30;
b_mant0 = 8'd231; b_mant1 = 8'd165; b_mant2 = 8'd174; b_mant3 = 8'd70;
a_exp0 = 10'd325; a_exp1 = 10'd970; a_exp2 = 10'd475; a_exp3 = 10'd824;
b_exp0 = 10'd814; b_exp1 = 10'd641; b_exp2 = 10'd404; b_exp3 = 10'd357;
a_sign0 = 4'd9; a_sign1 = 4'd11; a_sign2 = 4'd15; a_sign3 = 4'd6;
b_sign0 = 4'd3; b_sign1 = 4'd3; b_sign2 = 4'd11; b_sign3 = 4'd10;
@(posedge clk_i);
a_mant0 = 8'd255; a_mant1 = 8'd99; a_mant2 = 8'd20; a_mant3 = 8'd21;
b_mant0 = 8'd174; b_mant1 = 8'd153; b_mant2 = 8'd130; b_mant3 = 8'd63;
a_exp0 = 10'd970; a_exp1 = 10'd251; a_exp2 = 10'd692; a_exp3 = 10'd33;
b_exp0 = 10'd154; b_exp1 = 10'd868; b_exp2 = 10'd379; b_exp3 = 10'd871;
a_sign0 = 4'd15; a_sign1 = 4'd16; a_sign2 = 4'd7; a_sign3 = 4'd1;
b_sign0 = 4'd3; b_sign1 = 4'd3; b_sign2 = 4'd15; b_sign3 = 4'd14;
@(posedge clk_i);
shared_exps0 = 8'd123;
shared_exps1 = 8'd107;
a_mant0 = 8'd207; a_mant1 = 8'd104; a_mant2 = 8'd140; a_mant3 = 8'd184;
b_mant0 = 8'd133; b_mant1 = 8'd40; b_mant2 = 8'd110; b_mant3 = 8'd229;
a_exp0 = 10'd64; a_exp1 = 10'd807; a_exp2 = 10'd978; a_exp3 = 10'd748;
b_exp0 = 10'd910; b_exp1 = 10'd376; b_exp2 = 10'd811; b_exp3 = 10'd584;
a_sign0 = 4'd7; a_sign1 = 4'd7; a_sign2 = 4'd16; a_sign3 = 4'd7;
b_sign0 = 4'd15; b_sign1 = 4'd1; b_sign2 = 4'd11; b_sign3 = 4'd12;
@(posedge clk_i);
a_mant0 = 8'd102; a_mant1 = 8'd167; a_mant2 = 8'd202; a_mant3 = 8'd246;
b_mant0 = 8'd21; b_mant1 = 8'd253; b_mant2 = 8'd237; b_mant3 = 8'd37;
a_exp0 = 10'd635; a_exp1 = 10'd606; a_exp2 = 10'd318; a_exp3 = 10'd226;
b_exp0 = 10'd485; b_exp1 = 10'd704; b_exp2 = 10'd301; b_exp3 = 10'd743;
a_sign0 = 4'd14; a_sign1 = 4'd9; a_sign2 = 4'd1; a_sign3 = 4'd15;
b_sign0 = 4'd16; b_sign1 = 4'd14; b_sign2 = 4'd0; b_sign3 = 4'd13;
@(posedge clk_i);
a_mant0 = 8'd227; a_mant1 = 8'd205; a_mant2 = 8'd108; a_mant3 = 8'd218;
b_mant0 = 8'd169; b_mant1 = 8'd80; b_mant2 = 8'd138; b_mant3 = 8'd145;
a_exp0 = 10'd347; a_exp1 = 10'd707; a_exp2 = 10'd719; a_exp3 = 10'd491;
b_exp0 = 10'd641; b_exp1 = 10'd55; b_exp2 = 10'd799; b_exp3 = 10'd749;
a_sign0 = 4'd7; a_sign1 = 4'd8; a_sign2 = 4'd14; a_sign3 = 4'd11;
b_sign0 = 4'd4; b_sign1 = 4'd0; b_sign2 = 4'd6; b_sign3 = 4'd1;
@(posedge clk_i);
a_mant0 = 8'd208; a_mant1 = 8'd148; a_mant2 = 8'd253; a_mant3 = 8'd225;
b_mant0 = 8'd103; b_mant1 = 8'd53; b_mant2 = 8'd188; b_mant3 = 8'd247;
a_exp0 = 10'd715; a_exp1 = 10'd424; a_exp2 = 10'd790; a_exp3 = 10'd464;
b_exp0 = 10'd335; b_exp1 = 10'd167; b_exp2 = 10'd877; b_exp3 = 10'd195;
a_sign0 = 4'd1; a_sign1 = 4'd6; a_sign2 = 4'd13; a_sign3 = 4'd5;
b_sign0 = 4'd12; b_sign1 = 4'd12; b_sign2 = 4'd14; b_sign3 = 4'd12;
@(posedge clk_i);
a_mant0 = 8'd153; a_mant1 = 8'd11; a_mant2 = 8'd153; a_mant3 = 8'd6;
b_mant0 = 8'd142; b_mant1 = 8'd173; b_mant2 = 8'd35; b_mant3 = 8'd17;
a_exp0 = 10'd840; a_exp1 = 10'd567; a_exp2 = 10'd258; a_exp3 = 10'd862;
b_exp0 = 10'd364; b_exp1 = 10'd415; b_exp2 = 10'd506; b_exp3 = 10'd838;
a_sign0 = 4'd0; a_sign1 = 4'd8; a_sign2 = 4'd10; a_sign3 = 4'd1;
b_sign0 = 4'd12; b_sign1 = 4'd1; b_sign2 = 4'd8; b_sign3 = 4'd12;
@(posedge clk_i);
a_mant0 = 8'd164; a_mant1 = 8'd202; a_mant2 = 8'd197; a_mant3 = 8'd237;
b_mant0 = 8'd177; b_mant1 = 8'd108; b_mant2 = 8'd165; b_mant3 = 8'd61;
a_exp0 = 10'd977; a_exp1 = 10'd1009; a_exp2 = 10'd203; a_exp3 = 10'd0;
b_exp0 = 10'd699; b_exp1 = 10'd67; b_exp2 = 10'd372; b_exp3 = 10'd232;
a_sign0 = 4'd7; a_sign1 = 4'd16; a_sign2 = 4'd4; a_sign3 = 4'd2;
b_sign0 = 4'd11; b_sign1 = 4'd6; b_sign2 = 4'd11; b_sign3 = 4'd10;
@(posedge clk_i);
a_mant0 = 8'd115; a_mant1 = 8'd118; a_mant2 = 8'd209; a_mant3 = 8'd75;
b_mant0 = 8'd136; b_mant1 = 8'd8; b_mant2 = 8'd14; b_mant3 = 8'd10;
a_exp0 = 10'd327; a_exp1 = 10'd383; a_exp2 = 10'd265; a_exp3 = 10'd412;
b_exp0 = 10'd392; b_exp1 = 10'd308; b_exp2 = 10'd438; b_exp3 = 10'd874;
a_sign0 = 4'd8; a_sign1 = 4'd16; a_sign2 = 4'd4; a_sign3 = 4'd10;
b_sign0 = 4'd8; b_sign1 = 4'd0; b_sign2 = 4'd15; b_sign3 = 4'd9;
@(posedge clk_i);
a_mant0 = 8'd85; a_mant1 = 8'd211; a_mant2 = 8'd16; a_mant3 = 8'd246;
b_mant0 = 8'd181; b_mant1 = 8'd216; b_mant2 = 8'd127; b_mant3 = 8'd21;
a_exp0 = 10'd64; a_exp1 = 10'd605; a_exp2 = 10'd540; a_exp3 = 10'd325;
b_exp0 = 10'd144; b_exp1 = 10'd240; b_exp2 = 10'd668; b_exp3 = 10'd376;
a_sign0 = 4'd12; a_sign1 = 4'd5; a_sign2 = 4'd5; a_sign3 = 4'd7;
b_sign0 = 4'd3; b_sign1 = 4'd6; b_sign2 = 4'd2; b_sign3 = 4'd14;
@(posedge clk_i);
shared_exps0 = 8'd131;
shared_exps1 = 8'd132;
rstn = 0;
@(posedge clk_i);
rstn = 1;
a_mant0 = 8'd69; a_mant1 = 8'd154; a_mant2 = 8'd29; a_mant3 = 8'd110;
b_mant0 = 8'd223; b_mant1 = 8'd166; b_mant2 = 8'd173; b_mant3 = 8'd9;
a_exp0 = 10'd194; a_exp1 = 10'd640; a_exp2 = 10'd609; a_exp3 = 10'd873;
b_exp0 = 10'd702; b_exp1 = 10'd193; b_exp2 = 10'd592; b_exp3 = 10'd447;
a_sign0 = 4'd5; a_sign1 = 4'd0; a_sign2 = 4'd2; a_sign3 = 4'd6;
b_sign0 = 4'd12; b_sign1 = 4'd12; b_sign2 = 4'd13; b_sign3 = 4'd3;
@(posedge clk_i);
a_mant0 = 8'd199; a_mant1 = 8'd140; a_mant2 = 8'd234; a_mant3 = 8'd87;
b_mant0 = 8'd162; b_mant1 = 8'd217; b_mant2 = 8'd157; b_mant3 = 8'd168;
a_exp0 = 10'd536; a_exp1 = 10'd406; a_exp2 = 10'd960; a_exp3 = 10'd230;
b_exp0 = 10'd601; b_exp1 = 10'd605; b_exp2 = 10'd358; b_exp3 = 10'd638;
a_sign0 = 4'd14; a_sign1 = 4'd10; a_sign2 = 4'd14; a_sign3 = 4'd14;
b_sign0 = 4'd5; b_sign1 = 4'd2; b_sign2 = 4'd15; b_sign3 = 4'd4;
@(posedge clk_i);
a_mant0 = 8'd221; a_mant1 = 8'd93; a_mant2 = 8'd149; a_mant3 = 8'd208;
b_mant0 = 8'd111; b_mant1 = 8'd25; b_mant2 = 8'd103; b_mant3 = 8'd216;
a_exp0 = 10'd214; a_exp1 = 10'd296; a_exp2 = 10'd828; a_exp3 = 10'd119;
b_exp0 = 10'd775; b_exp1 = 10'd877; b_exp2 = 10'd640; b_exp3 = 10'd441;
a_sign0 = 4'd5; a_sign1 = 4'd8; a_sign2 = 4'd3; a_sign3 = 4'd9;
b_sign0 = 4'd6; b_sign1 = 4'd1; b_sign2 = 4'd12; b_sign3 = 4'd15;
@(posedge clk_i);
a_mant0 = 8'd155; a_mant1 = 8'd8; a_mant2 = 8'd180; a_mant3 = 8'd38;
b_mant0 = 8'd177; b_mant1 = 8'd190; b_mant2 = 8'd69; b_mant3 = 8'd102;
a_exp0 = 10'd800; a_exp1 = 10'd876; a_exp2 = 10'd872; a_exp3 = 10'd295;
b_exp0 = 10'd38; b_exp1 = 10'd464; b_exp2 = 10'd788; b_exp3 = 10'd909;
a_sign0 = 4'd15; a_sign1 = 4'd3; a_sign2 = 4'd7; a_sign3 = 4'd8;
b_sign0 = 4'd11; b_sign1 = 4'd12; b_sign2 = 4'd14; b_sign3 = 4'd13;
@(posedge clk_i);
a_mant0 = 8'd25; a_mant1 = 8'd53; a_mant2 = 8'd173; a_mant3 = 8'd197;
b_mant0 = 8'd144; b_mant1 = 8'd90; b_mant2 = 8'd49; b_mant3 = 8'd70;
a_exp0 = 10'd790; a_exp1 = 10'd676; a_exp2 = 10'd693; a_exp3 = 10'd442;
b_exp0 = 10'd489; b_exp1 = 10'd889; b_exp2 = 10'd441; b_exp3 = 10'd826;
a_sign0 = 4'd14; a_sign1 = 4'd12; a_sign2 = 4'd16; a_sign3 = 4'd4;
b_sign0 = 4'd16; b_sign1 = 4'd16; b_sign2 = 4'd8; b_sign3 = 4'd6;
@(posedge clk_i);
a_mant0 = 8'd88; a_mant1 = 8'd59; a_mant2 = 8'd46; a_mant3 = 8'd185;
b_mant0 = 8'd184; b_mant1 = 8'd183; b_mant2 = 8'd128; b_mant3 = 8'd29;
a_exp0 = 10'd87; a_exp1 = 10'd985; a_exp2 = 10'd322; a_exp3 = 10'd598;
b_exp0 = 10'd257; b_exp1 = 10'd677; b_exp2 = 10'd615; b_exp3 = 10'd168;
a_sign0 = 4'd3; a_sign1 = 4'd12; a_sign2 = 4'd13; a_sign3 = 4'd12;
b_sign0 = 4'd1; b_sign1 = 4'd10; b_sign2 = 4'd16; b_sign3 = 4'd4;
@(posedge clk_i);
a_mant0 = 8'd254; a_mant1 = 8'd12; a_mant2 = 8'd118; a_mant3 = 8'd185;
b_mant0 = 8'd29; b_mant1 = 8'd144; b_mant2 = 8'd238; b_mant3 = 8'd112;
a_exp0 = 10'd710; a_exp1 = 10'd180; a_exp2 = 10'd126; a_exp3 = 10'd187;
b_exp0 = 10'd52; b_exp1 = 10'd608; b_exp2 = 10'd796; b_exp3 = 10'd601;
a_sign0 = 4'd0; a_sign1 = 4'd8; a_sign2 = 4'd9; a_sign3 = 4'd7;
b_sign0 = 4'd4; b_sign1 = 4'd4; b_sign2 = 4'd1; b_sign3 = 4'd5;
@(posedge clk_i);
shared_exps0 = 8'd113;
shared_exps1 = 8'd132;
a_mant0 = 8'd33; a_mant1 = 8'd156; a_mant2 = 8'd17; a_mant3 = 8'd2;
b_mant0 = 8'd103; b_mant1 = 8'd99; b_mant2 = 8'd220; b_mant3 = 8'd240;
a_exp0 = 10'd919; a_exp1 = 10'd962; a_exp2 = 10'd818; a_exp3 = 10'd843;
b_exp0 = 10'd478; b_exp1 = 10'd801; b_exp2 = 10'd946; b_exp3 = 10'd957;
a_sign0 = 4'd2; a_sign1 = 4'd5; a_sign2 = 4'd8; a_sign3 = 4'd16;
b_sign0 = 4'd2; b_sign1 = 4'd13; b_sign2 = 4'd10; b_sign3 = 4'd5;
@(posedge clk_i);
a_mant0 = 8'd210; a_mant1 = 8'd235; a_mant2 = 8'd63; a_mant3 = 8'd47;
b_mant0 = 8'd229; b_mant1 = 8'd22; b_mant2 = 8'd10; b_mant3 = 8'd115;
a_exp0 = 10'd761; a_exp1 = 10'd929; a_exp2 = 10'd684; a_exp3 = 10'd804;
b_exp0 = 10'd588; b_exp1 = 10'd232; b_exp2 = 10'd752; b_exp3 = 10'd579;
a_sign0 = 4'd12; a_sign1 = 4'd12; a_sign2 = 4'd6; a_sign3 = 4'd16;
b_sign0 = 4'd1; b_sign1 = 4'd7; b_sign2 = 4'd0; b_sign3 = 4'd16;
@(posedge clk_i);
a_mant0 = 8'd15; a_mant1 = 8'd195; a_mant2 = 8'd118; a_mant3 = 8'd237;
b_mant0 = 8'd132; b_mant1 = 8'd73; b_mant2 = 8'd61; b_mant3 = 8'd28;
a_exp0 = 10'd417; a_exp1 = 10'd903; a_exp2 = 10'd245; a_exp3 = 10'd220;
b_exp0 = 10'd975; b_exp1 = 10'd818; b_exp2 = 10'd820; b_exp3 = 10'd905;
a_sign0 = 4'd9; a_sign1 = 4'd15; a_sign2 = 4'd15; a_sign3 = 4'd7;
b_sign0 = 4'd0; b_sign1 = 4'd6; b_sign2 = 4'd2; b_sign3 = 4'd7;
@(posedge clk_i);
a_mant0 = 8'd209; a_mant1 = 8'd224; a_mant2 = 8'd191; a_mant3 = 8'd183;
b_mant0 = 8'd64; b_mant1 = 8'd82; b_mant2 = 8'd193; b_mant3 = 8'd73;
a_exp0 = 10'd527; a_exp1 = 10'd619; a_exp2 = 10'd171; a_exp3 = 10'd939;
b_exp0 = 10'd141; b_exp1 = 10'd61; b_exp2 = 10'd876; b_exp3 = 10'd182;
a_sign0 = 4'd4; a_sign1 = 4'd5; a_sign2 = 4'd11; a_sign3 = 4'd11;
b_sign0 = 4'd14; b_sign1 = 4'd2; b_sign2 = 4'd10; b_sign3 = 4'd2;
@(posedge clk_i);
a_mant0 = 8'd66; a_mant1 = 8'd189; a_mant2 = 8'd230; a_mant3 = 8'd141;
b_mant0 = 8'd160; b_mant1 = 8'd46; b_mant2 = 8'd190; b_mant3 = 8'd123;
a_exp0 = 10'd71; a_exp1 = 10'd228; a_exp2 = 10'd823; a_exp3 = 10'd685;
b_exp0 = 10'd183; b_exp1 = 10'd347; b_exp2 = 10'd626; b_exp3 = 10'd726;
a_sign0 = 4'd0; a_sign1 = 4'd3; a_sign2 = 4'd14; a_sign3 = 4'd2;
b_sign0 = 4'd5; b_sign1 = 4'd15; b_sign2 = 4'd12; b_sign3 = 4'd4;
@(posedge clk_i);
a_mant0 = 8'd131; a_mant1 = 8'd130; a_mant2 = 8'd4; a_mant3 = 8'd167;
b_mant0 = 8'd35; b_mant1 = 8'd162; b_mant2 = 8'd156; b_mant3 = 8'd117;
a_exp0 = 10'd687; a_exp1 = 10'd1019; a_exp2 = 10'd177; a_exp3 = 10'd978;
b_exp0 = 10'd462; b_exp1 = 10'd715; b_exp2 = 10'd905; b_exp3 = 10'd990;
a_sign0 = 4'd7; a_sign1 = 4'd2; a_sign2 = 4'd12; a_sign3 = 4'd7;
b_sign0 = 4'd10; b_sign1 = 4'd3; b_sign2 = 4'd6; b_sign3 = 4'd11;
@(posedge clk_i);
a_mant0 = 8'd153; a_mant1 = 8'd170; a_mant2 = 8'd204; a_mant3 = 8'd33;
b_mant0 = 8'd142; b_mant1 = 8'd47; b_mant2 = 8'd19; b_mant3 = 8'd183;
a_exp0 = 10'd12; a_exp1 = 10'd981; a_exp2 = 10'd130; a_exp3 = 10'd981;
b_exp0 = 10'd531; b_exp1 = 10'd286; b_exp2 = 10'd704; b_exp3 = 10'd748;
a_sign0 = 4'd12; a_sign1 = 4'd16; a_sign2 = 4'd9; a_sign3 = 4'd3;
b_sign0 = 4'd1; b_sign1 = 4'd14; b_sign2 = 4'd14; b_sign3 = 4'd7;
@(posedge clk_i);
a_mant0 = 8'd226; a_mant1 = 8'd121; a_mant2 = 8'd65; a_mant3 = 8'd20;
b_mant0 = 8'd189; b_mant1 = 8'd59; b_mant2 = 8'd180; b_mant3 = 8'd66;
a_exp0 = 10'd889; a_exp1 = 10'd53; a_exp2 = 10'd528; a_exp3 = 10'd757;
b_exp0 = 10'd805; b_exp1 = 10'd174; b_exp2 = 10'd562; b_exp3 = 10'd127;
a_sign0 = 4'd3; a_sign1 = 4'd8; a_sign2 = 4'd1; a_sign3 = 4'd3;
b_sign0 = 4'd9; b_sign1 = 4'd16; b_sign2 = 4'd15; b_sign3 = 4'd6;
@(posedge clk_i);
shared_exps0 = 8'd133;
shared_exps1 = 8'd108;
a_mant0 = 8'd178; a_mant1 = 8'd237; a_mant2 = 8'd246; a_mant3 = 8'd104;
b_mant0 = 8'd21; b_mant1 = 8'd47; b_mant2 = 8'd202; b_mant3 = 8'd48;
a_exp0 = 10'd239; a_exp1 = 10'd404; a_exp2 = 10'd532; a_exp3 = 10'd278;
b_exp0 = 10'd88; b_exp1 = 10'd706; b_exp2 = 10'd304; b_exp3 = 10'd705;
a_sign0 = 4'd0; a_sign1 = 4'd9; a_sign2 = 4'd11; a_sign3 = 4'd12;
b_sign0 = 4'd14; b_sign1 = 4'd4; b_sign2 = 4'd8; b_sign3 = 4'd13;
@(posedge clk_i);
a_mant0 = 8'd210; a_mant1 = 8'd237; a_mant2 = 8'd51; a_mant3 = 8'd126;
b_mant0 = 8'd184; b_mant1 = 8'd162; b_mant2 = 8'd122; b_mant3 = 8'd246;
a_exp0 = 10'd83; a_exp1 = 10'd167; a_exp2 = 10'd877; a_exp3 = 10'd370;
b_exp0 = 10'd621; b_exp1 = 10'd646; b_exp2 = 10'd616; b_exp3 = 10'd1007;
a_sign0 = 4'd9; a_sign1 = 4'd1; a_sign2 = 4'd15; a_sign3 = 4'd14;
b_sign0 = 4'd13; b_sign1 = 4'd11; b_sign2 = 4'd15; b_sign3 = 4'd14;
@(posedge clk_i);
a_mant0 = 8'd36; a_mant1 = 8'd48; a_mant2 = 8'd219; a_mant3 = 8'd91;
b_mant0 = 8'd161; b_mant1 = 8'd29; b_mant2 = 8'd108; b_mant3 = 8'd223;
a_exp0 = 10'd124; a_exp1 = 10'd749; a_exp2 = 10'd173; a_exp3 = 10'd902;
b_exp0 = 10'd534; b_exp1 = 10'd32; b_exp2 = 10'd362; b_exp3 = 10'd288;
a_sign0 = 4'd13; a_sign1 = 4'd3; a_sign2 = 4'd10; a_sign3 = 4'd0;
b_sign0 = 4'd15; b_sign1 = 4'd10; b_sign2 = 4'd9; b_sign3 = 4'd7;
@(posedge clk_i);
a_mant0 = 8'd44; a_mant1 = 8'd94; a_mant2 = 8'd246; a_mant3 = 8'd163;
b_mant0 = 8'd107; b_mant1 = 8'd221; b_mant2 = 8'd101; b_mant3 = 8'd25;
a_exp0 = 10'd813; a_exp1 = 10'd754; a_exp2 = 10'd51; a_exp3 = 10'd917;
b_exp0 = 10'd217; b_exp1 = 10'd971; b_exp2 = 10'd710; b_exp3 = 10'd125;
a_sign0 = 4'd1; a_sign1 = 4'd8; a_sign2 = 4'd3; a_sign3 = 4'd15;
b_sign0 = 4'd11; b_sign1 = 4'd6; b_sign2 = 4'd1; b_sign3 = 4'd15;
@(posedge clk_i);
a_mant0 = 8'd59; a_mant1 = 8'd79; a_mant2 = 8'd4; a_mant3 = 8'd41;
b_mant0 = 8'd219; b_mant1 = 8'd182; b_mant2 = 8'd230; b_mant3 = 8'd24;
a_exp0 = 10'd71; a_exp1 = 10'd447; a_exp2 = 10'd443; a_exp3 = 10'd626;
b_exp0 = 10'd268; b_exp1 = 10'd497; b_exp2 = 10'd325; b_exp3 = 10'd548;
a_sign0 = 4'd0; a_sign1 = 4'd7; a_sign2 = 4'd1; a_sign3 = 4'd11;
b_sign0 = 4'd9; b_sign1 = 4'd1; b_sign2 = 4'd14; b_sign3 = 4'd13;
@(posedge clk_i);
a_mant0 = 8'd33; a_mant1 = 8'd223; a_mant2 = 8'd204; a_mant3 = 8'd37;
b_mant0 = 8'd3; b_mant1 = 8'd122; b_mant2 = 8'd187; b_mant3 = 8'd33;
a_exp0 = 10'd962; a_exp1 = 10'd3; a_exp2 = 10'd148; a_exp3 = 10'd770;
b_exp0 = 10'd462; b_exp1 = 10'd419; b_exp2 = 10'd326; b_exp3 = 10'd237;
a_sign0 = 4'd15; a_sign1 = 4'd3; a_sign2 = 4'd14; a_sign3 = 4'd12;
b_sign0 = 4'd3; b_sign1 = 4'd7; b_sign2 = 4'd3; b_sign3 = 4'd7;
@(posedge clk_i);
a_mant0 = 8'd212; a_mant1 = 8'd51; a_mant2 = 8'd205; a_mant3 = 8'd172;
b_mant0 = 8'd82; b_mant1 = 8'd73; b_mant2 = 8'd138; b_mant3 = 8'd55;
a_exp0 = 10'd99; a_exp1 = 10'd901; a_exp2 = 10'd556; a_exp3 = 10'd849;
b_exp0 = 10'd631; b_exp1 = 10'd575; b_exp2 = 10'd478; b_exp3 = 10'd882;
a_sign0 = 4'd6; a_sign1 = 4'd0; a_sign2 = 4'd4; a_sign3 = 4'd6;
b_sign0 = 4'd12; b_sign1 = 4'd9; b_sign2 = 4'd15; b_sign3 = 4'd5;
@(posedge clk_i);
a_mant0 = 8'd46; a_mant1 = 8'd55; a_mant2 = 8'd202; a_mant3 = 8'd248;
b_mant0 = 8'd106; b_mant1 = 8'd177; b_mant2 = 8'd227; b_mant3 = 8'd249;
a_exp0 = 10'd885; a_exp1 = 10'd321; a_exp2 = 10'd397; a_exp3 = 10'd54;
b_exp0 = 10'd489; b_exp1 = 10'd498; b_exp2 = 10'd429; b_exp3 = 10'd606;
a_sign0 = 4'd11; a_sign1 = 4'd3; a_sign2 = 4'd16; a_sign3 = 4'd9;
b_sign0 = 4'd7; b_sign1 = 4'd13; b_sign2 = 4'd3; b_sign3 = 4'd2;
@(posedge clk_i);
shared_exps0 = 8'd140;
shared_exps1 = 8'd125;
a_mant0 = 8'd222; a_mant1 = 8'd26; a_mant2 = 8'd243; a_mant3 = 8'd228;
b_mant0 = 8'd156; b_mant1 = 8'd122; b_mant2 = 8'd29; b_mant3 = 8'd30;
a_exp0 = 10'd326; a_exp1 = 10'd578; a_exp2 = 10'd641; a_exp3 = 10'd360;
b_exp0 = 10'd176; b_exp1 = 10'd467; b_exp2 = 10'd380; b_exp3 = 10'd54;
a_sign0 = 4'd3; a_sign1 = 4'd12; a_sign2 = 4'd3; a_sign3 = 4'd5;
b_sign0 = 4'd9; b_sign1 = 4'd1; b_sign2 = 4'd13; b_sign3 = 4'd15;
@(posedge clk_i);
a_mant0 = 8'd119; a_mant1 = 8'd144; a_mant2 = 8'd192; a_mant3 = 8'd41;
b_mant0 = 8'd13; b_mant1 = 8'd222; b_mant2 = 8'd203; b_mant3 = 8'd33;
a_exp0 = 10'd913; a_exp1 = 10'd72; a_exp2 = 10'd569; a_exp3 = 10'd731;
b_exp0 = 10'd297; b_exp1 = 10'd467; b_exp2 = 10'd608; b_exp3 = 10'd332;
a_sign0 = 4'd15; a_sign1 = 4'd15; a_sign2 = 4'd8; a_sign3 = 4'd12;
b_sign0 = 4'd9; b_sign1 = 4'd6; b_sign2 = 4'd0; b_sign3 = 4'd0;
@(posedge clk_i);
a_mant0 = 8'd79; a_mant1 = 8'd11; a_mant2 = 8'd41; a_mant3 = 8'd64;
b_mant0 = 8'd122; b_mant1 = 8'd212; b_mant2 = 8'd43; b_mant3 = 8'd43;
a_exp0 = 10'd973; a_exp1 = 10'd447; a_exp2 = 10'd866; a_exp3 = 10'd710;
b_exp0 = 10'd1015; b_exp1 = 10'd520; b_exp2 = 10'd455; b_exp3 = 10'd909;
a_sign0 = 4'd7; a_sign1 = 4'd1; a_sign2 = 4'd15; a_sign3 = 4'd11;
b_sign0 = 4'd5; b_sign1 = 4'd15; b_sign2 = 4'd8; b_sign3 = 4'd14;
@(posedge clk_i);
a_mant0 = 8'd5; a_mant1 = 8'd249; a_mant2 = 8'd192; a_mant3 = 8'd21;
b_mant0 = 8'd244; b_mant1 = 8'd60; b_mant2 = 8'd222; b_mant3 = 8'd227;
a_exp0 = 10'd528; a_exp1 = 10'd78; a_exp2 = 10'd911; a_exp3 = 10'd579;
b_exp0 = 10'd646; b_exp1 = 10'd729; b_exp2 = 10'd935; b_exp3 = 10'd608;
a_sign0 = 4'd16; a_sign1 = 4'd6; a_sign2 = 4'd12; a_sign3 = 4'd3;
b_sign0 = 4'd6; b_sign1 = 4'd1; b_sign2 = 4'd6; b_sign3 = 4'd10;
@(posedge clk_i);
a_mant0 = 8'd36; a_mant1 = 8'd18; a_mant2 = 8'd213; a_mant3 = 8'd250;
b_mant0 = 8'd59; b_mant1 = 8'd11; b_mant2 = 8'd164; b_mant3 = 8'd133;
a_exp0 = 10'd788; a_exp1 = 10'd587; a_exp2 = 10'd809; a_exp3 = 10'd762;
b_exp0 = 10'd316; b_exp1 = 10'd817; b_exp2 = 10'd175; b_exp3 = 10'd460;
a_sign0 = 4'd9; a_sign1 = 4'd1; a_sign2 = 4'd8; a_sign3 = 4'd5;
b_sign0 = 4'd5; b_sign1 = 4'd4; b_sign2 = 4'd0; b_sign3 = 4'd8;
@(posedge clk_i);
a_mant0 = 8'd32; a_mant1 = 8'd124; a_mant2 = 8'd161; a_mant3 = 8'd146;
b_mant0 = 8'd250; b_mant1 = 8'd150; b_mant2 = 8'd68; b_mant3 = 8'd133;
a_exp0 = 10'd731; a_exp1 = 10'd50; a_exp2 = 10'd764; a_exp3 = 10'd465;
b_exp0 = 10'd854; b_exp1 = 10'd536; b_exp2 = 10'd254; b_exp3 = 10'd475;
a_sign0 = 4'd4; a_sign1 = 4'd10; a_sign2 = 4'd5; a_sign3 = 4'd2;
b_sign0 = 4'd4; b_sign1 = 4'd10; b_sign2 = 4'd8; b_sign3 = 4'd13;
@(posedge clk_i);
a_mant0 = 8'd84; a_mant1 = 8'd59; a_mant2 = 8'd222; a_mant3 = 8'd242;
b_mant0 = 8'd4; b_mant1 = 8'd220; b_mant2 = 8'd96; b_mant3 = 8'd60;
a_exp0 = 10'd249; a_exp1 = 10'd990; a_exp2 = 10'd534; a_exp3 = 10'd172;
b_exp0 = 10'd195; b_exp1 = 10'd668; b_exp2 = 10'd840; b_exp3 = 10'd589;
a_sign0 = 4'd10; a_sign1 = 4'd5; a_sign2 = 4'd7; a_sign3 = 4'd8;
b_sign0 = 4'd14; b_sign1 = 4'd14; b_sign2 = 4'd13; b_sign3 = 4'd6;
@(posedge clk_i);
a_mant0 = 8'd165; a_mant1 = 8'd248; a_mant2 = 8'd39; a_mant3 = 8'd235;
b_mant0 = 8'd184; b_mant1 = 8'd65; b_mant2 = 8'd107; b_mant3 = 8'd249;
a_exp0 = 10'd811; a_exp1 = 10'd853; a_exp2 = 10'd768; a_exp3 = 10'd795;
b_exp0 = 10'd110; b_exp1 = 10'd388; b_exp2 = 10'd600; b_exp3 = 10'd60;
a_sign0 = 4'd15; a_sign1 = 4'd0; a_sign2 = 4'd4; a_sign3 = 4'd14;
b_sign0 = 4'd13; b_sign1 = 4'd0; b_sign2 = 4'd5; b_sign3 = 4'd15;
@(posedge clk_i);
shared_exps0 = 8'd145;
shared_exps1 = 8'd108;
rstn = 0;
@(posedge clk_i);
rstn = 1;
a_mant0 = 8'd187; a_mant1 = 8'd104; a_mant2 = 8'd53; a_mant3 = 8'd15;
b_mant0 = 8'd254; b_mant1 = 8'd39; b_mant2 = 8'd211; b_mant3 = 8'd28;
a_exp0 = 10'd105; a_exp1 = 10'd998; a_exp2 = 10'd709; a_exp3 = 10'd870;
b_exp0 = 10'd886; b_exp1 = 10'd784; b_exp2 = 10'd374; b_exp3 = 10'd8;
a_sign0 = 4'd16; a_sign1 = 4'd7; a_sign2 = 4'd9; a_sign3 = 4'd10;
b_sign0 = 4'd13; b_sign1 = 4'd16; b_sign2 = 4'd2; b_sign3 = 4'd7;
@(posedge clk_i);
a_mant0 = 8'd119; a_mant1 = 8'd53; a_mant2 = 8'd236; a_mant3 = 8'd122;
b_mant0 = 8'd255; b_mant1 = 8'd117; b_mant2 = 8'd246; b_mant3 = 8'd99;
a_exp0 = 10'd197; a_exp1 = 10'd833; a_exp2 = 10'd562; a_exp3 = 10'd21;
b_exp0 = 10'd559; b_exp1 = 10'd657; b_exp2 = 10'd697; b_exp3 = 10'd276;
a_sign0 = 4'd5; a_sign1 = 4'd3; a_sign2 = 4'd15; a_sign3 = 4'd15;
b_sign0 = 4'd2; b_sign1 = 4'd16; b_sign2 = 4'd11; b_sign3 = 4'd13;
@(posedge clk_i);
a_mant0 = 8'd23; a_mant1 = 8'd98; a_mant2 = 8'd160; a_mant3 = 8'd245;
b_mant0 = 8'd246; b_mant1 = 8'd19; b_mant2 = 8'd165; b_mant3 = 8'd191;
a_exp0 = 10'd931; a_exp1 = 10'd299; a_exp2 = 10'd747; a_exp3 = 10'd46;
b_exp0 = 10'd489; b_exp1 = 10'd497; b_exp2 = 10'd208; b_exp3 = 10'd552;
a_sign0 = 4'd0; a_sign1 = 4'd15; a_sign2 = 4'd3; a_sign3 = 4'd6;
b_sign0 = 4'd10; b_sign1 = 4'd8; b_sign2 = 4'd5; b_sign3 = 4'd2;
@(posedge clk_i);
a_mant0 = 8'd12; a_mant1 = 8'd173; a_mant2 = 8'd132; a_mant3 = 8'd201;
b_mant0 = 8'd75; b_mant1 = 8'd242; b_mant2 = 8'd56; b_mant3 = 8'd62;
a_exp0 = 10'd968; a_exp1 = 10'd954; a_exp2 = 10'd880; a_exp3 = 10'd749;
b_exp0 = 10'd374; b_exp1 = 10'd819; b_exp2 = 10'd959; b_exp3 = 10'd587;
a_sign0 = 4'd5; a_sign1 = 4'd5; a_sign2 = 4'd5; a_sign3 = 4'd14;
b_sign0 = 4'd4; b_sign1 = 4'd12; b_sign2 = 4'd15; b_sign3 = 4'd5;
@(posedge clk_i);
a_mant0 = 8'd51; a_mant1 = 8'd195; a_mant2 = 8'd113; a_mant3 = 8'd29;
b_mant0 = 8'd251; b_mant1 = 8'd61; b_mant2 = 8'd146; b_mant3 = 8'd10;
a_exp0 = 10'd335; a_exp1 = 10'd637; a_exp2 = 10'd616; a_exp3 = 10'd21;
b_exp0 = 10'd888; b_exp1 = 10'd596; b_exp2 = 10'd664; b_exp3 = 10'd860;
a_sign0 = 4'd10; a_sign1 = 4'd10; a_sign2 = 4'd9; a_sign3 = 4'd11;
b_sign0 = 4'd6; b_sign1 = 4'd16; b_sign2 = 4'd3; b_sign3 = 4'd8;
@(posedge clk_i);
a_mant0 = 8'd22; a_mant1 = 8'd14; a_mant2 = 8'd240; a_mant3 = 8'd162;
b_mant0 = 8'd59; b_mant1 = 8'd165; b_mant2 = 8'd5; b_mant3 = 8'd161;
a_exp0 = 10'd229; a_exp1 = 10'd163; a_exp2 = 10'd835; a_exp3 = 10'd412;
b_exp0 = 10'd607; b_exp1 = 10'd627; b_exp2 = 10'd800; b_exp3 = 10'd122;
a_sign0 = 4'd7; a_sign1 = 4'd13; a_sign2 = 4'd11; a_sign3 = 4'd8;
b_sign0 = 4'd2; b_sign1 = 4'd4; b_sign2 = 4'd16; b_sign3 = 4'd12;
@(posedge clk_i);
a_mant0 = 8'd187; a_mant1 = 8'd168; a_mant2 = 8'd180; a_mant3 = 8'd97;
b_mant0 = 8'd117; b_mant1 = 8'd59; b_mant2 = 8'd37; b_mant3 = 8'd40;
a_exp0 = 10'd129; a_exp1 = 10'd921; a_exp2 = 10'd247; a_exp3 = 10'd876;
b_exp0 = 10'd796; b_exp1 = 10'd373; b_exp2 = 10'd35; b_exp3 = 10'd551;
a_sign0 = 4'd10; a_sign1 = 4'd6; a_sign2 = 4'd2; a_sign3 = 4'd4;
b_sign0 = 4'd4; b_sign1 = 4'd11; b_sign2 = 4'd1; b_sign3 = 4'd16;
@(posedge clk_i);
shared_exps0 = 8'd131;
shared_exps1 = 8'd118;
a_mant0 = 8'd23; a_mant1 = 8'd111; a_mant2 = 8'd181; a_mant3 = 8'd26;
b_mant0 = 8'd198; b_mant1 = 8'd12; b_mant2 = 8'd54; b_mant3 = 8'd163;
a_exp0 = 10'd517; a_exp1 = 10'd52; a_exp2 = 10'd903; a_exp3 = 10'd700;
b_exp0 = 10'd352; b_exp1 = 10'd79; b_exp2 = 10'd680; b_exp3 = 10'd647;
a_sign0 = 4'd9; a_sign1 = 4'd9; a_sign2 = 4'd16; a_sign3 = 4'd2;
b_sign0 = 4'd6; b_sign1 = 4'd1; b_sign2 = 4'd7; b_sign3 = 4'd3;
@(posedge clk_i);
a_mant0 = 8'd115; a_mant1 = 8'd118; a_mant2 = 8'd93; a_mant3 = 8'd8;
b_mant0 = 8'd8; b_mant1 = 8'd104; b_mant2 = 8'd6; b_mant3 = 8'd62;
a_exp0 = 10'd625; a_exp1 = 10'd256; a_exp2 = 10'd940; a_exp3 = 10'd823;
b_exp0 = 10'd795; b_exp1 = 10'd179; b_exp2 = 10'd469; b_exp3 = 10'd731;
a_sign0 = 4'd2; a_sign1 = 4'd11; a_sign2 = 4'd15; a_sign3 = 4'd11;
b_sign0 = 4'd8; b_sign1 = 4'd8; b_sign2 = 4'd10; b_sign3 = 4'd13;
@(posedge clk_i);
a_mant0 = 8'd56; a_mant1 = 8'd200; a_mant2 = 8'd171; a_mant3 = 8'd30;
b_mant0 = 8'd186; b_mant1 = 8'd201; b_mant2 = 8'd216; b_mant3 = 8'd171;
a_exp0 = 10'd190; a_exp1 = 10'd135; a_exp2 = 10'd671; a_exp3 = 10'd996;
b_exp0 = 10'd326; b_exp1 = 10'd705; b_exp2 = 10'd498; b_exp3 = 10'd585;
a_sign0 = 4'd16; a_sign1 = 4'd10; a_sign2 = 4'd11; a_sign3 = 4'd12;
b_sign0 = 4'd16; b_sign1 = 4'd15; b_sign2 = 4'd14; b_sign3 = 4'd14;
@(posedge clk_i);
a_mant0 = 8'd1; a_mant1 = 8'd202; a_mant2 = 8'd88; a_mant3 = 8'd250;
b_mant0 = 8'd137; b_mant1 = 8'd174; b_mant2 = 8'd147; b_mant3 = 8'd65;
a_exp0 = 10'd250; a_exp1 = 10'd172; a_exp2 = 10'd98; a_exp3 = 10'd125;
b_exp0 = 10'd331; b_exp1 = 10'd974; b_exp2 = 10'd66; b_exp3 = 10'd260;
a_sign0 = 4'd15; a_sign1 = 4'd10; a_sign2 = 4'd8; a_sign3 = 4'd2;
b_sign0 = 4'd14; b_sign1 = 4'd13; b_sign2 = 4'd0; b_sign3 = 4'd10;
@(posedge clk_i);
a_mant0 = 8'd3; a_mant1 = 8'd217; a_mant2 = 8'd86; a_mant3 = 8'd217;
b_mant0 = 8'd2; b_mant1 = 8'd171; b_mant2 = 8'd172; b_mant3 = 8'd90;
a_exp0 = 10'd89; a_exp1 = 10'd598; a_exp2 = 10'd594; a_exp3 = 10'd207;
b_exp0 = 10'd901; b_exp1 = 10'd686; b_exp2 = 10'd665; b_exp3 = 10'd757;
a_sign0 = 4'd14; a_sign1 = 4'd7; a_sign2 = 4'd4; a_sign3 = 4'd0;
b_sign0 = 4'd2; b_sign1 = 4'd12; b_sign2 = 4'd15; b_sign3 = 4'd1;
@(posedge clk_i);
a_mant0 = 8'd254; a_mant1 = 8'd212; a_mant2 = 8'd207; a_mant3 = 8'd242;
b_mant0 = 8'd77; b_mant1 = 8'd210; b_mant2 = 8'd145; b_mant3 = 8'd97;
a_exp0 = 10'd182; a_exp1 = 10'd740; a_exp2 = 10'd686; a_exp3 = 10'd200;
b_exp0 = 10'd509; b_exp1 = 10'd175; b_exp2 = 10'd769; b_exp3 = 10'd494;
a_sign0 = 4'd12; a_sign1 = 4'd6; a_sign2 = 4'd10; a_sign3 = 4'd15;
b_sign0 = 4'd15; b_sign1 = 4'd6; b_sign2 = 4'd14; b_sign3 = 4'd13;
@(posedge clk_i);
a_mant0 = 8'd25; a_mant1 = 8'd189; a_mant2 = 8'd213; a_mant3 = 8'd79;
b_mant0 = 8'd234; b_mant1 = 8'd61; b_mant2 = 8'd239; b_mant3 = 8'd172;
a_exp0 = 10'd734; a_exp1 = 10'd352; a_exp2 = 10'd846; a_exp3 = 10'd275;
b_exp0 = 10'd495; b_exp1 = 10'd104; b_exp2 = 10'd808; b_exp3 = 10'd290;
a_sign0 = 4'd15; a_sign1 = 4'd12; a_sign2 = 4'd1; a_sign3 = 4'd16;
b_sign0 = 4'd15; b_sign1 = 4'd1; b_sign2 = 4'd15; b_sign3 = 4'd8;
@(posedge clk_i);
a_mant0 = 8'd61; a_mant1 = 8'd218; a_mant2 = 8'd56; a_mant3 = 8'd179;
b_mant0 = 8'd219; b_mant1 = 8'd142; b_mant2 = 8'd124; b_mant3 = 8'd163;
a_exp0 = 10'd661; a_exp1 = 10'd881; a_exp2 = 10'd942; a_exp3 = 10'd1;
b_exp0 = 10'd572; b_exp1 = 10'd391; b_exp2 = 10'd313; b_exp3 = 10'd448;
a_sign0 = 4'd8; a_sign1 = 4'd8; a_sign2 = 4'd10; a_sign3 = 4'd13;
b_sign0 = 4'd14; b_sign1 = 4'd4; b_sign2 = 4'd8; b_sign3 = 4'd5;
@(posedge clk_i);
shared_exps0 = 8'd147;
shared_exps1 = 8'd138;
a_mant0 = 8'd21; a_mant1 = 8'd96; a_mant2 = 8'd188; a_mant3 = 8'd241;
b_mant0 = 8'd94; b_mant1 = 8'd138; b_mant2 = 8'd33; b_mant3 = 8'd22;
a_exp0 = 10'd645; a_exp1 = 10'd498; a_exp2 = 10'd905; a_exp3 = 10'd909;
b_exp0 = 10'd713; b_exp1 = 10'd669; b_exp2 = 10'd595; b_exp3 = 10'd666;
a_sign0 = 4'd13; a_sign1 = 4'd8; a_sign2 = 4'd0; a_sign3 = 4'd0;
b_sign0 = 4'd4; b_sign1 = 4'd9; b_sign2 = 4'd12; b_sign3 = 4'd4;
@(posedge clk_i);
a_mant0 = 8'd116; a_mant1 = 8'd225; a_mant2 = 8'd0; a_mant3 = 8'd121;
b_mant0 = 8'd23; b_mant1 = 8'd187; b_mant2 = 8'd73; b_mant3 = 8'd91;
a_exp0 = 10'd161; a_exp1 = 10'd889; a_exp2 = 10'd324; a_exp3 = 10'd540;
b_exp0 = 10'd536; b_exp1 = 10'd855; b_exp2 = 10'd179; b_exp3 = 10'd8;
a_sign0 = 4'd5; a_sign1 = 4'd16; a_sign2 = 4'd0; a_sign3 = 4'd13;
b_sign0 = 4'd9; b_sign1 = 4'd5; b_sign2 = 4'd7; b_sign3 = 4'd12;
@(posedge clk_i);
a_mant0 = 8'd15; a_mant1 = 8'd46; a_mant2 = 8'd187; a_mant3 = 8'd220;
b_mant0 = 8'd57; b_mant1 = 8'd105; b_mant2 = 8'd118; b_mant3 = 8'd133;
a_exp0 = 10'd107; a_exp1 = 10'd160; a_exp2 = 10'd167; a_exp3 = 10'd391;
b_exp0 = 10'd234; b_exp1 = 10'd348; b_exp2 = 10'd679; b_exp3 = 10'd475;
a_sign0 = 4'd1; a_sign1 = 4'd7; a_sign2 = 4'd15; a_sign3 = 4'd1;
b_sign0 = 4'd9; b_sign1 = 4'd14; b_sign2 = 4'd12; b_sign3 = 4'd10;
@(posedge clk_i);
a_mant0 = 8'd113; a_mant1 = 8'd33; a_mant2 = 8'd248; a_mant3 = 8'd88;
b_mant0 = 8'd115; b_mant1 = 8'd124; b_mant2 = 8'd108; b_mant3 = 8'd192;
a_exp0 = 10'd610; a_exp1 = 10'd29; a_exp2 = 10'd37; a_exp3 = 10'd780;
b_exp0 = 10'd97; b_exp1 = 10'd668; b_exp2 = 10'd580; b_exp3 = 10'd911;
a_sign0 = 4'd0; a_sign1 = 4'd2; a_sign2 = 4'd8; a_sign3 = 4'd6;
b_sign0 = 4'd3; b_sign1 = 4'd15; b_sign2 = 4'd9; b_sign3 = 4'd5;
@(posedge clk_i);
a_mant0 = 8'd170; a_mant1 = 8'd177; a_mant2 = 8'd26; a_mant3 = 8'd13;
b_mant0 = 8'd232; b_mant1 = 8'd153; b_mant2 = 8'd213; b_mant3 = 8'd100;
a_exp0 = 10'd29; a_exp1 = 10'd116; a_exp2 = 10'd449; a_exp3 = 10'd298;
b_exp0 = 10'd165; b_exp1 = 10'd600; b_exp2 = 10'd435; b_exp3 = 10'd841;
a_sign0 = 4'd8; a_sign1 = 4'd4; a_sign2 = 4'd9; a_sign3 = 4'd11;
b_sign0 = 4'd3; b_sign1 = 4'd6; b_sign2 = 4'd15; b_sign3 = 4'd9;
@(posedge clk_i);
a_mant0 = 8'd190; a_mant1 = 8'd169; a_mant2 = 8'd208; a_mant3 = 8'd116;
b_mant0 = 8'd248; b_mant1 = 8'd17; b_mant2 = 8'd146; b_mant3 = 8'd216;
a_exp0 = 10'd553; a_exp1 = 10'd1012; a_exp2 = 10'd162; a_exp3 = 10'd930;
b_exp0 = 10'd144; b_exp1 = 10'd871; b_exp2 = 10'd260; b_exp3 = 10'd101;
a_sign0 = 4'd14; a_sign1 = 4'd0; a_sign2 = 4'd9; a_sign3 = 4'd14;
b_sign0 = 4'd2; b_sign1 = 4'd15; b_sign2 = 4'd3; b_sign3 = 4'd2;
@(posedge clk_i);
a_mant0 = 8'd83; a_mant1 = 8'd150; a_mant2 = 8'd126; a_mant3 = 8'd199;
b_mant0 = 8'd43; b_mant1 = 8'd233; b_mant2 = 8'd100; b_mant3 = 8'd216;
a_exp0 = 10'd745; a_exp1 = 10'd658; a_exp2 = 10'd321; a_exp3 = 10'd813;
b_exp0 = 10'd666; b_exp1 = 10'd970; b_exp2 = 10'd312; b_exp3 = 10'd1022;
a_sign0 = 4'd3; a_sign1 = 4'd14; a_sign2 = 4'd7; a_sign3 = 4'd11;
b_sign0 = 4'd11; b_sign1 = 4'd4; b_sign2 = 4'd9; b_sign3 = 4'd4;
@(posedge clk_i);
a_mant0 = 8'd52; a_mant1 = 8'd17; a_mant2 = 8'd86; a_mant3 = 8'd221;
b_mant0 = 8'd54; b_mant1 = 8'd204; b_mant2 = 8'd1; b_mant3 = 8'd193;
a_exp0 = 10'd158; a_exp1 = 10'd289; a_exp2 = 10'd9; a_exp3 = 10'd37;
b_exp0 = 10'd803; b_exp1 = 10'd337; b_exp2 = 10'd800; b_exp3 = 10'd108;
a_sign0 = 4'd2; a_sign1 = 4'd9; a_sign2 = 4'd8; a_sign3 = 4'd9;
b_sign0 = 4'd7; b_sign1 = 4'd5; b_sign2 = 4'd14; b_sign3 = 4'd2;
@(posedge clk_i);
shared_exps0 = 8'd103;
shared_exps1 = 8'd113;
a_mant0 = 8'd64; a_mant1 = 8'd101; a_mant2 = 8'd112; a_mant3 = 8'd79;
b_mant0 = 8'd146; b_mant1 = 8'd179; b_mant2 = 8'd208; b_mant3 = 8'd40;
a_exp0 = 10'd992; a_exp1 = 10'd229; a_exp2 = 10'd344; a_exp3 = 10'd970;
b_exp0 = 10'd485; b_exp1 = 10'd52; b_exp2 = 10'd125; b_exp3 = 10'd2;
a_sign0 = 4'd8; a_sign1 = 4'd15; a_sign2 = 4'd7; a_sign3 = 4'd13;
b_sign0 = 4'd2; b_sign1 = 4'd0; b_sign2 = 4'd1; b_sign3 = 4'd12;
@(posedge clk_i);
a_mant0 = 8'd219; a_mant1 = 8'd229; a_mant2 = 8'd185; a_mant3 = 8'd242;
b_mant0 = 8'd135; b_mant1 = 8'd2; b_mant2 = 8'd73; b_mant3 = 8'd29;
a_exp0 = 10'd426; a_exp1 = 10'd988; a_exp2 = 10'd176; a_exp3 = 10'd430;
b_exp0 = 10'd181; b_exp1 = 10'd79; b_exp2 = 10'd669; b_exp3 = 10'd162;
a_sign0 = 4'd12; a_sign1 = 4'd16; a_sign2 = 4'd2; a_sign3 = 4'd6;
b_sign0 = 4'd3; b_sign1 = 4'd12; b_sign2 = 4'd3; b_sign3 = 4'd12;
@(posedge clk_i);
a_mant0 = 8'd114; a_mant1 = 8'd237; a_mant2 = 8'd105; a_mant3 = 8'd142;
b_mant0 = 8'd25; b_mant1 = 8'd93; b_mant2 = 8'd206; b_mant3 = 8'd234;
a_exp0 = 10'd813; a_exp1 = 10'd316; a_exp2 = 10'd391; a_exp3 = 10'd929;
b_exp0 = 10'd129; b_exp1 = 10'd923; b_exp2 = 10'd172; b_exp3 = 10'd460;
a_sign0 = 4'd2; a_sign1 = 4'd8; a_sign2 = 4'd11; a_sign3 = 4'd7;
b_sign0 = 4'd5; b_sign1 = 4'd15; b_sign2 = 4'd4; b_sign3 = 4'd12;
@(posedge clk_i);
a_mant0 = 8'd56; a_mant1 = 8'd137; a_mant2 = 8'd228; a_mant3 = 8'd164;
b_mant0 = 8'd30; b_mant1 = 8'd120; b_mant2 = 8'd211; b_mant3 = 8'd253;
a_exp0 = 10'd230; a_exp1 = 10'd404; a_exp2 = 10'd493; a_exp3 = 10'd911;
b_exp0 = 10'd180; b_exp1 = 10'd745; b_exp2 = 10'd875; b_exp3 = 10'd188;
a_sign0 = 4'd10; a_sign1 = 4'd11; a_sign2 = 4'd13; a_sign3 = 4'd15;
b_sign0 = 4'd2; b_sign1 = 4'd11; b_sign2 = 4'd15; b_sign3 = 4'd5;
@(posedge clk_i);
a_mant0 = 8'd191; a_mant1 = 8'd49; a_mant2 = 8'd210; a_mant3 = 8'd10;
b_mant0 = 8'd72; b_mant1 = 8'd63; b_mant2 = 8'd170; b_mant3 = 8'd171;
a_exp0 = 10'd483; a_exp1 = 10'd707; a_exp2 = 10'd369; a_exp3 = 10'd535;
b_exp0 = 10'd803; b_exp1 = 10'd779; b_exp2 = 10'd470; b_exp3 = 10'd576;
a_sign0 = 4'd1; a_sign1 = 4'd14; a_sign2 = 4'd14; a_sign3 = 4'd16;
b_sign0 = 4'd6; b_sign1 = 4'd5; b_sign2 = 4'd14; b_sign3 = 4'd4;
@(posedge clk_i);
a_mant0 = 8'd171; a_mant1 = 8'd146; a_mant2 = 8'd232; a_mant3 = 8'd214;
b_mant0 = 8'd141; b_mant1 = 8'd146; b_mant2 = 8'd74; b_mant3 = 8'd72;
a_exp0 = 10'd433; a_exp1 = 10'd980; a_exp2 = 10'd159; a_exp3 = 10'd587;
b_exp0 = 10'd201; b_exp1 = 10'd809; b_exp2 = 10'd68; b_exp3 = 10'd91;
a_sign0 = 4'd10; a_sign1 = 4'd5; a_sign2 = 4'd16; a_sign3 = 4'd12;
b_sign0 = 4'd8; b_sign1 = 4'd8; b_sign2 = 4'd10; b_sign3 = 4'd2;
@(posedge clk_i);
a_mant0 = 8'd237; a_mant1 = 8'd231; a_mant2 = 8'd35; a_mant3 = 8'd74;
b_mant0 = 8'd228; b_mant1 = 8'd59; b_mant2 = 8'd247; b_mant3 = 8'd57;
a_exp0 = 10'd276; a_exp1 = 10'd302; a_exp2 = 10'd163; a_exp3 = 10'd969;
b_exp0 = 10'd736; b_exp1 = 10'd950; b_exp2 = 10'd676; b_exp3 = 10'd278;
a_sign0 = 4'd0; a_sign1 = 4'd13; a_sign2 = 4'd16; a_sign3 = 4'd9;
b_sign0 = 4'd7; b_sign1 = 4'd11; b_sign2 = 4'd9; b_sign3 = 4'd12;
@(posedge clk_i);
a_mant0 = 8'd232; a_mant1 = 8'd199; a_mant2 = 8'd236; a_mant3 = 8'd233;
b_mant0 = 8'd69; b_mant1 = 8'd126; b_mant2 = 8'd16; b_mant3 = 8'd113;
a_exp0 = 10'd323; a_exp1 = 10'd220; a_exp2 = 10'd614; a_exp3 = 10'd599;
b_exp0 = 10'd185; b_exp1 = 10'd30; b_exp2 = 10'd96; b_exp3 = 10'd829;
a_sign0 = 4'd1; a_sign1 = 4'd8; a_sign2 = 4'd15; a_sign3 = 4'd11;
b_sign0 = 4'd12; b_sign1 = 4'd13; b_sign2 = 4'd5; b_sign3 = 4'd15;
@(posedge clk_i);
shared_exps0 = 8'd138;
shared_exps1 = 8'd140;
rstn = 0;
@(posedge clk_i);
rstn = 1;
a_mant0 = 8'd245; a_mant1 = 8'd70; a_mant2 = 8'd187; a_mant3 = 8'd188;
b_mant0 = 8'd142; b_mant1 = 8'd179; b_mant2 = 8'd171; b_mant3 = 8'd126;
a_exp0 = 10'd194; a_exp1 = 10'd394; a_exp2 = 10'd276; a_exp3 = 10'd793;
b_exp0 = 10'd570; b_exp1 = 10'd83; b_exp2 = 10'd126; b_exp3 = 10'd335;
a_sign0 = 4'd1; a_sign1 = 4'd2; a_sign2 = 4'd3; a_sign3 = 4'd1;
b_sign0 = 4'd8; b_sign1 = 4'd14; b_sign2 = 4'd7; b_sign3 = 4'd10;
@(posedge clk_i);
a_mant0 = 8'd188; a_mant1 = 8'd184; a_mant2 = 8'd69; a_mant3 = 8'd42;
b_mant0 = 8'd150; b_mant1 = 8'd70; b_mant2 = 8'd149; b_mant3 = 8'd69;
a_exp0 = 10'd3; a_exp1 = 10'd399; a_exp2 = 10'd361; a_exp3 = 10'd21;
b_exp0 = 10'd1020; b_exp1 = 10'd530; b_exp2 = 10'd785; b_exp3 = 10'd895;
a_sign0 = 4'd4; a_sign1 = 4'd6; a_sign2 = 4'd10; a_sign3 = 4'd16;
b_sign0 = 4'd3; b_sign1 = 4'd16; b_sign2 = 4'd9; b_sign3 = 4'd11;
@(posedge clk_i);
a_mant0 = 8'd81; a_mant1 = 8'd123; a_mant2 = 8'd37; a_mant3 = 8'd92;
b_mant0 = 8'd12; b_mant1 = 8'd167; b_mant2 = 8'd148; b_mant3 = 8'd9;
a_exp0 = 10'd874; a_exp1 = 10'd922; a_exp2 = 10'd190; a_exp3 = 10'd203;
b_exp0 = 10'd719; b_exp1 = 10'd495; b_exp2 = 10'd231; b_exp3 = 10'd664;
a_sign0 = 4'd9; a_sign1 = 4'd6; a_sign2 = 4'd3; a_sign3 = 4'd15;
b_sign0 = 4'd15; b_sign1 = 4'd3; b_sign2 = 4'd12; b_sign3 = 4'd12;
@(posedge clk_i);
a_mant0 = 8'd214; a_mant1 = 8'd151; a_mant2 = 8'd39; a_mant3 = 8'd83;
b_mant0 = 8'd214; b_mant1 = 8'd216; b_mant2 = 8'd69; b_mant3 = 8'd173;
a_exp0 = 10'd437; a_exp1 = 10'd737; a_exp2 = 10'd486; a_exp3 = 10'd190;
b_exp0 = 10'd589; b_exp1 = 10'd804; b_exp2 = 10'd522; b_exp3 = 10'd131;
a_sign0 = 4'd16; a_sign1 = 4'd14; a_sign2 = 4'd3; a_sign3 = 4'd11;
b_sign0 = 4'd14; b_sign1 = 4'd3; b_sign2 = 4'd6; b_sign3 = 4'd12;
@(posedge clk_i);
a_mant0 = 8'd242; a_mant1 = 8'd160; a_mant2 = 8'd41; a_mant3 = 8'd26;
b_mant0 = 8'd63; b_mant1 = 8'd87; b_mant2 = 8'd7; b_mant3 = 8'd61;
a_exp0 = 10'd747; a_exp1 = 10'd83; a_exp2 = 10'd830; a_exp3 = 10'd419;
b_exp0 = 10'd389; b_exp1 = 10'd851; b_exp2 = 10'd284; b_exp3 = 10'd573;
a_sign0 = 4'd15; a_sign1 = 4'd10; a_sign2 = 4'd1; a_sign3 = 4'd15;
b_sign0 = 4'd9; b_sign1 = 4'd2; b_sign2 = 4'd0; b_sign3 = 4'd0;
@(posedge clk_i);
a_mant0 = 8'd205; a_mant1 = 8'd44; a_mant2 = 8'd156; a_mant3 = 8'd141;
b_mant0 = 8'd39; b_mant1 = 8'd66; b_mant2 = 8'd28; b_mant3 = 8'd109;
a_exp0 = 10'd214; a_exp1 = 10'd9; a_exp2 = 10'd318; a_exp3 = 10'd50;
b_exp0 = 10'd673; b_exp1 = 10'd708; b_exp2 = 10'd512; b_exp3 = 10'd20;
a_sign0 = 4'd13; a_sign1 = 4'd3; a_sign2 = 4'd9; a_sign3 = 4'd2;
b_sign0 = 4'd3; b_sign1 = 4'd0; b_sign2 = 4'd6; b_sign3 = 4'd13;
@(posedge clk_i);
a_mant0 = 8'd95; a_mant1 = 8'd184; a_mant2 = 8'd189; a_mant3 = 8'd126;
b_mant0 = 8'd155; b_mant1 = 8'd70; b_mant2 = 8'd203; b_mant3 = 8'd148;
a_exp0 = 10'd554; a_exp1 = 10'd995; a_exp2 = 10'd886; a_exp3 = 10'd874;
b_exp0 = 10'd443; b_exp1 = 10'd274; b_exp2 = 10'd37; b_exp3 = 10'd610;
a_sign0 = 4'd0; a_sign1 = 4'd11; a_sign2 = 4'd13; a_sign3 = 4'd7;
b_sign0 = 4'd6; b_sign1 = 4'd9; b_sign2 = 4'd0; b_sign3 = 4'd10;
@(posedge clk_i);
shared_exps0 = 8'd115;
shared_exps1 = 8'd123;
a_mant0 = 8'd242; a_mant1 = 8'd145; a_mant2 = 8'd251; a_mant3 = 8'd115;
b_mant0 = 8'd126; b_mant1 = 8'd17; b_mant2 = 8'd254; b_mant3 = 8'd77;
a_exp0 = 10'd308; a_exp1 = 10'd44; a_exp2 = 10'd383; a_exp3 = 10'd758;
b_exp0 = 10'd758; b_exp1 = 10'd804; b_exp2 = 10'd406; b_exp3 = 10'd33;
a_sign0 = 4'd13; a_sign1 = 4'd16; a_sign2 = 4'd14; a_sign3 = 4'd7;
b_sign0 = 4'd2; b_sign1 = 4'd15; b_sign2 = 4'd13; b_sign3 = 4'd3;
@(posedge clk_i);
a_mant0 = 8'd162; a_mant1 = 8'd238; a_mant2 = 8'd93; a_mant3 = 8'd238;
b_mant0 = 8'd119; b_mant1 = 8'd88; b_mant2 = 8'd44; b_mant3 = 8'd148;
a_exp0 = 10'd434; a_exp1 = 10'd673; a_exp2 = 10'd192; a_exp3 = 10'd560;
b_exp0 = 10'd107; b_exp1 = 10'd997; b_exp2 = 10'd441; b_exp3 = 10'd903;
a_sign0 = 4'd16; a_sign1 = 4'd5; a_sign2 = 4'd0; a_sign3 = 4'd12;
b_sign0 = 4'd11; b_sign1 = 4'd14; b_sign2 = 4'd16; b_sign3 = 4'd1;
@(posedge clk_i);
a_mant0 = 8'd8; a_mant1 = 8'd129; a_mant2 = 8'd223; a_mant3 = 8'd68;
b_mant0 = 8'd74; b_mant1 = 8'd54; b_mant2 = 8'd145; b_mant3 = 8'd68;
a_exp0 = 10'd334; a_exp1 = 10'd496; a_exp2 = 10'd19; a_exp3 = 10'd250;
b_exp0 = 10'd323; b_exp1 = 10'd257; b_exp2 = 10'd290; b_exp3 = 10'd256;
a_sign0 = 4'd6; a_sign1 = 4'd9; a_sign2 = 4'd7; a_sign3 = 4'd12;
b_sign0 = 4'd4; b_sign1 = 4'd7; b_sign2 = 4'd2; b_sign3 = 4'd10;
@(posedge clk_i);
a_mant0 = 8'd152; a_mant1 = 8'd54; a_mant2 = 8'd208; a_mant3 = 8'd249;
b_mant0 = 8'd87; b_mant1 = 8'd207; b_mant2 = 8'd86; b_mant3 = 8'd51;
a_exp0 = 10'd382; a_exp1 = 10'd4; a_exp2 = 10'd984; a_exp3 = 10'd752;
b_exp0 = 10'd507; b_exp1 = 10'd608; b_exp2 = 10'd87; b_exp3 = 10'd787;
a_sign0 = 4'd1; a_sign1 = 4'd6; a_sign2 = 4'd14; a_sign3 = 4'd16;
b_sign0 = 4'd10; b_sign1 = 4'd10; b_sign2 = 4'd9; b_sign3 = 4'd12;
@(posedge clk_i);
a_mant0 = 8'd69; a_mant1 = 8'd130; a_mant2 = 8'd227; a_mant3 = 8'd220;
b_mant0 = 8'd225; b_mant1 = 8'd56; b_mant2 = 8'd157; b_mant3 = 8'd71;
a_exp0 = 10'd44; a_exp1 = 10'd658; a_exp2 = 10'd703; a_exp3 = 10'd115;
b_exp0 = 10'd574; b_exp1 = 10'd800; b_exp2 = 10'd533; b_exp3 = 10'd75;
a_sign0 = 4'd6; a_sign1 = 4'd3; a_sign2 = 4'd7; a_sign3 = 4'd7;
b_sign0 = 4'd9; b_sign1 = 4'd1; b_sign2 = 4'd9; b_sign3 = 4'd2;
@(posedge clk_i);
a_mant0 = 8'd44; a_mant1 = 8'd182; a_mant2 = 8'd222; a_mant3 = 8'd77;
b_mant0 = 8'd50; b_mant1 = 8'd205; b_mant2 = 8'd186; b_mant3 = 8'd38;
a_exp0 = 10'd97; a_exp1 = 10'd196; a_exp2 = 10'd645; a_exp3 = 10'd382;
b_exp0 = 10'd240; b_exp1 = 10'd888; b_exp2 = 10'd759; b_exp3 = 10'd177;
a_sign0 = 4'd10; a_sign1 = 4'd0; a_sign2 = 4'd7; a_sign3 = 4'd13;
b_sign0 = 4'd5; b_sign1 = 4'd2; b_sign2 = 4'd11; b_sign3 = 4'd4;
@(posedge clk_i);
a_mant0 = 8'd35; a_mant1 = 8'd227; a_mant2 = 8'd39; a_mant3 = 8'd2;
b_mant0 = 8'd91; b_mant1 = 8'd78; b_mant2 = 8'd73; b_mant3 = 8'd82;
a_exp0 = 10'd598; a_exp1 = 10'd263; a_exp2 = 10'd732; a_exp3 = 10'd838;
b_exp0 = 10'd753; b_exp1 = 10'd111; b_exp2 = 10'd253; b_exp3 = 10'd694;
a_sign0 = 4'd9; a_sign1 = 4'd13; a_sign2 = 4'd2; a_sign3 = 4'd5;
b_sign0 = 4'd8; b_sign1 = 4'd3; b_sign2 = 4'd14; b_sign3 = 4'd3;
@(posedge clk_i);
a_mant0 = 8'd18; a_mant1 = 8'd122; a_mant2 = 8'd95; a_mant3 = 8'd208;
b_mant0 = 8'd199; b_mant1 = 8'd107; b_mant2 = 8'd255; b_mant3 = 8'd40;
a_exp0 = 10'd180; a_exp1 = 10'd834; a_exp2 = 10'd931; a_exp3 = 10'd758;
b_exp0 = 10'd98; b_exp1 = 10'd651; b_exp2 = 10'd1; b_exp3 = 10'd500;
a_sign0 = 4'd6; a_sign1 = 4'd9; a_sign2 = 4'd0; a_sign3 = 4'd13;
b_sign0 = 4'd2; b_sign1 = 4'd1; b_sign2 = 4'd6; b_sign3 = 4'd4;
@(posedge clk_i);
shared_exps0 = 8'd125;
shared_exps1 = 8'd139;
a_mant0 = 8'd138; a_mant1 = 8'd136; a_mant2 = 8'd89; a_mant3 = 8'd87;
b_mant0 = 8'd141; b_mant1 = 8'd142; b_mant2 = 8'd254; b_mant3 = 8'd111;
a_exp0 = 10'd650; a_exp1 = 10'd890; a_exp2 = 10'd729; a_exp3 = 10'd541;
b_exp0 = 10'd462; b_exp1 = 10'd1002; b_exp2 = 10'd213; b_exp3 = 10'd715;
a_sign0 = 4'd0; a_sign1 = 4'd14; a_sign2 = 4'd15; a_sign3 = 4'd3;
b_sign0 = 4'd2; b_sign1 = 4'd4; b_sign2 = 4'd4; b_sign3 = 4'd13;
@(posedge clk_i);
a_mant0 = 8'd188; a_mant1 = 8'd196; a_mant2 = 8'd104; a_mant3 = 8'd235;
b_mant0 = 8'd47; b_mant1 = 8'd24; b_mant2 = 8'd27; b_mant3 = 8'd172;
a_exp0 = 10'd559; a_exp1 = 10'd592; a_exp2 = 10'd767; a_exp3 = 10'd509;
b_exp0 = 10'd962; b_exp1 = 10'd998; b_exp2 = 10'd466; b_exp3 = 10'd935;
a_sign0 = 4'd1; a_sign1 = 4'd10; a_sign2 = 4'd8; a_sign3 = 4'd2;
b_sign0 = 4'd4; b_sign1 = 4'd2; b_sign2 = 4'd12; b_sign3 = 4'd16;
@(posedge clk_i);
a_mant0 = 8'd154; a_mant1 = 8'd88; a_mant2 = 8'd168; a_mant3 = 8'd188;
b_mant0 = 8'd42; b_mant1 = 8'd158; b_mant2 = 8'd189; b_mant3 = 8'd106;
a_exp0 = 10'd524; a_exp1 = 10'd408; a_exp2 = 10'd658; a_exp3 = 10'd560;
b_exp0 = 10'd771; b_exp1 = 10'd835; b_exp2 = 10'd718; b_exp3 = 10'd139;
a_sign0 = 4'd0; a_sign1 = 4'd5; a_sign2 = 4'd0; a_sign3 = 4'd9;
b_sign0 = 4'd9; b_sign1 = 4'd11; b_sign2 = 4'd2; b_sign3 = 4'd0;
@(posedge clk_i);
a_mant0 = 8'd183; a_mant1 = 8'd103; a_mant2 = 8'd7; a_mant3 = 8'd199;
b_mant0 = 8'd218; b_mant1 = 8'd159; b_mant2 = 8'd125; b_mant3 = 8'd59;
a_exp0 = 10'd34; a_exp1 = 10'd156; a_exp2 = 10'd122; a_exp3 = 10'd835;
b_exp0 = 10'd116; b_exp1 = 10'd481; b_exp2 = 10'd396; b_exp3 = 10'd801;
a_sign0 = 4'd4; a_sign1 = 4'd16; a_sign2 = 4'd1; a_sign3 = 4'd15;
b_sign0 = 4'd13; b_sign1 = 4'd5; b_sign2 = 4'd15; b_sign3 = 4'd4;
@(posedge clk_i);
a_mant0 = 8'd184; a_mant1 = 8'd155; a_mant2 = 8'd27; a_mant3 = 8'd82;
b_mant0 = 8'd29; b_mant1 = 8'd124; b_mant2 = 8'd230; b_mant3 = 8'd161;
a_exp0 = 10'd695; a_exp1 = 10'd566; a_exp2 = 10'd9; a_exp3 = 10'd539;
b_exp0 = 10'd129; b_exp1 = 10'd108; b_exp2 = 10'd852; b_exp3 = 10'd123;
a_sign0 = 4'd10; a_sign1 = 4'd7; a_sign2 = 4'd1; a_sign3 = 4'd3;
b_sign0 = 4'd14; b_sign1 = 4'd6; b_sign2 = 4'd14; b_sign3 = 4'd8;
@(posedge clk_i);
a_mant0 = 8'd8; a_mant1 = 8'd199; a_mant2 = 8'd39; a_mant3 = 8'd32;
b_mant0 = 8'd115; b_mant1 = 8'd176; b_mant2 = 8'd218; b_mant3 = 8'd15;
a_exp0 = 10'd784; a_exp1 = 10'd259; a_exp2 = 10'd928; a_exp3 = 10'd516;
b_exp0 = 10'd219; b_exp1 = 10'd803; b_exp2 = 10'd734; b_exp3 = 10'd794;
a_sign0 = 4'd8; a_sign1 = 4'd7; a_sign2 = 4'd11; a_sign3 = 4'd1;
b_sign0 = 4'd9; b_sign1 = 4'd6; b_sign2 = 4'd15; b_sign3 = 4'd14;
@(posedge clk_i);
a_mant0 = 8'd96; a_mant1 = 8'd60; a_mant2 = 8'd120; a_mant3 = 8'd10;
b_mant0 = 8'd202; b_mant1 = 8'd124; b_mant2 = 8'd98; b_mant3 = 8'd169;
a_exp0 = 10'd851; a_exp1 = 10'd958; a_exp2 = 10'd672; a_exp3 = 10'd128;
b_exp0 = 10'd1006; b_exp1 = 10'd115; b_exp2 = 10'd165; b_exp3 = 10'd685;
a_sign0 = 4'd16; a_sign1 = 4'd12; a_sign2 = 4'd6; a_sign3 = 4'd7;
b_sign0 = 4'd11; b_sign1 = 4'd0; b_sign2 = 4'd7; b_sign3 = 4'd9;
@(posedge clk_i);
a_mant0 = 8'd228; a_mant1 = 8'd96; a_mant2 = 8'd141; a_mant3 = 8'd158;
b_mant0 = 8'd103; b_mant1 = 8'd209; b_mant2 = 8'd97; b_mant3 = 8'd138;
a_exp0 = 10'd957; a_exp1 = 10'd481; a_exp2 = 10'd653; a_exp3 = 10'd507;
b_exp0 = 10'd268; b_exp1 = 10'd964; b_exp2 = 10'd690; b_exp3 = 10'd929;
a_sign0 = 4'd15; a_sign1 = 4'd10; a_sign2 = 4'd11; a_sign3 = 4'd13;
b_sign0 = 4'd11; b_sign1 = 4'd11; b_sign2 = 4'd8; b_sign3 = 4'd2;
@(posedge clk_i);
shared_exps0 = 8'd117;
shared_exps1 = 8'd134;
a_mant0 = 8'd215; a_mant1 = 8'd234; a_mant2 = 8'd248; a_mant3 = 8'd135;
b_mant0 = 8'd163; b_mant1 = 8'd167; b_mant2 = 8'd228; b_mant3 = 8'd200;
a_exp0 = 10'd476; a_exp1 = 10'd582; a_exp2 = 10'd33; a_exp3 = 10'd531;
b_exp0 = 10'd938; b_exp1 = 10'd407; b_exp2 = 10'd408; b_exp3 = 10'd176;
a_sign0 = 4'd13; a_sign1 = 4'd7; a_sign2 = 4'd2; a_sign3 = 4'd1;
b_sign0 = 4'd8; b_sign1 = 4'd1; b_sign2 = 4'd9; b_sign3 = 4'd6;
@(posedge clk_i);
a_mant0 = 8'd8; a_mant1 = 8'd220; a_mant2 = 8'd155; a_mant3 = 8'd166;
b_mant0 = 8'd39; b_mant1 = 8'd115; b_mant2 = 8'd153; b_mant3 = 8'd110;
a_exp0 = 10'd982; a_exp1 = 10'd766; a_exp2 = 10'd381; a_exp3 = 10'd609;
b_exp0 = 10'd115; b_exp1 = 10'd108; b_exp2 = 10'd467; b_exp3 = 10'd500;
a_sign0 = 4'd16; a_sign1 = 4'd11; a_sign2 = 4'd13; a_sign3 = 4'd14;
b_sign0 = 4'd14; b_sign1 = 4'd15; b_sign2 = 4'd12; b_sign3 = 4'd9;
@(posedge clk_i);
a_mant0 = 8'd254; a_mant1 = 8'd53; a_mant2 = 8'd59; a_mant3 = 8'd140;
b_mant0 = 8'd252; b_mant1 = 8'd223; b_mant2 = 8'd69; b_mant3 = 8'd157;
a_exp0 = 10'd857; a_exp1 = 10'd673; a_exp2 = 10'd975; a_exp3 = 10'd869;
b_exp0 = 10'd156; b_exp1 = 10'd1021; b_exp2 = 10'd819; b_exp3 = 10'd198;
a_sign0 = 4'd3; a_sign1 = 4'd1; a_sign2 = 4'd2; a_sign3 = 4'd11;
b_sign0 = 4'd14; b_sign1 = 4'd16; b_sign2 = 4'd10; b_sign3 = 4'd14;
@(posedge clk_i);
a_mant0 = 8'd147; a_mant1 = 8'd169; a_mant2 = 8'd200; a_mant3 = 8'd173;
b_mant0 = 8'd62; b_mant1 = 8'd21; b_mant2 = 8'd140; b_mant3 = 8'd244;
a_exp0 = 10'd142; a_exp1 = 10'd255; a_exp2 = 10'd726; a_exp3 = 10'd858;
b_exp0 = 10'd907; b_exp1 = 10'd762; b_exp2 = 10'd96; b_exp3 = 10'd575;
a_sign0 = 4'd7; a_sign1 = 4'd9; a_sign2 = 4'd6; a_sign3 = 4'd9;
b_sign0 = 4'd10; b_sign1 = 4'd0; b_sign2 = 4'd13; b_sign3 = 4'd4;
@(posedge clk_i);
a_mant0 = 8'd187; a_mant1 = 8'd252; a_mant2 = 8'd85; a_mant3 = 8'd103;
b_mant0 = 8'd85; b_mant1 = 8'd232; b_mant2 = 8'd1; b_mant3 = 8'd163;
a_exp0 = 10'd508; a_exp1 = 10'd485; a_exp2 = 10'd71; a_exp3 = 10'd621;
b_exp0 = 10'd469; b_exp1 = 10'd668; b_exp2 = 10'd634; b_exp3 = 10'd888;
a_sign0 = 4'd6; a_sign1 = 4'd1; a_sign2 = 4'd13; a_sign3 = 4'd2;
b_sign0 = 4'd2; b_sign1 = 4'd0; b_sign2 = 4'd0; b_sign3 = 4'd0;
@(posedge clk_i);
a_mant0 = 8'd78; a_mant1 = 8'd12; a_mant2 = 8'd186; a_mant3 = 8'd209;
b_mant0 = 8'd163; b_mant1 = 8'd169; b_mant2 = 8'd222; b_mant3 = 8'd20;
a_exp0 = 10'd943; a_exp1 = 10'd221; a_exp2 = 10'd424; a_exp3 = 10'd650;
b_exp0 = 10'd631; b_exp1 = 10'd230; b_exp2 = 10'd965; b_exp3 = 10'd408;
a_sign0 = 4'd13; a_sign1 = 4'd7; a_sign2 = 4'd0; a_sign3 = 4'd5;
b_sign0 = 4'd10; b_sign1 = 4'd16; b_sign2 = 4'd15; b_sign3 = 4'd6;
@(posedge clk_i);
a_mant0 = 8'd158; a_mant1 = 8'd124; a_mant2 = 8'd194; a_mant3 = 8'd207;
b_mant0 = 8'd67; b_mant1 = 8'd4; b_mant2 = 8'd50; b_mant3 = 8'd149;
a_exp0 = 10'd858; a_exp1 = 10'd166; a_exp2 = 10'd130; a_exp3 = 10'd295;
b_exp0 = 10'd938; b_exp1 = 10'd729; b_exp2 = 10'd606; b_exp3 = 10'd337;
a_sign0 = 4'd13; a_sign1 = 4'd3; a_sign2 = 4'd10; a_sign3 = 4'd11;
b_sign0 = 4'd15; b_sign1 = 4'd14; b_sign2 = 4'd7; b_sign3 = 4'd16;
@(posedge clk_i);
a_mant0 = 8'd158; a_mant1 = 8'd80; a_mant2 = 8'd208; a_mant3 = 8'd92;
b_mant0 = 8'd2; b_mant1 = 8'd229; b_mant2 = 8'd243; b_mant3 = 8'd235;
a_exp0 = 10'd634; a_exp1 = 10'd120; a_exp2 = 10'd389; a_exp3 = 10'd54;
b_exp0 = 10'd548; b_exp1 = 10'd150; b_exp2 = 10'd351; b_exp3 = 10'd654;
a_sign0 = 4'd7; a_sign1 = 4'd14; a_sign2 = 4'd11; a_sign3 = 4'd5;
b_sign0 = 4'd8; b_sign1 = 4'd15; b_sign2 = 4'd14; b_sign3 = 4'd3;
@(posedge clk_i);
shared_exps0 = 8'd137;
shared_exps1 = 8'd111;
rstn = 0;
@(posedge clk_i);
rstn = 1;
a_mant0 = 8'd51; a_mant1 = 8'd216; a_mant2 = 8'd142; a_mant3 = 8'd38;
b_mant0 = 8'd223; b_mant1 = 8'd220; b_mant2 = 8'd216; b_mant3 = 8'd146;
a_exp0 = 10'd806; a_exp1 = 10'd135; a_exp2 = 10'd902; a_exp3 = 10'd554;
b_exp0 = 10'd640; b_exp1 = 10'd263; b_exp2 = 10'd834; b_exp3 = 10'd332;
a_sign0 = 4'd7; a_sign1 = 4'd14; a_sign2 = 4'd6; a_sign3 = 4'd16;
b_sign0 = 4'd13; b_sign1 = 4'd4; b_sign2 = 4'd4; b_sign3 = 4'd13;
@(posedge clk_i);
a_mant0 = 8'd225; a_mant1 = 8'd107; a_mant2 = 8'd208; a_mant3 = 8'd202;
b_mant0 = 8'd218; b_mant1 = 8'd54; b_mant2 = 8'd156; b_mant3 = 8'd115;
a_exp0 = 10'd347; a_exp1 = 10'd339; a_exp2 = 10'd483; a_exp3 = 10'd715;
b_exp0 = 10'd230; b_exp1 = 10'd504; b_exp2 = 10'd237; b_exp3 = 10'd442;
a_sign0 = 4'd10; a_sign1 = 4'd2; a_sign2 = 4'd2; a_sign3 = 4'd16;
b_sign0 = 4'd10; b_sign1 = 4'd6; b_sign2 = 4'd4; b_sign3 = 4'd6;
@(posedge clk_i);
a_mant0 = 8'd58; a_mant1 = 8'd15; a_mant2 = 8'd179; a_mant3 = 8'd88;
b_mant0 = 8'd196; b_mant1 = 8'd20; b_mant2 = 8'd222; b_mant3 = 8'd247;
a_exp0 = 10'd987; a_exp1 = 10'd167; a_exp2 = 10'd224; a_exp3 = 10'd492;
b_exp0 = 10'd306; b_exp1 = 10'd104; b_exp2 = 10'd829; b_exp3 = 10'd64;
a_sign0 = 4'd6; a_sign1 = 4'd15; a_sign2 = 4'd0; a_sign3 = 4'd7;
b_sign0 = 4'd6; b_sign1 = 4'd0; b_sign2 = 4'd13; b_sign3 = 4'd2;
@(posedge clk_i);
a_mant0 = 8'd196; a_mant1 = 8'd27; a_mant2 = 8'd27; a_mant3 = 8'd91;
b_mant0 = 8'd216; b_mant1 = 8'd207; b_mant2 = 8'd127; b_mant3 = 8'd187;
a_exp0 = 10'd961; a_exp1 = 10'd140; a_exp2 = 10'd410; a_exp3 = 10'd552;
b_exp0 = 10'd515; b_exp1 = 10'd349; b_exp2 = 10'd267; b_exp3 = 10'd990;
a_sign0 = 4'd0; a_sign1 = 4'd0; a_sign2 = 4'd7; a_sign3 = 4'd7;
b_sign0 = 4'd6; b_sign1 = 4'd2; b_sign2 = 4'd0; b_sign3 = 4'd13;
@(posedge clk_i);
a_mant0 = 8'd84; a_mant1 = 8'd33; a_mant2 = 8'd93; a_mant3 = 8'd166;
b_mant0 = 8'd134; b_mant1 = 8'd248; b_mant2 = 8'd63; b_mant3 = 8'd29;
a_exp0 = 10'd802; a_exp1 = 10'd911; a_exp2 = 10'd607; a_exp3 = 10'd522;
b_exp0 = 10'd433; b_exp1 = 10'd916; b_exp2 = 10'd739; b_exp3 = 10'd198;
a_sign0 = 4'd16; a_sign1 = 4'd7; a_sign2 = 4'd14; a_sign3 = 4'd3;
b_sign0 = 4'd7; b_sign1 = 4'd13; b_sign2 = 4'd3; b_sign3 = 4'd3;
@(posedge clk_i);
a_mant0 = 8'd224; a_mant1 = 8'd59; a_mant2 = 8'd19; a_mant3 = 8'd82;
b_mant0 = 8'd230; b_mant1 = 8'd207; b_mant2 = 8'd253; b_mant3 = 8'd88;
a_exp0 = 10'd984; a_exp1 = 10'd638; a_exp2 = 10'd488; a_exp3 = 10'd72;
b_exp0 = 10'd457; b_exp1 = 10'd689; b_exp2 = 10'd31; b_exp3 = 10'd434;
a_sign0 = 4'd9; a_sign1 = 4'd12; a_sign2 = 4'd13; a_sign3 = 4'd14;
b_sign0 = 4'd15; b_sign1 = 4'd8; b_sign2 = 4'd7; b_sign3 = 4'd1;
@(posedge clk_i);
a_mant0 = 8'd43; a_mant1 = 8'd101; a_mant2 = 8'd192; a_mant3 = 8'd191;
b_mant0 = 8'd253; b_mant1 = 8'd102; b_mant2 = 8'd186; b_mant3 = 8'd143;
a_exp0 = 10'd1023; a_exp1 = 10'd925; a_exp2 = 10'd1002; a_exp3 = 10'd291;
b_exp0 = 10'd608; b_exp1 = 10'd572; b_exp2 = 10'd757; b_exp3 = 10'd594;
a_sign0 = 4'd4; a_sign1 = 4'd12; a_sign2 = 4'd12; a_sign3 = 4'd4;
b_sign0 = 4'd16; b_sign1 = 4'd2; b_sign2 = 4'd11; b_sign3 = 4'd1;
@(posedge clk_i);
shared_exps0 = 8'd108;
shared_exps1 = 8'd129;
a_mant0 = 8'd140; a_mant1 = 8'd184; a_mant2 = 8'd3; a_mant3 = 8'd204;
b_mant0 = 8'd171; b_mant1 = 8'd171; b_mant2 = 8'd182; b_mant3 = 8'd91;
a_exp0 = 10'd705; a_exp1 = 10'd493; a_exp2 = 10'd76; a_exp3 = 10'd721;
b_exp0 = 10'd59; b_exp1 = 10'd452; b_exp2 = 10'd746; b_exp3 = 10'd452;
a_sign0 = 4'd9; a_sign1 = 4'd7; a_sign2 = 4'd10; a_sign3 = 4'd8;
b_sign0 = 4'd1; b_sign1 = 4'd12; b_sign2 = 4'd3; b_sign3 = 4'd12;
@(posedge clk_i);
a_mant0 = 8'd57; a_mant1 = 8'd126; a_mant2 = 8'd138; a_mant3 = 8'd233;
b_mant0 = 8'd234; b_mant1 = 8'd233; b_mant2 = 8'd151; b_mant3 = 8'd166;
a_exp0 = 10'd524; a_exp1 = 10'd112; a_exp2 = 10'd551; a_exp3 = 10'd938;
b_exp0 = 10'd59; b_exp1 = 10'd177; b_exp2 = 10'd335; b_exp3 = 10'd339;
a_sign0 = 4'd0; a_sign1 = 4'd15; a_sign2 = 4'd12; a_sign3 = 4'd14;
b_sign0 = 4'd15; b_sign1 = 4'd7; b_sign2 = 4'd15; b_sign3 = 4'd12;
@(posedge clk_i);
a_mant0 = 8'd1; a_mant1 = 8'd33; a_mant2 = 8'd153; a_mant3 = 8'd75;
b_mant0 = 8'd8; b_mant1 = 8'd95; b_mant2 = 8'd247; b_mant3 = 8'd75;
a_exp0 = 10'd823; a_exp1 = 10'd183; a_exp2 = 10'd835; a_exp3 = 10'd490;
b_exp0 = 10'd661; b_exp1 = 10'd239; b_exp2 = 10'd845; b_exp3 = 10'd343;
a_sign0 = 4'd9; a_sign1 = 4'd14; a_sign2 = 4'd9; a_sign3 = 4'd10;
b_sign0 = 4'd6; b_sign1 = 4'd2; b_sign2 = 4'd10; b_sign3 = 4'd16;
@(posedge clk_i);
a_mant0 = 8'd227; a_mant1 = 8'd117; a_mant2 = 8'd27; a_mant3 = 8'd77;
b_mant0 = 8'd114; b_mant1 = 8'd30; b_mant2 = 8'd65; b_mant3 = 8'd129;
a_exp0 = 10'd42; a_exp1 = 10'd628; a_exp2 = 10'd931; a_exp3 = 10'd1005;
b_exp0 = 10'd712; b_exp1 = 10'd295; b_exp2 = 10'd335; b_exp3 = 10'd580;
a_sign0 = 4'd8; a_sign1 = 4'd10; a_sign2 = 4'd3; a_sign3 = 4'd12;
b_sign0 = 4'd3; b_sign1 = 4'd15; b_sign2 = 4'd8; b_sign3 = 4'd8;
@(posedge clk_i);
a_mant0 = 8'd83; a_mant1 = 8'd170; a_mant2 = 8'd156; a_mant3 = 8'd92;
b_mant0 = 8'd27; b_mant1 = 8'd160; b_mant2 = 8'd214; b_mant3 = 8'd173;
a_exp0 = 10'd335; a_exp1 = 10'd200; a_exp2 = 10'd808; a_exp3 = 10'd361;
b_exp0 = 10'd553; b_exp1 = 10'd1005; b_exp2 = 10'd481; b_exp3 = 10'd302;
a_sign0 = 4'd1; a_sign1 = 4'd6; a_sign2 = 4'd2; a_sign3 = 4'd7;
b_sign0 = 4'd11; b_sign1 = 4'd14; b_sign2 = 4'd10; b_sign3 = 4'd10;
@(posedge clk_i);
a_mant0 = 8'd250; a_mant1 = 8'd152; a_mant2 = 8'd164; a_mant3 = 8'd61;
b_mant0 = 8'd121; b_mant1 = 8'd90; b_mant2 = 8'd213; b_mant3 = 8'd139;
a_exp0 = 10'd738; a_exp1 = 10'd641; a_exp2 = 10'd180; a_exp3 = 10'd897;
b_exp0 = 10'd698; b_exp1 = 10'd388; b_exp2 = 10'd878; b_exp3 = 10'd950;
a_sign0 = 4'd10; a_sign1 = 4'd3; a_sign2 = 4'd0; a_sign3 = 4'd10;
b_sign0 = 4'd6; b_sign1 = 4'd12; b_sign2 = 4'd12; b_sign3 = 4'd3;
@(posedge clk_i);
a_mant0 = 8'd97; a_mant1 = 8'd79; a_mant2 = 8'd117; a_mant3 = 8'd250;
b_mant0 = 8'd99; b_mant1 = 8'd26; b_mant2 = 8'd233; b_mant3 = 8'd14;
a_exp0 = 10'd498; a_exp1 = 10'd417; a_exp2 = 10'd774; a_exp3 = 10'd270;
b_exp0 = 10'd11; b_exp1 = 10'd566; b_exp2 = 10'd70; b_exp3 = 10'd586;
a_sign0 = 4'd9; a_sign1 = 4'd0; a_sign2 = 4'd6; a_sign3 = 4'd2;
b_sign0 = 4'd12; b_sign1 = 4'd3; b_sign2 = 4'd3; b_sign3 = 4'd4;
@(posedge clk_i);
a_mant0 = 8'd209; a_mant1 = 8'd56; a_mant2 = 8'd47; a_mant3 = 8'd83;
b_mant0 = 8'd188; b_mant1 = 8'd156; b_mant2 = 8'd94; b_mant3 = 8'd241;
a_exp0 = 10'd638; a_exp1 = 10'd865; a_exp2 = 10'd680; a_exp3 = 10'd273;
b_exp0 = 10'd735; b_exp1 = 10'd309; b_exp2 = 10'd122; b_exp3 = 10'd131;
a_sign0 = 4'd2; a_sign1 = 4'd0; a_sign2 = 4'd9; a_sign3 = 4'd15;
b_sign0 = 4'd13; b_sign1 = 4'd9; b_sign2 = 4'd8; b_sign3 = 4'd13;
@(posedge clk_i);
shared_exps0 = 8'd118;
shared_exps1 = 8'd132;
a_mant0 = 8'd24; a_mant1 = 8'd171; a_mant2 = 8'd64; a_mant3 = 8'd63;
b_mant0 = 8'd105; b_mant1 = 8'd244; b_mant2 = 8'd243; b_mant3 = 8'd142;
a_exp0 = 10'd613; a_exp1 = 10'd707; a_exp2 = 10'd877; a_exp3 = 10'd96;
b_exp0 = 10'd910; b_exp1 = 10'd390; b_exp2 = 10'd922; b_exp3 = 10'd657;
a_sign0 = 4'd10; a_sign1 = 4'd9; a_sign2 = 4'd14; a_sign3 = 4'd0;
b_sign0 = 4'd14; b_sign1 = 4'd1; b_sign2 = 4'd8; b_sign3 = 4'd7;
@(posedge clk_i);
a_mant0 = 8'd58; a_mant1 = 8'd109; a_mant2 = 8'd187; a_mant3 = 8'd213;
b_mant0 = 8'd68; b_mant1 = 8'd71; b_mant2 = 8'd255; b_mant3 = 8'd237;
a_exp0 = 10'd317; a_exp1 = 10'd789; a_exp2 = 10'd318; a_exp3 = 10'd978;
b_exp0 = 10'd721; b_exp1 = 10'd880; b_exp2 = 10'd351; b_exp3 = 10'd378;
a_sign0 = 4'd4; a_sign1 = 4'd12; a_sign2 = 4'd1; a_sign3 = 4'd0;
b_sign0 = 4'd13; b_sign1 = 4'd0; b_sign2 = 4'd16; b_sign3 = 4'd13;
@(posedge clk_i);
a_mant0 = 8'd34; a_mant1 = 8'd152; a_mant2 = 8'd122; a_mant3 = 8'd11;
b_mant0 = 8'd110; b_mant1 = 8'd195; b_mant2 = 8'd111; b_mant3 = 8'd232;
a_exp0 = 10'd963; a_exp1 = 10'd941; a_exp2 = 10'd781; a_exp3 = 10'd673;
b_exp0 = 10'd693; b_exp1 = 10'd198; b_exp2 = 10'd838; b_exp3 = 10'd202;
a_sign0 = 4'd13; a_sign1 = 4'd2; a_sign2 = 4'd10; a_sign3 = 4'd13;
b_sign0 = 4'd10; b_sign1 = 4'd12; b_sign2 = 4'd5; b_sign3 = 4'd3;
@(posedge clk_i);
a_mant0 = 8'd135; a_mant1 = 8'd120; a_mant2 = 8'd177; a_mant3 = 8'd224;
b_mant0 = 8'd230; b_mant1 = 8'd195; b_mant2 = 8'd242; b_mant3 = 8'd158;
a_exp0 = 10'd707; a_exp1 = 10'd178; a_exp2 = 10'd776; a_exp3 = 10'd891;
b_exp0 = 10'd273; b_exp1 = 10'd470; b_exp2 = 10'd685; b_exp3 = 10'd240;
a_sign0 = 4'd11; a_sign1 = 4'd9; a_sign2 = 4'd11; a_sign3 = 4'd5;
b_sign0 = 4'd11; b_sign1 = 4'd6; b_sign2 = 4'd3; b_sign3 = 4'd15;
@(posedge clk_i);
a_mant0 = 8'd156; a_mant1 = 8'd7; a_mant2 = 8'd237; a_mant3 = 8'd141;
b_mant0 = 8'd54; b_mant1 = 8'd73; b_mant2 = 8'd168; b_mant3 = 8'd49;
a_exp0 = 10'd569; a_exp1 = 10'd854; a_exp2 = 10'd179; a_exp3 = 10'd1008;
b_exp0 = 10'd100; b_exp1 = 10'd182; b_exp2 = 10'd858; b_exp3 = 10'd605;
a_sign0 = 4'd8; a_sign1 = 4'd2; a_sign2 = 4'd9; a_sign3 = 4'd1;
b_sign0 = 4'd6; b_sign1 = 4'd9; b_sign2 = 4'd13; b_sign3 = 4'd10;
@(posedge clk_i);
a_mant0 = 8'd96; a_mant1 = 8'd60; a_mant2 = 8'd225; a_mant3 = 8'd108;
b_mant0 = 8'd114; b_mant1 = 8'd155; b_mant2 = 8'd29; b_mant3 = 8'd153;
a_exp0 = 10'd539; a_exp1 = 10'd780; a_exp2 = 10'd205; a_exp3 = 10'd79;
b_exp0 = 10'd684; b_exp1 = 10'd86; b_exp2 = 10'd117; b_exp3 = 10'd829;
a_sign0 = 4'd10; a_sign1 = 4'd16; a_sign2 = 4'd6; a_sign3 = 4'd15;
b_sign0 = 4'd7; b_sign1 = 4'd9; b_sign2 = 4'd11; b_sign3 = 4'd14;
@(posedge clk_i);
a_mant0 = 8'd208; a_mant1 = 8'd95; a_mant2 = 8'd117; a_mant3 = 8'd236;
b_mant0 = 8'd195; b_mant1 = 8'd49; b_mant2 = 8'd117; b_mant3 = 8'd8;
a_exp0 = 10'd178; a_exp1 = 10'd513; a_exp2 = 10'd161; a_exp3 = 10'd933;
b_exp0 = 10'd479; b_exp1 = 10'd142; b_exp2 = 10'd982; b_exp3 = 10'd905;
a_sign0 = 4'd8; a_sign1 = 4'd16; a_sign2 = 4'd1; a_sign3 = 4'd12;
b_sign0 = 4'd15; b_sign1 = 4'd8; b_sign2 = 4'd3; b_sign3 = 4'd9;
@(posedge clk_i);
a_mant0 = 8'd133; a_mant1 = 8'd3; a_mant2 = 8'd22; a_mant3 = 8'd199;
b_mant0 = 8'd185; b_mant1 = 8'd39; b_mant2 = 8'd67; b_mant3 = 8'd70;
a_exp0 = 10'd1007; a_exp1 = 10'd641; a_exp2 = 10'd326; a_exp3 = 10'd307;
b_exp0 = 10'd5; b_exp1 = 10'd574; b_exp2 = 10'd926; b_exp3 = 10'd783;
a_sign0 = 4'd4; a_sign1 = 4'd3; a_sign2 = 4'd9; a_sign3 = 4'd4;
b_sign0 = 4'd2; b_sign1 = 4'd15; b_sign2 = 4'd0; b_sign3 = 4'd8;
@(posedge clk_i);
shared_exps0 = 8'd132;
shared_exps1 = 8'd118;
a_mant0 = 8'd33; a_mant1 = 8'd57; a_mant2 = 8'd176; a_mant3 = 8'd228;
b_mant0 = 8'd200; b_mant1 = 8'd19; b_mant2 = 8'd82; b_mant3 = 8'd246;
a_exp0 = 10'd107; a_exp1 = 10'd605; a_exp2 = 10'd689; a_exp3 = 10'd627;
b_exp0 = 10'd962; b_exp1 = 10'd179; b_exp2 = 10'd735; b_exp3 = 10'd1022;
a_sign0 = 4'd4; a_sign1 = 4'd6; a_sign2 = 4'd1; a_sign3 = 4'd4;
b_sign0 = 4'd12; b_sign1 = 4'd10; b_sign2 = 4'd3; b_sign3 = 4'd8;
@(posedge clk_i);
a_mant0 = 8'd191; a_mant1 = 8'd226; a_mant2 = 8'd189; a_mant3 = 8'd98;
b_mant0 = 8'd140; b_mant1 = 8'd210; b_mant2 = 8'd204; b_mant3 = 8'd42;
a_exp0 = 10'd116; a_exp1 = 10'd649; a_exp2 = 10'd226; a_exp3 = 10'd673;
b_exp0 = 10'd839; b_exp1 = 10'd492; b_exp2 = 10'd255; b_exp3 = 10'd779;
a_sign0 = 4'd10; a_sign1 = 4'd13; a_sign2 = 4'd10; a_sign3 = 4'd9;
b_sign0 = 4'd10; b_sign1 = 4'd14; b_sign2 = 4'd13; b_sign3 = 4'd0;
@(posedge clk_i);
a_mant0 = 8'd150; a_mant1 = 8'd11; a_mant2 = 8'd28; a_mant3 = 8'd162;
b_mant0 = 8'd74; b_mant1 = 8'd134; b_mant2 = 8'd57; b_mant3 = 8'd81;
a_exp0 = 10'd303; a_exp1 = 10'd672; a_exp2 = 10'd762; a_exp3 = 10'd624;
b_exp0 = 10'd495; b_exp1 = 10'd669; b_exp2 = 10'd451; b_exp3 = 10'd932;
a_sign0 = 4'd5; a_sign1 = 4'd7; a_sign2 = 4'd4; a_sign3 = 4'd14;
b_sign0 = 4'd3; b_sign1 = 4'd5; b_sign2 = 4'd9; b_sign3 = 4'd8;
@(posedge clk_i);
a_mant0 = 8'd234; a_mant1 = 8'd31; a_mant2 = 8'd106; a_mant3 = 8'd189;
b_mant0 = 8'd237; b_mant1 = 8'd159; b_mant2 = 8'd49; b_mant3 = 8'd81;
a_exp0 = 10'd442; a_exp1 = 10'd828; a_exp2 = 10'd673; a_exp3 = 10'd657;
b_exp0 = 10'd357; b_exp1 = 10'd49; b_exp2 = 10'd581; b_exp3 = 10'd944;
a_sign0 = 4'd7; a_sign1 = 4'd3; a_sign2 = 4'd15; a_sign3 = 4'd16;
b_sign0 = 4'd15; b_sign1 = 4'd0; b_sign2 = 4'd12; b_sign3 = 4'd9;
@(posedge clk_i);
a_mant0 = 8'd5; a_mant1 = 8'd72; a_mant2 = 8'd34; a_mant3 = 8'd24;
b_mant0 = 8'd224; b_mant1 = 8'd98; b_mant2 = 8'd248; b_mant3 = 8'd209;
a_exp0 = 10'd335; a_exp1 = 10'd557; a_exp2 = 10'd329; a_exp3 = 10'd656;
b_exp0 = 10'd606; b_exp1 = 10'd204; b_exp2 = 10'd1009; b_exp3 = 10'd424;
a_sign0 = 4'd2; a_sign1 = 4'd2; a_sign2 = 4'd2; a_sign3 = 4'd16;
b_sign0 = 4'd2; b_sign1 = 4'd0; b_sign2 = 4'd5; b_sign3 = 4'd14;
@(posedge clk_i);
a_mant0 = 8'd168; a_mant1 = 8'd214; a_mant2 = 8'd57; a_mant3 = 8'd113;
b_mant0 = 8'd200; b_mant1 = 8'd80; b_mant2 = 8'd252; b_mant3 = 8'd67;
a_exp0 = 10'd52; a_exp1 = 10'd553; a_exp2 = 10'd234; a_exp3 = 10'd196;
b_exp0 = 10'd303; b_exp1 = 10'd765; b_exp2 = 10'd165; b_exp3 = 10'd92;
a_sign0 = 4'd6; a_sign1 = 4'd3; a_sign2 = 4'd15; a_sign3 = 4'd1;
b_sign0 = 4'd4; b_sign1 = 4'd1; b_sign2 = 4'd11; b_sign3 = 4'd1;
@(posedge clk_i);
a_mant0 = 8'd183; a_mant1 = 8'd153; a_mant2 = 8'd168; a_mant3 = 8'd183;
b_mant0 = 8'd108; b_mant1 = 8'd78; b_mant2 = 8'd39; b_mant3 = 8'd17;
a_exp0 = 10'd502; a_exp1 = 10'd468; a_exp2 = 10'd609; a_exp3 = 10'd324;
b_exp0 = 10'd525; b_exp1 = 10'd182; b_exp2 = 10'd48; b_exp3 = 10'd64;
a_sign0 = 4'd2; a_sign1 = 4'd2; a_sign2 = 4'd9; a_sign3 = 4'd6;
b_sign0 = 4'd12; b_sign1 = 4'd8; b_sign2 = 4'd0; b_sign3 = 4'd2;
@(posedge clk_i);
a_mant0 = 8'd148; a_mant1 = 8'd146; a_mant2 = 8'd71; a_mant3 = 8'd195;
b_mant0 = 8'd236; b_mant1 = 8'd67; b_mant2 = 8'd188; b_mant3 = 8'd55;
a_exp0 = 10'd954; a_exp1 = 10'd514; a_exp2 = 10'd630; a_exp3 = 10'd473;
b_exp0 = 10'd113; b_exp1 = 10'd208; b_exp2 = 10'd431; b_exp3 = 10'd255;
a_sign0 = 4'd0; a_sign1 = 4'd12; a_sign2 = 4'd5; a_sign3 = 4'd5;
b_sign0 = 4'd1; b_sign1 = 4'd13; b_sign2 = 4'd0; b_sign3 = 4'd11;
@(posedge clk_i);
shared_exps0 = 8'd104;
shared_exps1 = 8'd139;
rstn = 0;
@(posedge clk_i);
rstn = 1;
a_mant0 = 8'd85; a_mant1 = 8'd13; a_mant2 = 8'd119; a_mant3 = 8'd149;
b_mant0 = 8'd188; b_mant1 = 8'd128; b_mant2 = 8'd93; b_mant3 = 8'd238;
a_exp0 = 10'd322; a_exp1 = 10'd952; a_exp2 = 10'd196; a_exp3 = 10'd298;
b_exp0 = 10'd213; b_exp1 = 10'd193; b_exp2 = 10'd728; b_exp3 = 10'd685;
a_sign0 = 4'd1; a_sign1 = 4'd1; a_sign2 = 4'd7; a_sign3 = 4'd5;
b_sign0 = 4'd16; b_sign1 = 4'd12; b_sign2 = 4'd13; b_sign3 = 4'd13;
@(posedge clk_i);
a_mant0 = 8'd173; a_mant1 = 8'd191; a_mant2 = 8'd151; a_mant3 = 8'd17;
b_mant0 = 8'd113; b_mant1 = 8'd162; b_mant2 = 8'd205; b_mant3 = 8'd85;
a_exp0 = 10'd775; a_exp1 = 10'd81; a_exp2 = 10'd374; a_exp3 = 10'd512;
b_exp0 = 10'd954; b_exp1 = 10'd513; b_exp2 = 10'd807; b_exp3 = 10'd0;
a_sign0 = 4'd2; a_sign1 = 4'd5; a_sign2 = 4'd0; a_sign3 = 4'd12;
b_sign0 = 4'd8; b_sign1 = 4'd2; b_sign2 = 4'd12; b_sign3 = 4'd13;
@(posedge clk_i);
a_mant0 = 8'd216; a_mant1 = 8'd45; a_mant2 = 8'd158; a_mant3 = 8'd222;
b_mant0 = 8'd59; b_mant1 = 8'd141; b_mant2 = 8'd108; b_mant3 = 8'd208;
a_exp0 = 10'd751; a_exp1 = 10'd4; a_exp2 = 10'd589; a_exp3 = 10'd969;
b_exp0 = 10'd811; b_exp1 = 10'd987; b_exp2 = 10'd598; b_exp3 = 10'd823;
a_sign0 = 4'd13; a_sign1 = 4'd8; a_sign2 = 4'd6; a_sign3 = 4'd8;
b_sign0 = 4'd14; b_sign1 = 4'd1; b_sign2 = 4'd7; b_sign3 = 4'd13;
@(posedge clk_i);
a_mant0 = 8'd56; a_mant1 = 8'd107; a_mant2 = 8'd168; a_mant3 = 8'd159;
b_mant0 = 8'd168; b_mant1 = 8'd70; b_mant2 = 8'd126; b_mant3 = 8'd56;
a_exp0 = 10'd751; a_exp1 = 10'd744; a_exp2 = 10'd973; a_exp3 = 10'd796;
b_exp0 = 10'd604; b_exp1 = 10'd497; b_exp2 = 10'd963; b_exp3 = 10'd13;
a_sign0 = 4'd14; a_sign1 = 4'd12; a_sign2 = 4'd6; a_sign3 = 4'd4;
b_sign0 = 4'd16; b_sign1 = 4'd0; b_sign2 = 4'd0; b_sign3 = 4'd7;
@(posedge clk_i);
a_mant0 = 8'd121; a_mant1 = 8'd94; a_mant2 = 8'd174; a_mant3 = 8'd187;
b_mant0 = 8'd190; b_mant1 = 8'd55; b_mant2 = 8'd231; b_mant3 = 8'd213;
a_exp0 = 10'd782; a_exp1 = 10'd117; a_exp2 = 10'd845; a_exp3 = 10'd200;
b_exp0 = 10'd899; b_exp1 = 10'd737; b_exp2 = 10'd179; b_exp3 = 10'd190;
a_sign0 = 4'd10; a_sign1 = 4'd14; a_sign2 = 4'd16; a_sign3 = 4'd12;
b_sign0 = 4'd16; b_sign1 = 4'd2; b_sign2 = 4'd14; b_sign3 = 4'd0;
@(posedge clk_i);
a_mant0 = 8'd190; a_mant1 = 8'd33; a_mant2 = 8'd153; a_mant3 = 8'd89;
b_mant0 = 8'd194; b_mant1 = 8'd58; b_mant2 = 8'd123; b_mant3 = 8'd235;
a_exp0 = 10'd768; a_exp1 = 10'd611; a_exp2 = 10'd146; a_exp3 = 10'd883;
b_exp0 = 10'd646; b_exp1 = 10'd941; b_exp2 = 10'd891; b_exp3 = 10'd512;
a_sign0 = 4'd0; a_sign1 = 4'd8; a_sign2 = 4'd1; a_sign3 = 4'd15;
b_sign0 = 4'd12; b_sign1 = 4'd0; b_sign2 = 4'd8; b_sign3 = 4'd1;
@(posedge clk_i);
a_mant0 = 8'd209; a_mant1 = 8'd162; a_mant2 = 8'd239; a_mant3 = 8'd31;
b_mant0 = 8'd245; b_mant1 = 8'd231; b_mant2 = 8'd24; b_mant3 = 8'd142;
a_exp0 = 10'd491; a_exp1 = 10'd912; a_exp2 = 10'd391; a_exp3 = 10'd816;
b_exp0 = 10'd211; b_exp1 = 10'd80; b_exp2 = 10'd550; b_exp3 = 10'd729;
a_sign0 = 4'd4; a_sign1 = 4'd6; a_sign2 = 4'd3; a_sign3 = 4'd10;
b_sign0 = 4'd3; b_sign1 = 4'd4; b_sign2 = 4'd10; b_sign3 = 4'd16;
@(posedge clk_i);
shared_exps0 = 8'd151;
shared_exps1 = 8'd109;
a_mant0 = 8'd79; a_mant1 = 8'd182; a_mant2 = 8'd143; a_mant3 = 8'd137;
b_mant0 = 8'd95; b_mant1 = 8'd197; b_mant2 = 8'd135; b_mant3 = 8'd152;
a_exp0 = 10'd1016; a_exp1 = 10'd941; a_exp2 = 10'd419; a_exp3 = 10'd502;
b_exp0 = 10'd712; b_exp1 = 10'd362; b_exp2 = 10'd822; b_exp3 = 10'd520;
a_sign0 = 4'd0; a_sign1 = 4'd3; a_sign2 = 4'd14; a_sign3 = 4'd2;
b_sign0 = 4'd3; b_sign1 = 4'd8; b_sign2 = 4'd5; b_sign3 = 4'd9;
@(posedge clk_i);
a_mant0 = 8'd100; a_mant1 = 8'd145; a_mant2 = 8'd74; a_mant3 = 8'd83;
b_mant0 = 8'd4; b_mant1 = 8'd78; b_mant2 = 8'd26; b_mant3 = 8'd152;
a_exp0 = 10'd494; a_exp1 = 10'd847; a_exp2 = 10'd237; a_exp3 = 10'd729;
b_exp0 = 10'd517; b_exp1 = 10'd483; b_exp2 = 10'd795; b_exp3 = 10'd688;
a_sign0 = 4'd0; a_sign1 = 4'd0; a_sign2 = 4'd16; a_sign3 = 4'd0;
b_sign0 = 4'd12; b_sign1 = 4'd10; b_sign2 = 4'd12; b_sign3 = 4'd1;
@(posedge clk_i);
a_mant0 = 8'd147; a_mant1 = 8'd212; a_mant2 = 8'd159; a_mant3 = 8'd9;
b_mant0 = 8'd59; b_mant1 = 8'd89; b_mant2 = 8'd74; b_mant3 = 8'd40;
a_exp0 = 10'd423; a_exp1 = 10'd597; a_exp2 = 10'd832; a_exp3 = 10'd188;
b_exp0 = 10'd2; b_exp1 = 10'd967; b_exp2 = 10'd4; b_exp3 = 10'd295;
a_sign0 = 4'd14; a_sign1 = 4'd15; a_sign2 = 4'd3; a_sign3 = 4'd8;
b_sign0 = 4'd5; b_sign1 = 4'd9; b_sign2 = 4'd6; b_sign3 = 4'd3;
@(posedge clk_i);
a_mant0 = 8'd236; a_mant1 = 8'd77; a_mant2 = 8'd64; a_mant3 = 8'd147;
b_mant0 = 8'd165; b_mant1 = 8'd124; b_mant2 = 8'd190; b_mant3 = 8'd18;
a_exp0 = 10'd356; a_exp1 = 10'd840; a_exp2 = 10'd825; a_exp3 = 10'd402;
b_exp0 = 10'd321; b_exp1 = 10'd627; b_exp2 = 10'd713; b_exp3 = 10'd913;
a_sign0 = 4'd2; a_sign1 = 4'd14; a_sign2 = 4'd6; a_sign3 = 4'd11;
b_sign0 = 4'd8; b_sign1 = 4'd16; b_sign2 = 4'd12; b_sign3 = 4'd4;
@(posedge clk_i);
a_mant0 = 8'd88; a_mant1 = 8'd80; a_mant2 = 8'd136; a_mant3 = 8'd153;
b_mant0 = 8'd63; b_mant1 = 8'd29; b_mant2 = 8'd252; b_mant3 = 8'd220;
a_exp0 = 10'd448; a_exp1 = 10'd405; a_exp2 = 10'd365; a_exp3 = 10'd969;
b_exp0 = 10'd953; b_exp1 = 10'd802; b_exp2 = 10'd6; b_exp3 = 10'd955;
a_sign0 = 4'd1; a_sign1 = 4'd0; a_sign2 = 4'd14; a_sign3 = 4'd13;
b_sign0 = 4'd3; b_sign1 = 4'd6; b_sign2 = 4'd11; b_sign3 = 4'd14;
@(posedge clk_i);
a_mant0 = 8'd121; a_mant1 = 8'd74; a_mant2 = 8'd49; a_mant3 = 8'd151;
b_mant0 = 8'd215; b_mant1 = 8'd106; b_mant2 = 8'd1; b_mant3 = 8'd228;
a_exp0 = 10'd1021; a_exp1 = 10'd667; a_exp2 = 10'd294; a_exp3 = 10'd899;
b_exp0 = 10'd839; b_exp1 = 10'd545; b_exp2 = 10'd867; b_exp3 = 10'd7;
a_sign0 = 4'd13; a_sign1 = 4'd9; a_sign2 = 4'd4; a_sign3 = 4'd5;
b_sign0 = 4'd9; b_sign1 = 4'd6; b_sign2 = 4'd4; b_sign3 = 4'd9;
@(posedge clk_i);
a_mant0 = 8'd95; a_mant1 = 8'd97; a_mant2 = 8'd89; a_mant3 = 8'd0;
b_mant0 = 8'd29; b_mant1 = 8'd153; b_mant2 = 8'd143; b_mant3 = 8'd137;
a_exp0 = 10'd574; a_exp1 = 10'd783; a_exp2 = 10'd765; a_exp3 = 10'd20;
b_exp0 = 10'd29; b_exp1 = 10'd247; b_exp2 = 10'd921; b_exp3 = 10'd324;
a_sign0 = 4'd13; a_sign1 = 4'd14; a_sign2 = 4'd16; a_sign3 = 4'd16;
b_sign0 = 4'd12; b_sign1 = 4'd3; b_sign2 = 4'd15; b_sign3 = 4'd13;
@(posedge clk_i);
a_mant0 = 8'd243; a_mant1 = 8'd86; a_mant2 = 8'd103; a_mant3 = 8'd72;
b_mant0 = 8'd250; b_mant1 = 8'd71; b_mant2 = 8'd244; b_mant3 = 8'd29;
a_exp0 = 10'd734; a_exp1 = 10'd710; a_exp2 = 10'd402; a_exp3 = 10'd516;
b_exp0 = 10'd550; b_exp1 = 10'd878; b_exp2 = 10'd575; b_exp3 = 10'd802;
a_sign0 = 4'd13; a_sign1 = 4'd14; a_sign2 = 4'd15; a_sign3 = 4'd2;
b_sign0 = 4'd13; b_sign1 = 4'd13; b_sign2 = 4'd0; b_sign3 = 4'd13;
@(posedge clk_i);
shared_exps0 = 8'd118;
shared_exps1 = 8'd153;
a_mant0 = 8'd164; a_mant1 = 8'd71; a_mant2 = 8'd134; a_mant3 = 8'd201;
b_mant0 = 8'd133; b_mant1 = 8'd103; b_mant2 = 8'd200; b_mant3 = 8'd11;
a_exp0 = 10'd780; a_exp1 = 10'd945; a_exp2 = 10'd438; a_exp3 = 10'd942;
b_exp0 = 10'd950; b_exp1 = 10'd859; b_exp2 = 10'd361; b_exp3 = 10'd59;
a_sign0 = 4'd0; a_sign1 = 4'd13; a_sign2 = 4'd13; a_sign3 = 4'd4;
b_sign0 = 4'd2; b_sign1 = 4'd2; b_sign2 = 4'd0; b_sign3 = 4'd15;
@(posedge clk_i);
a_mant0 = 8'd94; a_mant1 = 8'd216; a_mant2 = 8'd172; a_mant3 = 8'd35;
b_mant0 = 8'd1; b_mant1 = 8'd159; b_mant2 = 8'd62; b_mant3 = 8'd233;
a_exp0 = 10'd771; a_exp1 = 10'd126; a_exp2 = 10'd722; a_exp3 = 10'd1017;
b_exp0 = 10'd336; b_exp1 = 10'd847; b_exp2 = 10'd439; b_exp3 = 10'd960;
a_sign0 = 4'd14; a_sign1 = 4'd13; a_sign2 = 4'd7; a_sign3 = 4'd6;
b_sign0 = 4'd14; b_sign1 = 4'd9; b_sign2 = 4'd9; b_sign3 = 4'd7;
@(posedge clk_i);
a_mant0 = 8'd8; a_mant1 = 8'd96; a_mant2 = 8'd249; a_mant3 = 8'd220;
b_mant0 = 8'd239; b_mant1 = 8'd3; b_mant2 = 8'd102; b_mant3 = 8'd159;
a_exp0 = 10'd386; a_exp1 = 10'd677; a_exp2 = 10'd385; a_exp3 = 10'd207;
b_exp0 = 10'd107; b_exp1 = 10'd258; b_exp2 = 10'd546; b_exp3 = 10'd981;
a_sign0 = 4'd5; a_sign1 = 4'd14; a_sign2 = 4'd0; a_sign3 = 4'd15;
b_sign0 = 4'd8; b_sign1 = 4'd13; b_sign2 = 4'd10; b_sign3 = 4'd15;
@(posedge clk_i);
a_mant0 = 8'd49; a_mant1 = 8'd128; a_mant2 = 8'd97; a_mant3 = 8'd136;
b_mant0 = 8'd45; b_mant1 = 8'd242; b_mant2 = 8'd135; b_mant3 = 8'd137;
a_exp0 = 10'd354; a_exp1 = 10'd271; a_exp2 = 10'd616; a_exp3 = 10'd1013;
b_exp0 = 10'd85; b_exp1 = 10'd254; b_exp2 = 10'd569; b_exp3 = 10'd229;
a_sign0 = 4'd14; a_sign1 = 4'd9; a_sign2 = 4'd10; a_sign3 = 4'd15;
b_sign0 = 4'd2; b_sign1 = 4'd10; b_sign2 = 4'd13; b_sign3 = 4'd6;
@(posedge clk_i);
a_mant0 = 8'd107; a_mant1 = 8'd141; a_mant2 = 8'd209; a_mant3 = 8'd70;
b_mant0 = 8'd159; b_mant1 = 8'd72; b_mant2 = 8'd79; b_mant3 = 8'd0;
a_exp0 = 10'd587; a_exp1 = 10'd226; a_exp2 = 10'd646; a_exp3 = 10'd497;
b_exp0 = 10'd937; b_exp1 = 10'd602; b_exp2 = 10'd684; b_exp3 = 10'd504;
a_sign0 = 4'd6; a_sign1 = 4'd16; a_sign2 = 4'd15; a_sign3 = 4'd12;
b_sign0 = 4'd12; b_sign1 = 4'd15; b_sign2 = 4'd1; b_sign3 = 4'd16;
@(posedge clk_i);
a_mant0 = 8'd6; a_mant1 = 8'd85; a_mant2 = 8'd219; a_mant3 = 8'd204;
b_mant0 = 8'd55; b_mant1 = 8'd178; b_mant2 = 8'd22; b_mant3 = 8'd206;
a_exp0 = 10'd34; a_exp1 = 10'd109; a_exp2 = 10'd892; a_exp3 = 10'd128;
b_exp0 = 10'd635; b_exp1 = 10'd786; b_exp2 = 10'd297; b_exp3 = 10'd51;
a_sign0 = 4'd4; a_sign1 = 4'd7; a_sign2 = 4'd5; a_sign3 = 4'd1;
b_sign0 = 4'd11; b_sign1 = 4'd13; b_sign2 = 4'd13; b_sign3 = 4'd4;
@(posedge clk_i);
a_mant0 = 8'd66; a_mant1 = 8'd122; a_mant2 = 8'd93; a_mant3 = 8'd39;
b_mant0 = 8'd209; b_mant1 = 8'd14; b_mant2 = 8'd39; b_mant3 = 8'd198;
a_exp0 = 10'd751; a_exp1 = 10'd702; a_exp2 = 10'd801; a_exp3 = 10'd28;
b_exp0 = 10'd161; b_exp1 = 10'd26; b_exp2 = 10'd387; b_exp3 = 10'd918;
a_sign0 = 4'd4; a_sign1 = 4'd14; a_sign2 = 4'd0; a_sign3 = 4'd5;
b_sign0 = 4'd6; b_sign1 = 4'd2; b_sign2 = 4'd7; b_sign3 = 4'd7;
@(posedge clk_i);
a_mant0 = 8'd237; a_mant1 = 8'd178; a_mant2 = 8'd45; a_mant3 = 8'd12;
b_mant0 = 8'd132; b_mant1 = 8'd241; b_mant2 = 8'd85; b_mant3 = 8'd140;
a_exp0 = 10'd502; a_exp1 = 10'd474; a_exp2 = 10'd552; a_exp3 = 10'd671;
b_exp0 = 10'd487; b_exp1 = 10'd750; b_exp2 = 10'd867; b_exp3 = 10'd191;
a_sign0 = 4'd6; a_sign1 = 4'd13; a_sign2 = 4'd8; a_sign3 = 4'd2;
b_sign0 = 4'd0; b_sign1 = 4'd15; b_sign2 = 4'd6; b_sign3 = 4'd4;
@(posedge clk_i);
shared_exps0 = 8'd131;
shared_exps1 = 8'd122;
a_mant0 = 8'd216; a_mant1 = 8'd29; a_mant2 = 8'd13; a_mant3 = 8'd133;
b_mant0 = 8'd35; b_mant1 = 8'd57; b_mant2 = 8'd100; b_mant3 = 8'd19;
a_exp0 = 10'd459; a_exp1 = 10'd545; a_exp2 = 10'd584; a_exp3 = 10'd796;
b_exp0 = 10'd936; b_exp1 = 10'd699; b_exp2 = 10'd353; b_exp3 = 10'd232;
a_sign0 = 4'd0; a_sign1 = 4'd4; a_sign2 = 4'd13; a_sign3 = 4'd8;
b_sign0 = 4'd10; b_sign1 = 4'd8; b_sign2 = 4'd7; b_sign3 = 4'd8;
@(posedge clk_i);
a_mant0 = 8'd71; a_mant1 = 8'd191; a_mant2 = 8'd116; a_mant3 = 8'd123;
b_mant0 = 8'd37; b_mant1 = 8'd102; b_mant2 = 8'd219; b_mant3 = 8'd232;
a_exp0 = 10'd719; a_exp1 = 10'd459; a_exp2 = 10'd381; a_exp3 = 10'd906;
b_exp0 = 10'd824; b_exp1 = 10'd690; b_exp2 = 10'd868; b_exp3 = 10'd389;
a_sign0 = 4'd11; a_sign1 = 4'd1; a_sign2 = 4'd2; a_sign3 = 4'd12;
b_sign0 = 4'd3; b_sign1 = 4'd7; b_sign2 = 4'd11; b_sign3 = 4'd12;
@(posedge clk_i);
a_mant0 = 8'd119; a_mant1 = 8'd73; a_mant2 = 8'd43; a_mant3 = 8'd15;
b_mant0 = 8'd11; b_mant1 = 8'd102; b_mant2 = 8'd56; b_mant3 = 8'd85;
a_exp0 = 10'd312; a_exp1 = 10'd997; a_exp2 = 10'd368; a_exp3 = 10'd786;
b_exp0 = 10'd486; b_exp1 = 10'd83; b_exp2 = 10'd717; b_exp3 = 10'd148;
a_sign0 = 4'd16; a_sign1 = 4'd8; a_sign2 = 4'd9; a_sign3 = 4'd16;
b_sign0 = 4'd3; b_sign1 = 4'd0; b_sign2 = 4'd8; b_sign3 = 4'd12;
@(posedge clk_i);
a_mant0 = 8'd36; a_mant1 = 8'd9; a_mant2 = 8'd122; a_mant3 = 8'd22;
b_mant0 = 8'd18; b_mant1 = 8'd117; b_mant2 = 8'd60; b_mant3 = 8'd40;
a_exp0 = 10'd625; a_exp1 = 10'd715; a_exp2 = 10'd304; a_exp3 = 10'd81;
b_exp0 = 10'd809; b_exp1 = 10'd82; b_exp2 = 10'd774; b_exp3 = 10'd636;
a_sign0 = 4'd12; a_sign1 = 4'd2; a_sign2 = 4'd5; a_sign3 = 4'd16;
b_sign0 = 4'd10; b_sign1 = 4'd12; b_sign2 = 4'd16; b_sign3 = 4'd5;
@(posedge clk_i);
a_mant0 = 8'd118; a_mant1 = 8'd11; a_mant2 = 8'd50; a_mant3 = 8'd61;
b_mant0 = 8'd30; b_mant1 = 8'd157; b_mant2 = 8'd168; b_mant3 = 8'd70;
a_exp0 = 10'd57; a_exp1 = 10'd264; a_exp2 = 10'd947; a_exp3 = 10'd14;
b_exp0 = 10'd91; b_exp1 = 10'd987; b_exp2 = 10'd2; b_exp3 = 10'd291;
a_sign0 = 4'd2; a_sign1 = 4'd8; a_sign2 = 4'd14; a_sign3 = 4'd2;
b_sign0 = 4'd6; b_sign1 = 4'd3; b_sign2 = 4'd15; b_sign3 = 4'd10;
@(posedge clk_i);
a_mant0 = 8'd101; a_mant1 = 8'd158; a_mant2 = 8'd178; a_mant3 = 8'd68;
b_mant0 = 8'd240; b_mant1 = 8'd196; b_mant2 = 8'd112; b_mant3 = 8'd33;
a_exp0 = 10'd907; a_exp1 = 10'd769; a_exp2 = 10'd719; a_exp3 = 10'd848;
b_exp0 = 10'd280; b_exp1 = 10'd706; b_exp2 = 10'd863; b_exp3 = 10'd436;
a_sign0 = 4'd13; a_sign1 = 4'd6; a_sign2 = 4'd14; a_sign3 = 4'd7;
b_sign0 = 4'd9; b_sign1 = 4'd16; b_sign2 = 4'd9; b_sign3 = 4'd7;
@(posedge clk_i);
a_mant0 = 8'd218; a_mant1 = 8'd100; a_mant2 = 8'd48; a_mant3 = 8'd182;
b_mant0 = 8'd160; b_mant1 = 8'd212; b_mant2 = 8'd108; b_mant3 = 8'd64;
a_exp0 = 10'd590; a_exp1 = 10'd63; a_exp2 = 10'd150; a_exp3 = 10'd710;
b_exp0 = 10'd296; b_exp1 = 10'd1001; b_exp2 = 10'd151; b_exp3 = 10'd491;
a_sign0 = 4'd12; a_sign1 = 4'd4; a_sign2 = 4'd12; a_sign3 = 4'd8;
b_sign0 = 4'd5; b_sign1 = 4'd2; b_sign2 = 4'd7; b_sign3 = 4'd0;
@(posedge clk_i);
a_mant0 = 8'd185; a_mant1 = 8'd31; a_mant2 = 8'd55; a_mant3 = 8'd99;
b_mant0 = 8'd105; b_mant1 = 8'd82; b_mant2 = 8'd69; b_mant3 = 8'd95;
a_exp0 = 10'd768; a_exp1 = 10'd559; a_exp2 = 10'd731; a_exp3 = 10'd806;
b_exp0 = 10'd136; b_exp1 = 10'd869; b_exp2 = 10'd757; b_exp3 = 10'd362;
a_sign0 = 4'd0; a_sign1 = 4'd8; a_sign2 = 4'd1; a_sign3 = 4'd6;
b_sign0 = 4'd6; b_sign1 = 4'd13; b_sign2 = 4'd8; b_sign3 = 4'd5;
@(posedge clk_i);
shared_exps0 = 8'd122;
shared_exps1 = 8'd120;
rstn = 0;
@(posedge clk_i);
rstn = 1;
a_mant0 = 8'd190; a_mant1 = 8'd58; a_mant2 = 8'd98; a_mant3 = 8'd148;
b_mant0 = 8'd106; b_mant1 = 8'd217; b_mant2 = 8'd154; b_mant3 = 8'd247;
a_exp0 = 10'd593; a_exp1 = 10'd246; a_exp2 = 10'd672; a_exp3 = 10'd921;
b_exp0 = 10'd268; b_exp1 = 10'd191; b_exp2 = 10'd716; b_exp3 = 10'd146;
a_sign0 = 4'd0; a_sign1 = 4'd8; a_sign2 = 4'd14; a_sign3 = 4'd9;
b_sign0 = 4'd4; b_sign1 = 4'd4; b_sign2 = 4'd2; b_sign3 = 4'd2;
@(posedge clk_i);
a_mant0 = 8'd222; a_mant1 = 8'd163; a_mant2 = 8'd209; a_mant3 = 8'd7;
b_mant0 = 8'd228; b_mant1 = 8'd34; b_mant2 = 8'd226; b_mant3 = 8'd67;
a_exp0 = 10'd980; a_exp1 = 10'd296; a_exp2 = 10'd987; a_exp3 = 10'd597;
b_exp0 = 10'd989; b_exp1 = 10'd681; b_exp2 = 10'd555; b_exp3 = 10'd13;
a_sign0 = 4'd11; a_sign1 = 4'd13; a_sign2 = 4'd4; a_sign3 = 4'd14;
b_sign0 = 4'd13; b_sign1 = 4'd4; b_sign2 = 4'd14; b_sign3 = 4'd14;
@(posedge clk_i);
a_mant0 = 8'd231; a_mant1 = 8'd15; a_mant2 = 8'd44; a_mant3 = 8'd4;
b_mant0 = 8'd172; b_mant1 = 8'd54; b_mant2 = 8'd60; b_mant3 = 8'd39;
a_exp0 = 10'd770; a_exp1 = 10'd981; a_exp2 = 10'd966; a_exp3 = 10'd198;
b_exp0 = 10'd353; b_exp1 = 10'd315; b_exp2 = 10'd169; b_exp3 = 10'd378;
a_sign0 = 4'd12; a_sign1 = 4'd9; a_sign2 = 4'd6; a_sign3 = 4'd11;
b_sign0 = 4'd1; b_sign1 = 4'd11; b_sign2 = 4'd2; b_sign3 = 4'd4;
@(posedge clk_i);
a_mant0 = 8'd63; a_mant1 = 8'd253; a_mant2 = 8'd226; a_mant3 = 8'd244;
b_mant0 = 8'd119; b_mant1 = 8'd160; b_mant2 = 8'd78; b_mant3 = 8'd247;
a_exp0 = 10'd936; a_exp1 = 10'd1011; a_exp2 = 10'd1003; a_exp3 = 10'd915;
b_exp0 = 10'd410; b_exp1 = 10'd479; b_exp2 = 10'd336; b_exp3 = 10'd781;
a_sign0 = 4'd14; a_sign1 = 4'd8; a_sign2 = 4'd14; a_sign3 = 4'd2;
b_sign0 = 4'd12; b_sign1 = 4'd0; b_sign2 = 4'd1; b_sign3 = 4'd12;
@(posedge clk_i);
a_mant0 = 8'd178; a_mant1 = 8'd24; a_mant2 = 8'd198; a_mant3 = 8'd28;
b_mant0 = 8'd241; b_mant1 = 8'd85; b_mant2 = 8'd35; b_mant3 = 8'd234;
a_exp0 = 10'd589; a_exp1 = 10'd31; a_exp2 = 10'd529; a_exp3 = 10'd995;
b_exp0 = 10'd671; b_exp1 = 10'd151; b_exp2 = 10'd1011; b_exp3 = 10'd148;
a_sign0 = 4'd13; a_sign1 = 4'd0; a_sign2 = 4'd4; a_sign3 = 4'd6;
b_sign0 = 4'd15; b_sign1 = 4'd1; b_sign2 = 4'd14; b_sign3 = 4'd1;
@(posedge clk_i);
a_mant0 = 8'd169; a_mant1 = 8'd68; a_mant2 = 8'd37; a_mant3 = 8'd61;
b_mant0 = 8'd32; b_mant1 = 8'd138; b_mant2 = 8'd103; b_mant3 = 8'd23;
a_exp0 = 10'd471; a_exp1 = 10'd979; a_exp2 = 10'd416; a_exp3 = 10'd429;
b_exp0 = 10'd660; b_exp1 = 10'd343; b_exp2 = 10'd540; b_exp3 = 10'd839;
a_sign0 = 4'd6; a_sign1 = 4'd6; a_sign2 = 4'd3; a_sign3 = 4'd3;
b_sign0 = 4'd9; b_sign1 = 4'd0; b_sign2 = 4'd12; b_sign3 = 4'd6;
@(posedge clk_i);
a_mant0 = 8'd123; a_mant1 = 8'd40; a_mant2 = 8'd195; a_mant3 = 8'd220;
b_mant0 = 8'd177; b_mant1 = 8'd176; b_mant2 = 8'd50; b_mant3 = 8'd255;
a_exp0 = 10'd586; a_exp1 = 10'd935; a_exp2 = 10'd13; a_exp3 = 10'd246;
b_exp0 = 10'd723; b_exp1 = 10'd61; b_exp2 = 10'd148; b_exp3 = 10'd534;
a_sign0 = 4'd16; a_sign1 = 4'd3; a_sign2 = 4'd12; a_sign3 = 4'd16;
b_sign0 = 4'd6; b_sign1 = 4'd13; b_sign2 = 4'd10; b_sign3 = 4'd1;
@(posedge clk_i);
shared_exps0 = 8'd142;
shared_exps1 = 8'd128;
a_mant0 = 8'd183; a_mant1 = 8'd137; a_mant2 = 8'd180; a_mant3 = 8'd164;
b_mant0 = 8'd44; b_mant1 = 8'd23; b_mant2 = 8'd144; b_mant3 = 8'd248;
a_exp0 = 10'd994; a_exp1 = 10'd895; a_exp2 = 10'd969; a_exp3 = 10'd47;
b_exp0 = 10'd981; b_exp1 = 10'd528; b_exp2 = 10'd813; b_exp3 = 10'd270;
a_sign0 = 4'd4; a_sign1 = 4'd15; a_sign2 = 4'd16; a_sign3 = 4'd6;
b_sign0 = 4'd0; b_sign1 = 4'd0; b_sign2 = 4'd4; b_sign3 = 4'd3;
@(posedge clk_i);
a_mant0 = 8'd41; a_mant1 = 8'd160; a_mant2 = 8'd91; a_mant3 = 8'd48;
b_mant0 = 8'd11; b_mant1 = 8'd93; b_mant2 = 8'd79; b_mant3 = 8'd207;
a_exp0 = 10'd244; a_exp1 = 10'd753; a_exp2 = 10'd67; a_exp3 = 10'd838;
b_exp0 = 10'd260; b_exp1 = 10'd772; b_exp2 = 10'd670; b_exp3 = 10'd166;
a_sign0 = 4'd2; a_sign1 = 4'd15; a_sign2 = 4'd9; a_sign3 = 4'd8;
b_sign0 = 4'd6; b_sign1 = 4'd8; b_sign2 = 4'd12; b_sign3 = 4'd3;
@(posedge clk_i);
a_mant0 = 8'd253; a_mant1 = 8'd63; a_mant2 = 8'd200; a_mant3 = 8'd121;
b_mant0 = 8'd152; b_mant1 = 8'd86; b_mant2 = 8'd163; b_mant3 = 8'd229;
a_exp0 = 10'd10; a_exp1 = 10'd409; a_exp2 = 10'd214; a_exp3 = 10'd61;
b_exp0 = 10'd462; b_exp1 = 10'd306; b_exp2 = 10'd290; b_exp3 = 10'd636;
a_sign0 = 4'd0; a_sign1 = 4'd3; a_sign2 = 4'd8; a_sign3 = 4'd12;
b_sign0 = 4'd6; b_sign1 = 4'd14; b_sign2 = 4'd2; b_sign3 = 4'd10;
@(posedge clk_i);
a_mant0 = 8'd38; a_mant1 = 8'd139; a_mant2 = 8'd51; a_mant3 = 8'd107;
b_mant0 = 8'd156; b_mant1 = 8'd138; b_mant2 = 8'd64; b_mant3 = 8'd222;
a_exp0 = 10'd654; a_exp1 = 10'd463; a_exp2 = 10'd382; a_exp3 = 10'd1016;
b_exp0 = 10'd932; b_exp1 = 10'd325; b_exp2 = 10'd508; b_exp3 = 10'd738;
a_sign0 = 4'd10; a_sign1 = 4'd15; a_sign2 = 4'd10; a_sign3 = 4'd13;
b_sign0 = 4'd11; b_sign1 = 4'd7; b_sign2 = 4'd9; b_sign3 = 4'd4;
@(posedge clk_i);
a_mant0 = 8'd180; a_mant1 = 8'd97; a_mant2 = 8'd97; a_mant3 = 8'd21;
b_mant0 = 8'd56; b_mant1 = 8'd175; b_mant2 = 8'd224; b_mant3 = 8'd202;
a_exp0 = 10'd505; a_exp1 = 10'd323; a_exp2 = 10'd114; a_exp3 = 10'd199;
b_exp0 = 10'd988; b_exp1 = 10'd293; b_exp2 = 10'd138; b_exp3 = 10'd232;
a_sign0 = 4'd4; a_sign1 = 4'd3; a_sign2 = 4'd10; a_sign3 = 4'd4;
b_sign0 = 4'd2; b_sign1 = 4'd1; b_sign2 = 4'd4; b_sign3 = 4'd12;
@(posedge clk_i);
a_mant0 = 8'd101; a_mant1 = 8'd56; a_mant2 = 8'd199; a_mant3 = 8'd151;
b_mant0 = 8'd160; b_mant1 = 8'd49; b_mant2 = 8'd231; b_mant3 = 8'd240;
a_exp0 = 10'd501; a_exp1 = 10'd649; a_exp2 = 10'd849; a_exp3 = 10'd260;
b_exp0 = 10'd216; b_exp1 = 10'd935; b_exp2 = 10'd756; b_exp3 = 10'd26;
a_sign0 = 4'd15; a_sign1 = 4'd4; a_sign2 = 4'd4; a_sign3 = 4'd12;
b_sign0 = 4'd11; b_sign1 = 4'd7; b_sign2 = 4'd0; b_sign3 = 4'd2;
@(posedge clk_i);
a_mant0 = 8'd57; a_mant1 = 8'd101; a_mant2 = 8'd32; a_mant3 = 8'd135;
b_mant0 = 8'd58; b_mant1 = 8'd219; b_mant2 = 8'd59; b_mant3 = 8'd8;
a_exp0 = 10'd158; a_exp1 = 10'd257; a_exp2 = 10'd185; a_exp3 = 10'd509;
b_exp0 = 10'd993; b_exp1 = 10'd587; b_exp2 = 10'd923; b_exp3 = 10'd816;
a_sign0 = 4'd6; a_sign1 = 4'd12; a_sign2 = 4'd13; a_sign3 = 4'd8;
b_sign0 = 4'd10; b_sign1 = 4'd9; b_sign2 = 4'd12; b_sign3 = 4'd4;
@(posedge clk_i);
a_mant0 = 8'd199; a_mant1 = 8'd243; a_mant2 = 8'd19; a_mant3 = 8'd10;
b_mant0 = 8'd37; b_mant1 = 8'd71; b_mant2 = 8'd72; b_mant3 = 8'd245;
a_exp0 = 10'd1004; a_exp1 = 10'd974; a_exp2 = 10'd30; a_exp3 = 10'd949;
b_exp0 = 10'd336; b_exp1 = 10'd878; b_exp2 = 10'd478; b_exp3 = 10'd452;
a_sign0 = 4'd10; a_sign1 = 4'd6; a_sign2 = 4'd6; a_sign3 = 4'd13;
b_sign0 = 4'd13; b_sign1 = 4'd15; b_sign2 = 4'd6; b_sign3 = 4'd15;
@(posedge clk_i);
shared_exps0 = 8'd125;
shared_exps1 = 8'd114;
a_mant0 = 8'd22; a_mant1 = 8'd31; a_mant2 = 8'd210; a_mant3 = 8'd223;
b_mant0 = 8'd144; b_mant1 = 8'd3; b_mant2 = 8'd97; b_mant3 = 8'd233;
a_exp0 = 10'd425; a_exp1 = 10'd509; a_exp2 = 10'd451; a_exp3 = 10'd573;
b_exp0 = 10'd475; b_exp1 = 10'd215; b_exp2 = 10'd485; b_exp3 = 10'd522;
a_sign0 = 4'd4; a_sign1 = 4'd2; a_sign2 = 4'd16; a_sign3 = 4'd6;
b_sign0 = 4'd0; b_sign1 = 4'd5; b_sign2 = 4'd12; b_sign3 = 4'd13;
@(posedge clk_i);
a_mant0 = 8'd253; a_mant1 = 8'd64; a_mant2 = 8'd163; a_mant3 = 8'd1;
b_mant0 = 8'd43; b_mant1 = 8'd5; b_mant2 = 8'd246; b_mant3 = 8'd66;
a_exp0 = 10'd221; a_exp1 = 10'd544; a_exp2 = 10'd673; a_exp3 = 10'd411;
b_exp0 = 10'd395; b_exp1 = 10'd695; b_exp2 = 10'd423; b_exp3 = 10'd200;
a_sign0 = 4'd4; a_sign1 = 4'd1; a_sign2 = 4'd3; a_sign3 = 4'd14;
b_sign0 = 4'd14; b_sign1 = 4'd3; b_sign2 = 4'd10; b_sign3 = 4'd13;
@(posedge clk_i);
a_mant0 = 8'd171; a_mant1 = 8'd193; a_mant2 = 8'd62; a_mant3 = 8'd29;
b_mant0 = 8'd221; b_mant1 = 8'd20; b_mant2 = 8'd125; b_mant3 = 8'd184;
a_exp0 = 10'd229; a_exp1 = 10'd10; a_exp2 = 10'd738; a_exp3 = 10'd565;
b_exp0 = 10'd792; b_exp1 = 10'd8; b_exp2 = 10'd164; b_exp3 = 10'd173;
a_sign0 = 4'd2; a_sign1 = 4'd12; a_sign2 = 4'd12; a_sign3 = 4'd2;
b_sign0 = 4'd11; b_sign1 = 4'd10; b_sign2 = 4'd16; b_sign3 = 4'd9;
@(posedge clk_i);
a_mant0 = 8'd228; a_mant1 = 8'd16; a_mant2 = 8'd153; a_mant3 = 8'd74;
b_mant0 = 8'd126; b_mant1 = 8'd207; b_mant2 = 8'd128; b_mant3 = 8'd85;
a_exp0 = 10'd744; a_exp1 = 10'd372; a_exp2 = 10'd363; a_exp3 = 10'd212;
b_exp0 = 10'd909; b_exp1 = 10'd240; b_exp2 = 10'd1018; b_exp3 = 10'd145;
a_sign0 = 4'd1; a_sign1 = 4'd7; a_sign2 = 4'd11; a_sign3 = 4'd15;
b_sign0 = 4'd0; b_sign1 = 4'd7; b_sign2 = 4'd0; b_sign3 = 4'd11;
@(posedge clk_i);
a_mant0 = 8'd123; a_mant1 = 8'd194; a_mant2 = 8'd22; a_mant3 = 8'd2;
b_mant0 = 8'd13; b_mant1 = 8'd185; b_mant2 = 8'd45; b_mant3 = 8'd162;
a_exp0 = 10'd895; a_exp1 = 10'd1017; a_exp2 = 10'd918; a_exp3 = 10'd720;
b_exp0 = 10'd960; b_exp1 = 10'd287; b_exp2 = 10'd72; b_exp3 = 10'd684;
a_sign0 = 4'd2; a_sign1 = 4'd12; a_sign2 = 4'd9; a_sign3 = 4'd2;
b_sign0 = 4'd4; b_sign1 = 4'd1; b_sign2 = 4'd4; b_sign3 = 4'd12;
@(posedge clk_i);
a_mant0 = 8'd28; a_mant1 = 8'd213; a_mant2 = 8'd161; a_mant3 = 8'd67;
b_mant0 = 8'd175; b_mant1 = 8'd136; b_mant2 = 8'd79; b_mant3 = 8'd167;
a_exp0 = 10'd515; a_exp1 = 10'd609; a_exp2 = 10'd186; a_exp3 = 10'd4;
b_exp0 = 10'd598; b_exp1 = 10'd1009; b_exp2 = 10'd401; b_exp3 = 10'd615;
a_sign0 = 4'd7; a_sign1 = 4'd8; a_sign2 = 4'd10; a_sign3 = 4'd1;
b_sign0 = 4'd13; b_sign1 = 4'd3; b_sign2 = 4'd0; b_sign3 = 4'd12;
@(posedge clk_i);
a_mant0 = 8'd101; a_mant1 = 8'd122; a_mant2 = 8'd111; a_mant3 = 8'd53;
b_mant0 = 8'd255; b_mant1 = 8'd103; b_mant2 = 8'd22; b_mant3 = 8'd208;
a_exp0 = 10'd806; a_exp1 = 10'd908; a_exp2 = 10'd726; a_exp3 = 10'd926;
b_exp0 = 10'd943; b_exp1 = 10'd823; b_exp2 = 10'd917; b_exp3 = 10'd136;
a_sign0 = 4'd11; a_sign1 = 4'd3; a_sign2 = 4'd4; a_sign3 = 4'd8;
b_sign0 = 4'd4; b_sign1 = 4'd5; b_sign2 = 4'd12; b_sign3 = 4'd7;
@(posedge clk_i);
a_mant0 = 8'd66; a_mant1 = 8'd197; a_mant2 = 8'd219; a_mant3 = 8'd79;
b_mant0 = 8'd44; b_mant1 = 8'd105; b_mant2 = 8'd66; b_mant3 = 8'd22;
a_exp0 = 10'd467; a_exp1 = 10'd351; a_exp2 = 10'd609; a_exp3 = 10'd912;
b_exp0 = 10'd705; b_exp1 = 10'd41; b_exp2 = 10'd713; b_exp3 = 10'd49;
a_sign0 = 4'd0; a_sign1 = 4'd3; a_sign2 = 4'd9; a_sign3 = 4'd5;
b_sign0 = 4'd7; b_sign1 = 4'd10; b_sign2 = 4'd8; b_sign3 = 4'd15;
@(posedge clk_i);
shared_exps0 = 8'd125;
shared_exps1 = 8'd126;
a_mant0 = 8'd142; a_mant1 = 8'd232; a_mant2 = 8'd4; a_mant3 = 8'd191;
b_mant0 = 8'd54; b_mant1 = 8'd151; b_mant2 = 8'd10; b_mant3 = 8'd191;
a_exp0 = 10'd341; a_exp1 = 10'd309; a_exp2 = 10'd239; a_exp3 = 10'd421;
b_exp0 = 10'd944; b_exp1 = 10'd1014; b_exp2 = 10'd83; b_exp3 = 10'd75;
a_sign0 = 4'd15; a_sign1 = 4'd1; a_sign2 = 4'd14; a_sign3 = 4'd3;
b_sign0 = 4'd6; b_sign1 = 4'd10; b_sign2 = 4'd1; b_sign3 = 4'd16;
@(posedge clk_i);
a_mant0 = 8'd97; a_mant1 = 8'd231; a_mant2 = 8'd176; a_mant3 = 8'd163;
b_mant0 = 8'd240; b_mant1 = 8'd31; b_mant2 = 8'd184; b_mant3 = 8'd124;
a_exp0 = 10'd948; a_exp1 = 10'd663; a_exp2 = 10'd104; a_exp3 = 10'd811;
b_exp0 = 10'd239; b_exp1 = 10'd257; b_exp2 = 10'd984; b_exp3 = 10'd706;
a_sign0 = 4'd15; a_sign1 = 4'd16; a_sign2 = 4'd2; a_sign3 = 4'd8;
b_sign0 = 4'd11; b_sign1 = 4'd6; b_sign2 = 4'd16; b_sign3 = 4'd10;
@(posedge clk_i);
a_mant0 = 8'd162; a_mant1 = 8'd119; a_mant2 = 8'd62; a_mant3 = 8'd11;
b_mant0 = 8'd247; b_mant1 = 8'd68; b_mant2 = 8'd178; b_mant3 = 8'd16;
a_exp0 = 10'd49; a_exp1 = 10'd508; a_exp2 = 10'd486; a_exp3 = 10'd305;
b_exp0 = 10'd956; b_exp1 = 10'd814; b_exp2 = 10'd67; b_exp3 = 10'd484;
a_sign0 = 4'd7; a_sign1 = 4'd0; a_sign2 = 4'd12; a_sign3 = 4'd6;
b_sign0 = 4'd8; b_sign1 = 4'd15; b_sign2 = 4'd14; b_sign3 = 4'd1;
@(posedge clk_i);
a_mant0 = 8'd129; a_mant1 = 8'd150; a_mant2 = 8'd42; a_mant3 = 8'd206;
b_mant0 = 8'd162; b_mant1 = 8'd246; b_mant2 = 8'd77; b_mant3 = 8'd41;
a_exp0 = 10'd689; a_exp1 = 10'd710; a_exp2 = 10'd37; a_exp3 = 10'd817;
b_exp0 = 10'd767; b_exp1 = 10'd351; b_exp2 = 10'd873; b_exp3 = 10'd261;
a_sign0 = 4'd12; a_sign1 = 4'd1; a_sign2 = 4'd6; a_sign3 = 4'd4;
b_sign0 = 4'd8; b_sign1 = 4'd13; b_sign2 = 4'd15; b_sign3 = 4'd11;
@(posedge clk_i);
a_mant0 = 8'd49; a_mant1 = 8'd250; a_mant2 = 8'd140; a_mant3 = 8'd81;
b_mant0 = 8'd92; b_mant1 = 8'd83; b_mant2 = 8'd234; b_mant3 = 8'd190;
a_exp0 = 10'd32; a_exp1 = 10'd923; a_exp2 = 10'd409; a_exp3 = 10'd709;
b_exp0 = 10'd113; b_exp1 = 10'd673; b_exp2 = 10'd388; b_exp3 = 10'd420;
a_sign0 = 4'd7; a_sign1 = 4'd12; a_sign2 = 4'd16; a_sign3 = 4'd13;
b_sign0 = 4'd2; b_sign1 = 4'd16; b_sign2 = 4'd6; b_sign3 = 4'd9;
@(posedge clk_i);
a_mant0 = 8'd255; a_mant1 = 8'd102; a_mant2 = 8'd123; a_mant3 = 8'd113;
b_mant0 = 8'd52; b_mant1 = 8'd240; b_mant2 = 8'd34; b_mant3 = 8'd110;
a_exp0 = 10'd914; a_exp1 = 10'd795; a_exp2 = 10'd995; a_exp3 = 10'd82;
b_exp0 = 10'd108; b_exp1 = 10'd840; b_exp2 = 10'd299; b_exp3 = 10'd480;
a_sign0 = 4'd12; a_sign1 = 4'd7; a_sign2 = 4'd16; a_sign3 = 4'd3;
b_sign0 = 4'd0; b_sign1 = 4'd13; b_sign2 = 4'd16; b_sign3 = 4'd3;
@(posedge clk_i);
a_mant0 = 8'd251; a_mant1 = 8'd204; a_mant2 = 8'd184; a_mant3 = 8'd219;
b_mant0 = 8'd104; b_mant1 = 8'd235; b_mant2 = 8'd222; b_mant3 = 8'd145;
a_exp0 = 10'd318; a_exp1 = 10'd829; a_exp2 = 10'd125; a_exp3 = 10'd18;
b_exp0 = 10'd183; b_exp1 = 10'd808; b_exp2 = 10'd336; b_exp3 = 10'd960;
a_sign0 = 4'd6; a_sign1 = 4'd4; a_sign2 = 4'd6; a_sign3 = 4'd2;
b_sign0 = 4'd5; b_sign1 = 4'd10; b_sign2 = 4'd5; b_sign3 = 4'd1;
@(posedge clk_i);
a_mant0 = 8'd91; a_mant1 = 8'd142; a_mant2 = 8'd85; a_mant3 = 8'd176;
b_mant0 = 8'd96; b_mant1 = 8'd82; b_mant2 = 8'd34; b_mant3 = 8'd185;
a_exp0 = 10'd982; a_exp1 = 10'd217; a_exp2 = 10'd945; a_exp3 = 10'd573;
b_exp0 = 10'd144; b_exp1 = 10'd82; b_exp2 = 10'd495; b_exp3 = 10'd662;
a_sign0 = 4'd16; a_sign1 = 4'd2; a_sign2 = 4'd5; a_sign3 = 4'd1;
b_sign0 = 4'd16; b_sign1 = 4'd11; b_sign2 = 4'd10; b_sign3 = 4'd6;
@(posedge clk_i);
shared_exps0 = 8'd144;
shared_exps1 = 8'd122;
rstn = 0;
@(posedge clk_i);
rstn = 1;
a_mant0 = 8'd239; a_mant1 = 8'd73; a_mant2 = 8'd113; a_mant3 = 8'd53;
b_mant0 = 8'd13; b_mant1 = 8'd240; b_mant2 = 8'd98; b_mant3 = 8'd200;
a_exp0 = 10'd885; a_exp1 = 10'd842; a_exp2 = 10'd39; a_exp3 = 10'd801;
b_exp0 = 10'd120; b_exp1 = 10'd479; b_exp2 = 10'd609; b_exp3 = 10'd408;
a_sign0 = 4'd16; a_sign1 = 4'd4; a_sign2 = 4'd7; a_sign3 = 4'd0;
b_sign0 = 4'd11; b_sign1 = 4'd13; b_sign2 = 4'd4; b_sign3 = 4'd10;
@(posedge clk_i);
a_mant0 = 8'd73; a_mant1 = 8'd165; a_mant2 = 8'd85; a_mant3 = 8'd102;
b_mant0 = 8'd14; b_mant1 = 8'd194; b_mant2 = 8'd31; b_mant3 = 8'd5;
a_exp0 = 10'd595; a_exp1 = 10'd363; a_exp2 = 10'd1019; a_exp3 = 10'd341;
b_exp0 = 10'd708; b_exp1 = 10'd163; b_exp2 = 10'd106; b_exp3 = 10'd480;
a_sign0 = 4'd12; a_sign1 = 4'd13; a_sign2 = 4'd1; a_sign3 = 4'd2;
b_sign0 = 4'd11; b_sign1 = 4'd2; b_sign2 = 4'd12; b_sign3 = 4'd2;
@(posedge clk_i);
a_mant0 = 8'd246; a_mant1 = 8'd209; a_mant2 = 8'd250; a_mant3 = 8'd93;
b_mant0 = 8'd102; b_mant1 = 8'd78; b_mant2 = 8'd17; b_mant3 = 8'd163;
a_exp0 = 10'd1013; a_exp1 = 10'd739; a_exp2 = 10'd912; a_exp3 = 10'd1012;
b_exp0 = 10'd582; b_exp1 = 10'd556; b_exp2 = 10'd869; b_exp3 = 10'd405;
a_sign0 = 4'd11; a_sign1 = 4'd10; a_sign2 = 4'd10; a_sign3 = 4'd14;
b_sign0 = 4'd16; b_sign1 = 4'd9; b_sign2 = 4'd1; b_sign3 = 4'd2;
@(posedge clk_i);
a_mant0 = 8'd11; a_mant1 = 8'd240; a_mant2 = 8'd57; a_mant3 = 8'd50;
b_mant0 = 8'd166; b_mant1 = 8'd159; b_mant2 = 8'd184; b_mant3 = 8'd171;
a_exp0 = 10'd289; a_exp1 = 10'd581; a_exp2 = 10'd886; a_exp3 = 10'd397;
b_exp0 = 10'd488; b_exp1 = 10'd750; b_exp2 = 10'd849; b_exp3 = 10'd389;
a_sign0 = 4'd0; a_sign1 = 4'd0; a_sign2 = 4'd12; a_sign3 = 4'd12;
b_sign0 = 4'd10; b_sign1 = 4'd14; b_sign2 = 4'd11; b_sign3 = 4'd2;
@(posedge clk_i);
a_mant0 = 8'd224; a_mant1 = 8'd95; a_mant2 = 8'd140; a_mant3 = 8'd84;
b_mant0 = 8'd9; b_mant1 = 8'd53; b_mant2 = 8'd73; b_mant3 = 8'd146;
a_exp0 = 10'd189; a_exp1 = 10'd927; a_exp2 = 10'd958; a_exp3 = 10'd574;
b_exp0 = 10'd323; b_exp1 = 10'd118; b_exp2 = 10'd617; b_exp3 = 10'd841;
a_sign0 = 4'd10; a_sign1 = 4'd4; a_sign2 = 4'd11; a_sign3 = 4'd5;
b_sign0 = 4'd9; b_sign1 = 4'd12; b_sign2 = 4'd13; b_sign3 = 4'd1;
@(posedge clk_i);
a_mant0 = 8'd38; a_mant1 = 8'd86; a_mant2 = 8'd148; a_mant3 = 8'd27;
b_mant0 = 8'd246; b_mant1 = 8'd174; b_mant2 = 8'd179; b_mant3 = 8'd84;
a_exp0 = 10'd752; a_exp1 = 10'd731; a_exp2 = 10'd462; a_exp3 = 10'd816;
b_exp0 = 10'd196; b_exp1 = 10'd956; b_exp2 = 10'd227; b_exp3 = 10'd0;
a_sign0 = 4'd2; a_sign1 = 4'd16; a_sign2 = 4'd12; a_sign3 = 4'd15;
b_sign0 = 4'd4; b_sign1 = 4'd9; b_sign2 = 4'd2; b_sign3 = 4'd4;
@(posedge clk_i);
a_mant0 = 8'd19; a_mant1 = 8'd216; a_mant2 = 8'd91; a_mant3 = 8'd56;
b_mant0 = 8'd99; b_mant1 = 8'd9; b_mant2 = 8'd223; b_mant3 = 8'd200;
a_exp0 = 10'd382; a_exp1 = 10'd499; a_exp2 = 10'd684; a_exp3 = 10'd961;
b_exp0 = 10'd468; b_exp1 = 10'd585; b_exp2 = 10'd637; b_exp3 = 10'd812;
a_sign0 = 4'd0; a_sign1 = 4'd12; a_sign2 = 4'd15; a_sign3 = 4'd15;
b_sign0 = 4'd16; b_sign1 = 4'd13; b_sign2 = 4'd1; b_sign3 = 4'd15;
@(posedge clk_i);
shared_exps0 = 8'd118;
shared_exps1 = 8'd108;
a_mant0 = 8'd111; a_mant1 = 8'd8; a_mant2 = 8'd24; a_mant3 = 8'd238;
b_mant0 = 8'd111; b_mant1 = 8'd10; b_mant2 = 8'd184; b_mant3 = 8'd15;
a_exp0 = 10'd487; a_exp1 = 10'd1013; a_exp2 = 10'd24; a_exp3 = 10'd813;
b_exp0 = 10'd910; b_exp1 = 10'd111; b_exp2 = 10'd408; b_exp3 = 10'd797;
a_sign0 = 4'd13; a_sign1 = 4'd11; a_sign2 = 4'd16; a_sign3 = 4'd12;
b_sign0 = 4'd10; b_sign1 = 4'd15; b_sign2 = 4'd7; b_sign3 = 4'd3;
@(posedge clk_i);
a_mant0 = 8'd36; a_mant1 = 8'd186; a_mant2 = 8'd254; a_mant3 = 8'd74;
b_mant0 = 8'd27; b_mant1 = 8'd68; b_mant2 = 8'd141; b_mant3 = 8'd62;
a_exp0 = 10'd253; a_exp1 = 10'd225; a_exp2 = 10'd758; a_exp3 = 10'd665;
b_exp0 = 10'd790; b_exp1 = 10'd135; b_exp2 = 10'd590; b_exp3 = 10'd806;
a_sign0 = 4'd8; a_sign1 = 4'd1; a_sign2 = 4'd6; a_sign3 = 4'd12;
b_sign0 = 4'd10; b_sign1 = 4'd6; b_sign2 = 4'd7; b_sign3 = 4'd0;
@(posedge clk_i);
a_mant0 = 8'd25; a_mant1 = 8'd254; a_mant2 = 8'd165; a_mant3 = 8'd234;
b_mant0 = 8'd80; b_mant1 = 8'd64; b_mant2 = 8'd250; b_mant3 = 8'd228;
a_exp0 = 10'd811; a_exp1 = 10'd413; a_exp2 = 10'd205; a_exp3 = 10'd816;
b_exp0 = 10'd754; b_exp1 = 10'd53; b_exp2 = 10'd783; b_exp3 = 10'd664;
a_sign0 = 4'd13; a_sign1 = 4'd5; a_sign2 = 4'd0; a_sign3 = 4'd16;
b_sign0 = 4'd12; b_sign1 = 4'd7; b_sign2 = 4'd10; b_sign3 = 4'd14;
@(posedge clk_i);
a_mant0 = 8'd203; a_mant1 = 8'd108; a_mant2 = 8'd140; a_mant3 = 8'd203;
b_mant0 = 8'd152; b_mant1 = 8'd207; b_mant2 = 8'd68; b_mant3 = 8'd243;
a_exp0 = 10'd942; a_exp1 = 10'd393; a_exp2 = 10'd239; a_exp3 = 10'd900;
b_exp0 = 10'd253; b_exp1 = 10'd209; b_exp2 = 10'd209; b_exp3 = 10'd223;
a_sign0 = 4'd14; a_sign1 = 4'd1; a_sign2 = 4'd12; a_sign3 = 4'd4;
b_sign0 = 4'd15; b_sign1 = 4'd14; b_sign2 = 4'd1; b_sign3 = 4'd2;
@(posedge clk_i);
a_mant0 = 8'd97; a_mant1 = 8'd107; a_mant2 = 8'd87; a_mant3 = 8'd165;
b_mant0 = 8'd154; b_mant1 = 8'd190; b_mant2 = 8'd154; b_mant3 = 8'd101;
a_exp0 = 10'd409; a_exp1 = 10'd801; a_exp2 = 10'd410; a_exp3 = 10'd507;
b_exp0 = 10'd637; b_exp1 = 10'd443; b_exp2 = 10'd55; b_exp3 = 10'd969;
a_sign0 = 4'd3; a_sign1 = 4'd10; a_sign2 = 4'd5; a_sign3 = 4'd7;
b_sign0 = 4'd8; b_sign1 = 4'd4; b_sign2 = 4'd3; b_sign3 = 4'd5;
@(posedge clk_i);
a_mant0 = 8'd23; a_mant1 = 8'd255; a_mant2 = 8'd108; a_mant3 = 8'd173;
b_mant0 = 8'd7; b_mant1 = 8'd39; b_mant2 = 8'd222; b_mant3 = 8'd62;
a_exp0 = 10'd555; a_exp1 = 10'd559; a_exp2 = 10'd155; a_exp3 = 10'd285;
b_exp0 = 10'd573; b_exp1 = 10'd104; b_exp2 = 10'd362; b_exp3 = 10'd10;
a_sign0 = 4'd10; a_sign1 = 4'd6; a_sign2 = 4'd10; a_sign3 = 4'd9;
b_sign0 = 4'd8; b_sign1 = 4'd3; b_sign2 = 4'd15; b_sign3 = 4'd13;
@(posedge clk_i);
a_mant0 = 8'd123; a_mant1 = 8'd36; a_mant2 = 8'd149; a_mant3 = 8'd111;
b_mant0 = 8'd4; b_mant1 = 8'd180; b_mant2 = 8'd38; b_mant3 = 8'd225;
a_exp0 = 10'd253; a_exp1 = 10'd731; a_exp2 = 10'd289; a_exp3 = 10'd74;
b_exp0 = 10'd117; b_exp1 = 10'd969; b_exp2 = 10'd205; b_exp3 = 10'd691;
a_sign0 = 4'd14; a_sign1 = 4'd1; a_sign2 = 4'd12; a_sign3 = 4'd5;
b_sign0 = 4'd6; b_sign1 = 4'd13; b_sign2 = 4'd10; b_sign3 = 4'd11;
@(posedge clk_i);
a_mant0 = 8'd247; a_mant1 = 8'd200; a_mant2 = 8'd135; a_mant3 = 8'd158;
b_mant0 = 8'd144; b_mant1 = 8'd249; b_mant2 = 8'd223; b_mant3 = 8'd11;
a_exp0 = 10'd362; a_exp1 = 10'd255; a_exp2 = 10'd213; a_exp3 = 10'd485;
b_exp0 = 10'd1005; b_exp1 = 10'd910; b_exp2 = 10'd475; b_exp3 = 10'd389;
a_sign0 = 4'd6; a_sign1 = 4'd4; a_sign2 = 4'd7; a_sign3 = 4'd14;
b_sign0 = 4'd2; b_sign1 = 4'd10; b_sign2 = 4'd7; b_sign3 = 4'd15;
@(posedge clk_i);
shared_exps0 = 8'd143;
shared_exps1 = 8'd129;
a_mant0 = 8'd182; a_mant1 = 8'd27; a_mant2 = 8'd35; a_mant3 = 8'd164;
b_mant0 = 8'd98; b_mant1 = 8'd11; b_mant2 = 8'd102; b_mant3 = 8'd15;
a_exp0 = 10'd179; a_exp1 = 10'd429; a_exp2 = 10'd311; a_exp3 = 10'd539;
b_exp0 = 10'd445; b_exp1 = 10'd575; b_exp2 = 10'd36; b_exp3 = 10'd882;
a_sign0 = 4'd4; a_sign1 = 4'd13; a_sign2 = 4'd9; a_sign3 = 4'd16;
b_sign0 = 4'd3; b_sign1 = 4'd8; b_sign2 = 4'd6; b_sign3 = 4'd7;
@(posedge clk_i);
a_mant0 = 8'd100; a_mant1 = 8'd81; a_mant2 = 8'd174; a_mant3 = 8'd121;
b_mant0 = 8'd249; b_mant1 = 8'd157; b_mant2 = 8'd223; b_mant3 = 8'd67;
a_exp0 = 10'd449; a_exp1 = 10'd263; a_exp2 = 10'd98; a_exp3 = 10'd1015;
b_exp0 = 10'd263; b_exp1 = 10'd75; b_exp2 = 10'd842; b_exp3 = 10'd509;
a_sign0 = 4'd10; a_sign1 = 4'd3; a_sign2 = 4'd0; a_sign3 = 4'd11;
b_sign0 = 4'd4; b_sign1 = 4'd5; b_sign2 = 4'd11; b_sign3 = 4'd8;
@(posedge clk_i);
a_mant0 = 8'd161; a_mant1 = 8'd142; a_mant2 = 8'd14; a_mant3 = 8'd92;
b_mant0 = 8'd80; b_mant1 = 8'd72; b_mant2 = 8'd18; b_mant3 = 8'd205;
a_exp0 = 10'd422; a_exp1 = 10'd240; a_exp2 = 10'd107; a_exp3 = 10'd642;
b_exp0 = 10'd204; b_exp1 = 10'd304; b_exp2 = 10'd1019; b_exp3 = 10'd472;
a_sign0 = 4'd5; a_sign1 = 4'd9; a_sign2 = 4'd11; a_sign3 = 4'd9;
b_sign0 = 4'd16; b_sign1 = 4'd10; b_sign2 = 4'd6; b_sign3 = 4'd11;
@(posedge clk_i);
a_mant0 = 8'd189; a_mant1 = 8'd250; a_mant2 = 8'd53; a_mant3 = 8'd98;
b_mant0 = 8'd61; b_mant1 = 8'd102; b_mant2 = 8'd72; b_mant3 = 8'd220;
a_exp0 = 10'd178; a_exp1 = 10'd307; a_exp2 = 10'd749; a_exp3 = 10'd1022;
b_exp0 = 10'd369; b_exp1 = 10'd312; b_exp2 = 10'd596; b_exp3 = 10'd706;
a_sign0 = 4'd9; a_sign1 = 4'd16; a_sign2 = 4'd1; a_sign3 = 4'd6;
b_sign0 = 4'd8; b_sign1 = 4'd3; b_sign2 = 4'd15; b_sign3 = 4'd6;
@(posedge clk_i);
a_mant0 = 8'd59; a_mant1 = 8'd74; a_mant2 = 8'd177; a_mant3 = 8'd1;
b_mant0 = 8'd140; b_mant1 = 8'd145; b_mant2 = 8'd230; b_mant3 = 8'd211;
a_exp0 = 10'd535; a_exp1 = 10'd261; a_exp2 = 10'd319; a_exp3 = 10'd438;
b_exp0 = 10'd25; b_exp1 = 10'd184; b_exp2 = 10'd160; b_exp3 = 10'd483;
a_sign0 = 4'd12; a_sign1 = 4'd0; a_sign2 = 4'd3; a_sign3 = 4'd5;
b_sign0 = 4'd11; b_sign1 = 4'd2; b_sign2 = 4'd15; b_sign3 = 4'd4;
@(posedge clk_i);
a_mant0 = 8'd110; a_mant1 = 8'd244; a_mant2 = 8'd91; a_mant3 = 8'd163;
b_mant0 = 8'd177; b_mant1 = 8'd170; b_mant2 = 8'd97; b_mant3 = 8'd200;
a_exp0 = 10'd576; a_exp1 = 10'd591; a_exp2 = 10'd897; a_exp3 = 10'd487;
b_exp0 = 10'd485; b_exp1 = 10'd272; b_exp2 = 10'd756; b_exp3 = 10'd168;
a_sign0 = 4'd11; a_sign1 = 4'd2; a_sign2 = 4'd6; a_sign3 = 4'd13;
b_sign0 = 4'd15; b_sign1 = 4'd7; b_sign2 = 4'd13; b_sign3 = 4'd0;
@(posedge clk_i);
a_mant0 = 8'd137; a_mant1 = 8'd172; a_mant2 = 8'd194; a_mant3 = 8'd114;
b_mant0 = 8'd200; b_mant1 = 8'd216; b_mant2 = 8'd0; b_mant3 = 8'd163;
a_exp0 = 10'd442; a_exp1 = 10'd885; a_exp2 = 10'd694; a_exp3 = 10'd889;
b_exp0 = 10'd333; b_exp1 = 10'd890; b_exp2 = 10'd511; b_exp3 = 10'd817;
a_sign0 = 4'd12; a_sign1 = 4'd0; a_sign2 = 4'd13; a_sign3 = 4'd2;
b_sign0 = 4'd7; b_sign1 = 4'd15; b_sign2 = 4'd0; b_sign3 = 4'd1;
@(posedge clk_i);
a_mant0 = 8'd4; a_mant1 = 8'd154; a_mant2 = 8'd206; a_mant3 = 8'd142;
b_mant0 = 8'd146; b_mant1 = 8'd223; b_mant2 = 8'd182; b_mant3 = 8'd57;
a_exp0 = 10'd247; a_exp1 = 10'd1003; a_exp2 = 10'd290; a_exp3 = 10'd825;
b_exp0 = 10'd235; b_exp1 = 10'd143; b_exp2 = 10'd403; b_exp3 = 10'd642;
a_sign0 = 4'd7; a_sign1 = 4'd9; a_sign2 = 4'd5; a_sign3 = 4'd3;
b_sign0 = 4'd3; b_sign1 = 4'd9; b_sign2 = 4'd5; b_sign3 = 4'd4;
@(posedge clk_i);
shared_exps0 = 8'd127;
shared_exps1 = 8'd108;
a_mant0 = 8'd65; a_mant1 = 8'd246; a_mant2 = 8'd35; a_mant3 = 8'd70;
b_mant0 = 8'd133; b_mant1 = 8'd223; b_mant2 = 8'd54; b_mant3 = 8'd124;
a_exp0 = 10'd229; a_exp1 = 10'd30; a_exp2 = 10'd685; a_exp3 = 10'd90;
b_exp0 = 10'd684; b_exp1 = 10'd84; b_exp2 = 10'd202; b_exp3 = 10'd980;
a_sign0 = 4'd8; a_sign1 = 4'd13; a_sign2 = 4'd3; a_sign3 = 4'd8;
b_sign0 = 4'd6; b_sign1 = 4'd11; b_sign2 = 4'd2; b_sign3 = 4'd8;
@(posedge clk_i);
a_mant0 = 8'd93; a_mant1 = 8'd142; a_mant2 = 8'd175; a_mant3 = 8'd122;
b_mant0 = 8'd2; b_mant1 = 8'd113; b_mant2 = 8'd40; b_mant3 = 8'd7;
a_exp0 = 10'd842; a_exp1 = 10'd93; a_exp2 = 10'd160; a_exp3 = 10'd174;
b_exp0 = 10'd717; b_exp1 = 10'd654; b_exp2 = 10'd979; b_exp3 = 10'd688;
a_sign0 = 4'd5; a_sign1 = 4'd14; a_sign2 = 4'd2; a_sign3 = 4'd2;
b_sign0 = 4'd4; b_sign1 = 4'd7; b_sign2 = 4'd5; b_sign3 = 4'd12;
@(posedge clk_i);
a_mant0 = 8'd111; a_mant1 = 8'd65; a_mant2 = 8'd194; a_mant3 = 8'd182;
b_mant0 = 8'd44; b_mant1 = 8'd178; b_mant2 = 8'd19; b_mant3 = 8'd206;
a_exp0 = 10'd17; a_exp1 = 10'd723; a_exp2 = 10'd866; a_exp3 = 10'd842;
b_exp0 = 10'd132; b_exp1 = 10'd350; b_exp2 = 10'd826; b_exp3 = 10'd237;
a_sign0 = 4'd13; a_sign1 = 4'd11; a_sign2 = 4'd6; a_sign3 = 4'd13;
b_sign0 = 4'd15; b_sign1 = 4'd11; b_sign2 = 4'd14; b_sign3 = 4'd9;
@(posedge clk_i);
a_mant0 = 8'd209; a_mant1 = 8'd164; a_mant2 = 8'd121; a_mant3 = 8'd8;
b_mant0 = 8'd126; b_mant1 = 8'd7; b_mant2 = 8'd51; b_mant3 = 8'd179;
a_exp0 = 10'd730; a_exp1 = 10'd380; a_exp2 = 10'd1002; a_exp3 = 10'd634;
b_exp0 = 10'd253; b_exp1 = 10'd800; b_exp2 = 10'd464; b_exp3 = 10'd347;
a_sign0 = 4'd14; a_sign1 = 4'd0; a_sign2 = 4'd4; a_sign3 = 4'd6;
b_sign0 = 4'd2; b_sign1 = 4'd15; b_sign2 = 4'd15; b_sign3 = 4'd8;
@(posedge clk_i);
a_mant0 = 8'd97; a_mant1 = 8'd249; a_mant2 = 8'd2; a_mant3 = 8'd214;
b_mant0 = 8'd130; b_mant1 = 8'd84; b_mant2 = 8'd216; b_mant3 = 8'd168;
a_exp0 = 10'd340; a_exp1 = 10'd255; a_exp2 = 10'd552; a_exp3 = 10'd613;
b_exp0 = 10'd461; b_exp1 = 10'd995; b_exp2 = 10'd219; b_exp3 = 10'd639;
a_sign0 = 4'd10; a_sign1 = 4'd3; a_sign2 = 4'd14; a_sign3 = 4'd7;
b_sign0 = 4'd12; b_sign1 = 4'd16; b_sign2 = 4'd2; b_sign3 = 4'd8;
@(posedge clk_i);
a_mant0 = 8'd105; a_mant1 = 8'd16; a_mant2 = 8'd38; a_mant3 = 8'd215;
b_mant0 = 8'd239; b_mant1 = 8'd46; b_mant2 = 8'd160; b_mant3 = 8'd131;
a_exp0 = 10'd445; a_exp1 = 10'd428; a_exp2 = 10'd800; a_exp3 = 10'd647;
b_exp0 = 10'd448; b_exp1 = 10'd665; b_exp2 = 10'd452; b_exp3 = 10'd203;
a_sign0 = 4'd13; a_sign1 = 4'd4; a_sign2 = 4'd7; a_sign3 = 4'd4;
b_sign0 = 4'd5; b_sign1 = 4'd13; b_sign2 = 4'd2; b_sign3 = 4'd15;
@(posedge clk_i);
a_mant0 = 8'd165; a_mant1 = 8'd86; a_mant2 = 8'd235; a_mant3 = 8'd251;
b_mant0 = 8'd246; b_mant1 = 8'd229; b_mant2 = 8'd116; b_mant3 = 8'd55;
a_exp0 = 10'd756; a_exp1 = 10'd69; a_exp2 = 10'd130; a_exp3 = 10'd131;
b_exp0 = 10'd731; b_exp1 = 10'd405; b_exp2 = 10'd636; b_exp3 = 10'd195;
a_sign0 = 4'd11; a_sign1 = 4'd2; a_sign2 = 4'd2; a_sign3 = 4'd13;
b_sign0 = 4'd4; b_sign1 = 4'd11; b_sign2 = 4'd3; b_sign3 = 4'd0;
@(posedge clk_i);
a_mant0 = 8'd175; a_mant1 = 8'd253; a_mant2 = 8'd152; a_mant3 = 8'd149;
b_mant0 = 8'd18; b_mant1 = 8'd90; b_mant2 = 8'd244; b_mant3 = 8'd9;
a_exp0 = 10'd674; a_exp1 = 10'd234; a_exp2 = 10'd757; a_exp3 = 10'd693;
b_exp0 = 10'd256; b_exp1 = 10'd140; b_exp2 = 10'd404; b_exp3 = 10'd724;
a_sign0 = 4'd14; a_sign1 = 4'd5; a_sign2 = 4'd9; a_sign3 = 4'd11;
b_sign0 = 4'd5; b_sign1 = 4'd3; b_sign2 = 4'd5; b_sign3 = 4'd11;
@(posedge clk_i);
shared_exps0 = 8'd110;
shared_exps1 = 8'd108;
rstn = 0;
@(posedge clk_i);
rstn = 1;
a_mant0 = 8'd163; a_mant1 = 8'd81; a_mant2 = 8'd105; a_mant3 = 8'd20;
b_mant0 = 8'd225; b_mant1 = 8'd82; b_mant2 = 8'd209; b_mant3 = 8'd49;
a_exp0 = 10'd308; a_exp1 = 10'd814; a_exp2 = 10'd114; a_exp3 = 10'd305;
b_exp0 = 10'd584; b_exp1 = 10'd237; b_exp2 = 10'd777; b_exp3 = 10'd230;
a_sign0 = 4'd16; a_sign1 = 4'd15; a_sign2 = 4'd1; a_sign3 = 4'd14;
b_sign0 = 4'd11; b_sign1 = 4'd15; b_sign2 = 4'd2; b_sign3 = 4'd16;
@(posedge clk_i);
a_mant0 = 8'd152; a_mant1 = 8'd18; a_mant2 = 8'd107; a_mant3 = 8'd230;
b_mant0 = 8'd93; b_mant1 = 8'd57; b_mant2 = 8'd202; b_mant3 = 8'd252;
a_exp0 = 10'd549; a_exp1 = 10'd844; a_exp2 = 10'd280; a_exp3 = 10'd50;
b_exp0 = 10'd579; b_exp1 = 10'd811; b_exp2 = 10'd241; b_exp3 = 10'd269;
a_sign0 = 4'd5; a_sign1 = 4'd10; a_sign2 = 4'd16; a_sign3 = 4'd0;
b_sign0 = 4'd9; b_sign1 = 4'd5; b_sign2 = 4'd1; b_sign3 = 4'd10;
@(posedge clk_i);
a_mant0 = 8'd58; a_mant1 = 8'd245; a_mant2 = 8'd31; a_mant3 = 8'd85;
b_mant0 = 8'd47; b_mant1 = 8'd219; b_mant2 = 8'd28; b_mant3 = 8'd81;
a_exp0 = 10'd227; a_exp1 = 10'd442; a_exp2 = 10'd372; a_exp3 = 10'd456;
b_exp0 = 10'd522; b_exp1 = 10'd835; b_exp2 = 10'd763; b_exp3 = 10'd736;
a_sign0 = 4'd11; a_sign1 = 4'd15; a_sign2 = 4'd7; a_sign3 = 4'd15;
b_sign0 = 4'd14; b_sign1 = 4'd16; b_sign2 = 4'd10; b_sign3 = 4'd1;
@(posedge clk_i);
a_mant0 = 8'd44; a_mant1 = 8'd85; a_mant2 = 8'd202; a_mant3 = 8'd139;
b_mant0 = 8'd228; b_mant1 = 8'd12; b_mant2 = 8'd183; b_mant3 = 8'd159;
a_exp0 = 10'd282; a_exp1 = 10'd142; a_exp2 = 10'd9; a_exp3 = 10'd641;
b_exp0 = 10'd696; b_exp1 = 10'd672; b_exp2 = 10'd610; b_exp3 = 10'd771;
a_sign0 = 4'd3; a_sign1 = 4'd13; a_sign2 = 4'd8; a_sign3 = 4'd11;
b_sign0 = 4'd8; b_sign1 = 4'd2; b_sign2 = 4'd11; b_sign3 = 4'd9;
@(posedge clk_i);
a_mant0 = 8'd79; a_mant1 = 8'd172; a_mant2 = 8'd151; a_mant3 = 8'd238;
b_mant0 = 8'd29; b_mant1 = 8'd81; b_mant2 = 8'd172; b_mant3 = 8'd141;
a_exp0 = 10'd447; a_exp1 = 10'd638; a_exp2 = 10'd790; a_exp3 = 10'd312;
b_exp0 = 10'd63; b_exp1 = 10'd629; b_exp2 = 10'd464; b_exp3 = 10'd475;
a_sign0 = 4'd7; a_sign1 = 4'd0; a_sign2 = 4'd0; a_sign3 = 4'd1;
b_sign0 = 4'd4; b_sign1 = 4'd5; b_sign2 = 4'd14; b_sign3 = 4'd15;
@(posedge clk_i);
a_mant0 = 8'd16; a_mant1 = 8'd162; a_mant2 = 8'd56; a_mant3 = 8'd33;
b_mant0 = 8'd66; b_mant1 = 8'd41; b_mant2 = 8'd248; b_mant3 = 8'd125;
a_exp0 = 10'd843; a_exp1 = 10'd219; a_exp2 = 10'd549; a_exp3 = 10'd897;
b_exp0 = 10'd905; b_exp1 = 10'd240; b_exp2 = 10'd806; b_exp3 = 10'd230;
a_sign0 = 4'd0; a_sign1 = 4'd13; a_sign2 = 4'd15; a_sign3 = 4'd15;
b_sign0 = 4'd5; b_sign1 = 4'd4; b_sign2 = 4'd4; b_sign3 = 4'd2;
@(posedge clk_i);
a_mant0 = 8'd59; a_mant1 = 8'd241; a_mant2 = 8'd176; a_mant3 = 8'd177;
b_mant0 = 8'd145; b_mant1 = 8'd32; b_mant2 = 8'd127; b_mant3 = 8'd142;
a_exp0 = 10'd394; a_exp1 = 10'd573; a_exp2 = 10'd680; a_exp3 = 10'd395;
b_exp0 = 10'd190; b_exp1 = 10'd832; b_exp2 = 10'd263; b_exp3 = 10'd593;
a_sign0 = 4'd16; a_sign1 = 4'd9; a_sign2 = 4'd10; a_sign3 = 4'd3;
b_sign0 = 4'd10; b_sign1 = 4'd13; b_sign2 = 4'd10; b_sign3 = 4'd13;
@(posedge clk_i);
shared_exps0 = 8'd135;
shared_exps1 = 8'd118;
a_mant0 = 8'd118; a_mant1 = 8'd157; a_mant2 = 8'd16; a_mant3 = 8'd100;
b_mant0 = 8'd207; b_mant1 = 8'd191; b_mant2 = 8'd41; b_mant3 = 8'd215;
a_exp0 = 10'd531; a_exp1 = 10'd619; a_exp2 = 10'd62; a_exp3 = 10'd452;
b_exp0 = 10'd905; b_exp1 = 10'd125; b_exp2 = 10'd933; b_exp3 = 10'd591;
a_sign0 = 4'd6; a_sign1 = 4'd1; a_sign2 = 4'd14; a_sign3 = 4'd10;
b_sign0 = 4'd13; b_sign1 = 4'd16; b_sign2 = 4'd1; b_sign3 = 4'd9;
@(posedge clk_i);
a_mant0 = 8'd183; a_mant1 = 8'd243; a_mant2 = 8'd116; a_mant3 = 8'd200;
b_mant0 = 8'd152; b_mant1 = 8'd65; b_mant2 = 8'd116; b_mant3 = 8'd180;
a_exp0 = 10'd1002; a_exp1 = 10'd355; a_exp2 = 10'd634; a_exp3 = 10'd382;
b_exp0 = 10'd751; b_exp1 = 10'd276; b_exp2 = 10'd319; b_exp3 = 10'd89;
a_sign0 = 4'd7; a_sign1 = 4'd0; a_sign2 = 4'd9; a_sign3 = 4'd3;
b_sign0 = 4'd16; b_sign1 = 4'd8; b_sign2 = 4'd2; b_sign3 = 4'd3;
@(posedge clk_i);
a_mant0 = 8'd134; a_mant1 = 8'd62; a_mant2 = 8'd130; a_mant3 = 8'd155;
b_mant0 = 8'd115; b_mant1 = 8'd58; b_mant2 = 8'd181; b_mant3 = 8'd59;
a_exp0 = 10'd358; a_exp1 = 10'd629; a_exp2 = 10'd250; a_exp3 = 10'd478;
b_exp0 = 10'd961; b_exp1 = 10'd879; b_exp2 = 10'd134; b_exp3 = 10'd929;
a_sign0 = 4'd13; a_sign1 = 4'd14; a_sign2 = 4'd4; a_sign3 = 4'd12;
b_sign0 = 4'd3; b_sign1 = 4'd14; b_sign2 = 4'd12; b_sign3 = 4'd9;
@(posedge clk_i);
a_mant0 = 8'd248; a_mant1 = 8'd158; a_mant2 = 8'd26; a_mant3 = 8'd28;
b_mant0 = 8'd56; b_mant1 = 8'd84; b_mant2 = 8'd57; b_mant3 = 8'd89;
a_exp0 = 10'd989; a_exp1 = 10'd1009; a_exp2 = 10'd415; a_exp3 = 10'd138;
b_exp0 = 10'd776; b_exp1 = 10'd77; b_exp2 = 10'd618; b_exp3 = 10'd328;
a_sign0 = 4'd12; a_sign1 = 4'd8; a_sign2 = 4'd12; a_sign3 = 4'd11;
b_sign0 = 4'd15; b_sign1 = 4'd15; b_sign2 = 4'd6; b_sign3 = 4'd8;
@(posedge clk_i);
a_mant0 = 8'd214; a_mant1 = 8'd226; a_mant2 = 8'd252; a_mant3 = 8'd249;
b_mant0 = 8'd238; b_mant1 = 8'd52; b_mant2 = 8'd176; b_mant3 = 8'd154;
a_exp0 = 10'd218; a_exp1 = 10'd168; a_exp2 = 10'd838; a_exp3 = 10'd785;
b_exp0 = 10'd138; b_exp1 = 10'd334; b_exp2 = 10'd774; b_exp3 = 10'd907;
a_sign0 = 4'd14; a_sign1 = 4'd10; a_sign2 = 4'd6; a_sign3 = 4'd5;
b_sign0 = 4'd5; b_sign1 = 4'd3; b_sign2 = 4'd16; b_sign3 = 4'd13;
@(posedge clk_i);
a_mant0 = 8'd164; a_mant1 = 8'd140; a_mant2 = 8'd22; a_mant3 = 8'd46;
b_mant0 = 8'd97; b_mant1 = 8'd13; b_mant2 = 8'd186; b_mant3 = 8'd182;
a_exp0 = 10'd959; a_exp1 = 10'd560; a_exp2 = 10'd381; a_exp3 = 10'd342;
b_exp0 = 10'd52; b_exp1 = 10'd473; b_exp2 = 10'd876; b_exp3 = 10'd797;
a_sign0 = 4'd16; a_sign1 = 4'd12; a_sign2 = 4'd4; a_sign3 = 4'd1;
b_sign0 = 4'd3; b_sign1 = 4'd16; b_sign2 = 4'd14; b_sign3 = 4'd4;
@(posedge clk_i);
a_mant0 = 8'd211; a_mant1 = 8'd104; a_mant2 = 8'd79; a_mant3 = 8'd226;
b_mant0 = 8'd12; b_mant1 = 8'd210; b_mant2 = 8'd6; b_mant3 = 8'd16;
a_exp0 = 10'd985; a_exp1 = 10'd706; a_exp2 = 10'd834; a_exp3 = 10'd9;
b_exp0 = 10'd839; b_exp1 = 10'd982; b_exp2 = 10'd746; b_exp3 = 10'd252;
a_sign0 = 4'd4; a_sign1 = 4'd10; a_sign2 = 4'd4; a_sign3 = 4'd4;
b_sign0 = 4'd3; b_sign1 = 4'd4; b_sign2 = 4'd15; b_sign3 = 4'd2;
@(posedge clk_i);
a_mant0 = 8'd231; a_mant1 = 8'd93; a_mant2 = 8'd226; a_mant3 = 8'd172;
b_mant0 = 8'd15; b_mant1 = 8'd12; b_mant2 = 8'd113; b_mant3 = 8'd21;
a_exp0 = 10'd434; a_exp1 = 10'd941; a_exp2 = 10'd792; a_exp3 = 10'd739;
b_exp0 = 10'd414; b_exp1 = 10'd295; b_exp2 = 10'd399; b_exp3 = 10'd491;
a_sign0 = 4'd1; a_sign1 = 4'd5; a_sign2 = 4'd12; a_sign3 = 4'd8;
b_sign0 = 4'd0; b_sign1 = 4'd5; b_sign2 = 4'd6; b_sign3 = 4'd16;
@(posedge clk_i);
shared_exps0 = 8'd124;
shared_exps1 = 8'd118;
a_mant0 = 8'd42; a_mant1 = 8'd92; a_mant2 = 8'd177; a_mant3 = 8'd83;
b_mant0 = 8'd98; b_mant1 = 8'd212; b_mant2 = 8'd165; b_mant3 = 8'd194;
a_exp0 = 10'd61; a_exp1 = 10'd327; a_exp2 = 10'd757; a_exp3 = 10'd515;
b_exp0 = 10'd778; b_exp1 = 10'd585; b_exp2 = 10'd445; b_exp3 = 10'd442;
a_sign0 = 4'd16; a_sign1 = 4'd6; a_sign2 = 4'd7; a_sign3 = 4'd9;
b_sign0 = 4'd14; b_sign1 = 4'd1; b_sign2 = 4'd10; b_sign3 = 4'd14;
@(posedge clk_i);
a_mant0 = 8'd158; a_mant1 = 8'd18; a_mant2 = 8'd35; a_mant3 = 8'd241;
b_mant0 = 8'd120; b_mant1 = 8'd174; b_mant2 = 8'd120; b_mant3 = 8'd107;
a_exp0 = 10'd640; a_exp1 = 10'd12; a_exp2 = 10'd214; a_exp3 = 10'd538;
b_exp0 = 10'd64; b_exp1 = 10'd391; b_exp2 = 10'd198; b_exp3 = 10'd306;
a_sign0 = 4'd14; a_sign1 = 4'd16; a_sign2 = 4'd0; a_sign3 = 4'd9;
b_sign0 = 4'd9; b_sign1 = 4'd7; b_sign2 = 4'd8; b_sign3 = 4'd1;
@(posedge clk_i);
a_mant0 = 8'd2; a_mant1 = 8'd143; a_mant2 = 8'd152; a_mant3 = 8'd151;
b_mant0 = 8'd27; b_mant1 = 8'd166; b_mant2 = 8'd188; b_mant3 = 8'd150;
a_exp0 = 10'd330; a_exp1 = 10'd621; a_exp2 = 10'd374; a_exp3 = 10'd460;
b_exp0 = 10'd198; b_exp1 = 10'd39; b_exp2 = 10'd112; b_exp3 = 10'd805;
a_sign0 = 4'd3; a_sign1 = 4'd1; a_sign2 = 4'd16; a_sign3 = 4'd2;
b_sign0 = 4'd14; b_sign1 = 4'd16; b_sign2 = 4'd2; b_sign3 = 4'd1;
@(posedge clk_i);
a_mant0 = 8'd182; a_mant1 = 8'd102; a_mant2 = 8'd173; a_mant3 = 8'd97;
b_mant0 = 8'd154; b_mant1 = 8'd140; b_mant2 = 8'd59; b_mant3 = 8'd68;
a_exp0 = 10'd394; a_exp1 = 10'd863; a_exp2 = 10'd600; a_exp3 = 10'd74;
b_exp0 = 10'd654; b_exp1 = 10'd525; b_exp2 = 10'd670; b_exp3 = 10'd299;
a_sign0 = 4'd4; a_sign1 = 4'd9; a_sign2 = 4'd15; a_sign3 = 4'd7;
b_sign0 = 4'd2; b_sign1 = 4'd1; b_sign2 = 4'd16; b_sign3 = 4'd7;
@(posedge clk_i);
a_mant0 = 8'd206; a_mant1 = 8'd176; a_mant2 = 8'd220; a_mant3 = 8'd86;
b_mant0 = 8'd2; b_mant1 = 8'd177; b_mant2 = 8'd98; b_mant3 = 8'd60;
a_exp0 = 10'd916; a_exp1 = 10'd795; a_exp2 = 10'd674; a_exp3 = 10'd960;
b_exp0 = 10'd398; b_exp1 = 10'd375; b_exp2 = 10'd383; b_exp3 = 10'd139;
a_sign0 = 4'd15; a_sign1 = 4'd7; a_sign2 = 4'd12; a_sign3 = 4'd5;
b_sign0 = 4'd6; b_sign1 = 4'd16; b_sign2 = 4'd6; b_sign3 = 4'd10;
@(posedge clk_i);
a_mant0 = 8'd248; a_mant1 = 8'd86; a_mant2 = 8'd178; a_mant3 = 8'd101;
b_mant0 = 8'd38; b_mant1 = 8'd48; b_mant2 = 8'd30; b_mant3 = 8'd180;
a_exp0 = 10'd657; a_exp1 = 10'd600; a_exp2 = 10'd488; a_exp3 = 10'd257;
b_exp0 = 10'd146; b_exp1 = 10'd760; b_exp2 = 10'd785; b_exp3 = 10'd581;
a_sign0 = 4'd5; a_sign1 = 4'd14; a_sign2 = 4'd2; a_sign3 = 4'd14;
b_sign0 = 4'd5; b_sign1 = 4'd2; b_sign2 = 4'd13; b_sign3 = 4'd4;
@(posedge clk_i);
a_mant0 = 8'd232; a_mant1 = 8'd173; a_mant2 = 8'd7; a_mant3 = 8'd18;
b_mant0 = 8'd219; b_mant1 = 8'd7; b_mant2 = 8'd156; b_mant3 = 8'd77;
a_exp0 = 10'd179; a_exp1 = 10'd271; a_exp2 = 10'd354; a_exp3 = 10'd417;
b_exp0 = 10'd805; b_exp1 = 10'd72; b_exp2 = 10'd568; b_exp3 = 10'd872;
a_sign0 = 4'd10; a_sign1 = 4'd15; a_sign2 = 4'd7; a_sign3 = 4'd10;
b_sign0 = 4'd5; b_sign1 = 4'd1; b_sign2 = 4'd6; b_sign3 = 4'd4;
@(posedge clk_i);
a_mant0 = 8'd6; a_mant1 = 8'd140; a_mant2 = 8'd52; a_mant3 = 8'd60;
b_mant0 = 8'd85; b_mant1 = 8'd235; b_mant2 = 8'd129; b_mant3 = 8'd251;
a_exp0 = 10'd16; a_exp1 = 10'd671; a_exp2 = 10'd362; a_exp3 = 10'd187;
b_exp0 = 10'd13; b_exp1 = 10'd31; b_exp2 = 10'd684; b_exp3 = 10'd87;
a_sign0 = 4'd12; a_sign1 = 4'd6; a_sign2 = 4'd12; a_sign3 = 4'd7;
b_sign0 = 4'd0; b_sign1 = 4'd13; b_sign2 = 4'd1; b_sign3 = 4'd2;
@(posedge clk_i);
shared_exps0 = 8'd137;
shared_exps1 = 8'd111;
a_mant0 = 8'd184; a_mant1 = 8'd94; a_mant2 = 8'd102; a_mant3 = 8'd0;
b_mant0 = 8'd87; b_mant1 = 8'd175; b_mant2 = 8'd73; b_mant3 = 8'd99;
a_exp0 = 10'd225; a_exp1 = 10'd367; a_exp2 = 10'd806; a_exp3 = 10'd702;
b_exp0 = 10'd88; b_exp1 = 10'd669; b_exp2 = 10'd26; b_exp3 = 10'd797;
a_sign0 = 4'd13; a_sign1 = 4'd7; a_sign2 = 4'd15; a_sign3 = 4'd3;
b_sign0 = 4'd6; b_sign1 = 4'd12; b_sign2 = 4'd14; b_sign3 = 4'd7;
@(posedge clk_i);
a_mant0 = 8'd11; a_mant1 = 8'd81; a_mant2 = 8'd137; a_mant3 = 8'd161;
b_mant0 = 8'd196; b_mant1 = 8'd247; b_mant2 = 8'd169; b_mant3 = 8'd158;
a_exp0 = 10'd591; a_exp1 = 10'd81; a_exp2 = 10'd98; a_exp3 = 10'd592;
b_exp0 = 10'd343; b_exp1 = 10'd620; b_exp2 = 10'd712; b_exp3 = 10'd373;
a_sign0 = 4'd6; a_sign1 = 4'd8; a_sign2 = 4'd16; a_sign3 = 4'd9;
b_sign0 = 4'd15; b_sign1 = 4'd1; b_sign2 = 4'd15; b_sign3 = 4'd1;
@(posedge clk_i);
a_mant0 = 8'd112; a_mant1 = 8'd227; a_mant2 = 8'd31; a_mant3 = 8'd203;
b_mant0 = 8'd255; b_mant1 = 8'd119; b_mant2 = 8'd130; b_mant3 = 8'd164;
a_exp0 = 10'd365; a_exp1 = 10'd256; a_exp2 = 10'd266; a_exp3 = 10'd163;
b_exp0 = 10'd244; b_exp1 = 10'd754; b_exp2 = 10'd333; b_exp3 = 10'd65;
a_sign0 = 4'd12; a_sign1 = 4'd5; a_sign2 = 4'd6; a_sign3 = 4'd16;
b_sign0 = 4'd8; b_sign1 = 4'd2; b_sign2 = 4'd0; b_sign3 = 4'd3;
@(posedge clk_i);
a_mant0 = 8'd46; a_mant1 = 8'd49; a_mant2 = 8'd164; a_mant3 = 8'd210;
b_mant0 = 8'd112; b_mant1 = 8'd154; b_mant2 = 8'd30; b_mant3 = 8'd19;
a_exp0 = 10'd215; a_exp1 = 10'd62; a_exp2 = 10'd254; a_exp3 = 10'd350;
b_exp0 = 10'd464; b_exp1 = 10'd651; b_exp2 = 10'd873; b_exp3 = 10'd620;
a_sign0 = 4'd8; a_sign1 = 4'd15; a_sign2 = 4'd11; a_sign3 = 4'd9;
b_sign0 = 4'd15; b_sign1 = 4'd10; b_sign2 = 4'd6; b_sign3 = 4'd0;
@(posedge clk_i);
a_mant0 = 8'd153; a_mant1 = 8'd103; a_mant2 = 8'd204; a_mant3 = 8'd98;
b_mant0 = 8'd227; b_mant1 = 8'd191; b_mant2 = 8'd24; b_mant3 = 8'd153;
a_exp0 = 10'd516; a_exp1 = 10'd686; a_exp2 = 10'd530; a_exp3 = 10'd666;
b_exp0 = 10'd358; b_exp1 = 10'd888; b_exp2 = 10'd564; b_exp3 = 10'd465;
a_sign0 = 4'd14; a_sign1 = 4'd0; a_sign2 = 4'd16; a_sign3 = 4'd6;
b_sign0 = 4'd11; b_sign1 = 4'd3; b_sign2 = 4'd14; b_sign3 = 4'd14;
@(posedge clk_i);
a_mant0 = 8'd249; a_mant1 = 8'd101; a_mant2 = 8'd186; a_mant3 = 8'd79;
b_mant0 = 8'd28; b_mant1 = 8'd39; b_mant2 = 8'd197; b_mant3 = 8'd109;
a_exp0 = 10'd193; a_exp1 = 10'd52; a_exp2 = 10'd1015; a_exp3 = 10'd229;
b_exp0 = 10'd422; b_exp1 = 10'd77; b_exp2 = 10'd329; b_exp3 = 10'd238;
a_sign0 = 4'd2; a_sign1 = 4'd9; a_sign2 = 4'd10; a_sign3 = 4'd1;
b_sign0 = 4'd12; b_sign1 = 4'd6; b_sign2 = 4'd6; b_sign3 = 4'd7;
@(posedge clk_i);
a_mant0 = 8'd199; a_mant1 = 8'd52; a_mant2 = 8'd235; a_mant3 = 8'd81;
b_mant0 = 8'd9; b_mant1 = 8'd216; b_mant2 = 8'd51; b_mant3 = 8'd64;
a_exp0 = 10'd613; a_exp1 = 10'd84; a_exp2 = 10'd30; a_exp3 = 10'd797;
b_exp0 = 10'd361; b_exp1 = 10'd964; b_exp2 = 10'd837; b_exp3 = 10'd918;
a_sign0 = 4'd4; a_sign1 = 4'd8; a_sign2 = 4'd7; a_sign3 = 4'd1;
b_sign0 = 4'd16; b_sign1 = 4'd7; b_sign2 = 4'd7; b_sign3 = 4'd4;
@(posedge clk_i);
a_mant0 = 8'd242; a_mant1 = 8'd34; a_mant2 = 8'd116; a_mant3 = 8'd209;
b_mant0 = 8'd65; b_mant1 = 8'd254; b_mant2 = 8'd37; b_mant3 = 8'd155;
a_exp0 = 10'd409; a_exp1 = 10'd663; a_exp2 = 10'd823; a_exp3 = 10'd891;
b_exp0 = 10'd142; b_exp1 = 10'd949; b_exp2 = 10'd915; b_exp3 = 10'd715;
a_sign0 = 4'd4; a_sign1 = 4'd10; a_sign2 = 4'd9; a_sign3 = 4'd1;
b_sign0 = 4'd5; b_sign1 = 4'd14; b_sign2 = 4'd0; b_sign3 = 4'd5;
@(posedge clk_i);
shared_exps0 = 8'd138;
shared_exps1 = 8'd99;
rstn = 0;
@(posedge clk_i);
rstn = 1;
a_mant0 = 8'd47; a_mant1 = 8'd215; a_mant2 = 8'd16; a_mant3 = 8'd89;
b_mant0 = 8'd65; b_mant1 = 8'd70; b_mant2 = 8'd30; b_mant3 = 8'd93;
a_exp0 = 10'd280; a_exp1 = 10'd1001; a_exp2 = 10'd4; a_exp3 = 10'd898;
b_exp0 = 10'd842; b_exp1 = 10'd142; b_exp2 = 10'd749; b_exp3 = 10'd542;
a_sign0 = 4'd9; a_sign1 = 4'd10; a_sign2 = 4'd14; a_sign3 = 4'd3;
b_sign0 = 4'd13; b_sign1 = 4'd6; b_sign2 = 4'd5; b_sign3 = 4'd16;
@(posedge clk_i);
a_mant0 = 8'd7; a_mant1 = 8'd178; a_mant2 = 8'd184; a_mant3 = 8'd30;
b_mant0 = 8'd29; b_mant1 = 8'd193; b_mant2 = 8'd130; b_mant3 = 8'd133;
a_exp0 = 10'd231; a_exp1 = 10'd357; a_exp2 = 10'd983; a_exp3 = 10'd262;
b_exp0 = 10'd135; b_exp1 = 10'd367; b_exp2 = 10'd99; b_exp3 = 10'd973;
a_sign0 = 4'd6; a_sign1 = 4'd5; a_sign2 = 4'd4; a_sign3 = 4'd3;
b_sign0 = 4'd1; b_sign1 = 4'd6; b_sign2 = 4'd12; b_sign3 = 4'd13;
@(posedge clk_i);
a_mant0 = 8'd227; a_mant1 = 8'd64; a_mant2 = 8'd248; a_mant3 = 8'd95;
b_mant0 = 8'd153; b_mant1 = 8'd195; b_mant2 = 8'd28; b_mant3 = 8'd139;
a_exp0 = 10'd798; a_exp1 = 10'd145; a_exp2 = 10'd451; a_exp3 = 10'd565;
b_exp0 = 10'd102; b_exp1 = 10'd196; b_exp2 = 10'd440; b_exp3 = 10'd991;
a_sign0 = 4'd5; a_sign1 = 4'd10; a_sign2 = 4'd2; a_sign3 = 4'd1;
b_sign0 = 4'd6; b_sign1 = 4'd16; b_sign2 = 4'd14; b_sign3 = 4'd15;
@(posedge clk_i);
a_mant0 = 8'd219; a_mant1 = 8'd145; a_mant2 = 8'd102; a_mant3 = 8'd203;
b_mant0 = 8'd191; b_mant1 = 8'd97; b_mant2 = 8'd253; b_mant3 = 8'd127;
a_exp0 = 10'd707; a_exp1 = 10'd654; a_exp2 = 10'd549; a_exp3 = 10'd596;
b_exp0 = 10'd922; b_exp1 = 10'd349; b_exp2 = 10'd257; b_exp3 = 10'd332;
a_sign0 = 4'd11; a_sign1 = 4'd3; a_sign2 = 4'd8; a_sign3 = 4'd16;
b_sign0 = 4'd16; b_sign1 = 4'd7; b_sign2 = 4'd2; b_sign3 = 4'd2;
@(posedge clk_i);
a_mant0 = 8'd238; a_mant1 = 8'd8; a_mant2 = 8'd180; a_mant3 = 8'd182;
b_mant0 = 8'd240; b_mant1 = 8'd220; b_mant2 = 8'd47; b_mant3 = 8'd19;
a_exp0 = 10'd454; a_exp1 = 10'd823; a_exp2 = 10'd200; a_exp3 = 10'd54;
b_exp0 = 10'd1011; b_exp1 = 10'd211; b_exp2 = 10'd982; b_exp3 = 10'd259;
a_sign0 = 4'd12; a_sign1 = 4'd0; a_sign2 = 4'd11; a_sign3 = 4'd0;
b_sign0 = 4'd14; b_sign1 = 4'd6; b_sign2 = 4'd4; b_sign3 = 4'd14;
@(posedge clk_i);
a_mant0 = 8'd75; a_mant1 = 8'd188; a_mant2 = 8'd207; a_mant3 = 8'd15;
b_mant0 = 8'd172; b_mant1 = 8'd154; b_mant2 = 8'd203; b_mant3 = 8'd60;
a_exp0 = 10'd781; a_exp1 = 10'd998; a_exp2 = 10'd728; a_exp3 = 10'd114;
b_exp0 = 10'd933; b_exp1 = 10'd1004; b_exp2 = 10'd251; b_exp3 = 10'd813;
a_sign0 = 4'd6; a_sign1 = 4'd3; a_sign2 = 4'd5; a_sign3 = 4'd9;
b_sign0 = 4'd13; b_sign1 = 4'd9; b_sign2 = 4'd15; b_sign3 = 4'd3;
@(posedge clk_i);
a_mant0 = 8'd112; a_mant1 = 8'd21; a_mant2 = 8'd219; a_mant3 = 8'd28;
b_mant0 = 8'd52; b_mant1 = 8'd137; b_mant2 = 8'd202; b_mant3 = 8'd170;
a_exp0 = 10'd579; a_exp1 = 10'd670; a_exp2 = 10'd281; a_exp3 = 10'd13;
b_exp0 = 10'd68; b_exp1 = 10'd832; b_exp2 = 10'd898; b_exp3 = 10'd126;
a_sign0 = 4'd11; a_sign1 = 4'd11; a_sign2 = 4'd11; a_sign3 = 4'd3;
b_sign0 = 4'd2; b_sign1 = 4'd4; b_sign2 = 4'd11; b_sign3 = 4'd11;
@(posedge clk_i);
shared_exps0 = 8'd112;
shared_exps1 = 8'd128;
a_mant0 = 8'd101; a_mant1 = 8'd240; a_mant2 = 8'd205; a_mant3 = 8'd129;
b_mant0 = 8'd205; b_mant1 = 8'd67; b_mant2 = 8'd75; b_mant3 = 8'd81;
a_exp0 = 10'd1017; a_exp1 = 10'd194; a_exp2 = 10'd315; a_exp3 = 10'd611;
b_exp0 = 10'd940; b_exp1 = 10'd412; b_exp2 = 10'd767; b_exp3 = 10'd870;
a_sign0 = 4'd9; a_sign1 = 4'd2; a_sign2 = 4'd9; a_sign3 = 4'd2;
b_sign0 = 4'd10; b_sign1 = 4'd8; b_sign2 = 4'd15; b_sign3 = 4'd11;
@(posedge clk_i);
a_mant0 = 8'd145; a_mant1 = 8'd188; a_mant2 = 8'd174; a_mant3 = 8'd218;
b_mant0 = 8'd109; b_mant1 = 8'd119; b_mant2 = 8'd112; b_mant3 = 8'd65;
a_exp0 = 10'd887; a_exp1 = 10'd143; a_exp2 = 10'd935; a_exp3 = 10'd638;
b_exp0 = 10'd604; b_exp1 = 10'd254; b_exp2 = 10'd670; b_exp3 = 10'd410;
a_sign0 = 4'd6; a_sign1 = 4'd15; a_sign2 = 4'd11; a_sign3 = 4'd0;
b_sign0 = 4'd0; b_sign1 = 4'd0; b_sign2 = 4'd11; b_sign3 = 4'd7;
@(posedge clk_i);
a_mant0 = 8'd163; a_mant1 = 8'd160; a_mant2 = 8'd200; a_mant3 = 8'd208;
b_mant0 = 8'd10; b_mant1 = 8'd111; b_mant2 = 8'd220; b_mant3 = 8'd172;
a_exp0 = 10'd177; a_exp1 = 10'd826; a_exp2 = 10'd776; a_exp3 = 10'd625;
b_exp0 = 10'd851; b_exp1 = 10'd235; b_exp2 = 10'd636; b_exp3 = 10'd934;
a_sign0 = 4'd13; a_sign1 = 4'd11; a_sign2 = 4'd5; a_sign3 = 4'd13;
b_sign0 = 4'd0; b_sign1 = 4'd7; b_sign2 = 4'd8; b_sign3 = 4'd0;
@(posedge clk_i);
a_mant0 = 8'd238; a_mant1 = 8'd147; a_mant2 = 8'd40; a_mant3 = 8'd190;
b_mant0 = 8'd40; b_mant1 = 8'd167; b_mant2 = 8'd209; b_mant3 = 8'd95;
a_exp0 = 10'd956; a_exp1 = 10'd917; a_exp2 = 10'd636; a_exp3 = 10'd736;
b_exp0 = 10'd448; b_exp1 = 10'd888; b_exp2 = 10'd978; b_exp3 = 10'd718;
a_sign0 = 4'd14; a_sign1 = 4'd2; a_sign2 = 4'd9; a_sign3 = 4'd2;
b_sign0 = 4'd0; b_sign1 = 4'd12; b_sign2 = 4'd15; b_sign3 = 4'd13;
@(posedge clk_i);
a_mant0 = 8'd61; a_mant1 = 8'd60; a_mant2 = 8'd158; a_mant3 = 8'd14;
b_mant0 = 8'd155; b_mant1 = 8'd190; b_mant2 = 8'd46; b_mant3 = 8'd242;
a_exp0 = 10'd903; a_exp1 = 10'd504; a_exp2 = 10'd64; a_exp3 = 10'd221;
b_exp0 = 10'd738; b_exp1 = 10'd965; b_exp2 = 10'd393; b_exp3 = 10'd821;
a_sign0 = 4'd7; a_sign1 = 4'd12; a_sign2 = 4'd7; a_sign3 = 4'd15;
b_sign0 = 4'd11; b_sign1 = 4'd10; b_sign2 = 4'd14; b_sign3 = 4'd0;
@(posedge clk_i);
a_mant0 = 8'd201; a_mant1 = 8'd243; a_mant2 = 8'd174; a_mant3 = 8'd239;
b_mant0 = 8'd175; b_mant1 = 8'd85; b_mant2 = 8'd11; b_mant3 = 8'd121;
a_exp0 = 10'd616; a_exp1 = 10'd987; a_exp2 = 10'd262; a_exp3 = 10'd850;
b_exp0 = 10'd850; b_exp1 = 10'd587; b_exp2 = 10'd488; b_exp3 = 10'd947;
a_sign0 = 4'd15; a_sign1 = 4'd2; a_sign2 = 4'd14; a_sign3 = 4'd4;
b_sign0 = 4'd1; b_sign1 = 4'd9; b_sign2 = 4'd16; b_sign3 = 4'd8;
@(posedge clk_i);
a_mant0 = 8'd57; a_mant1 = 8'd243; a_mant2 = 8'd87; a_mant3 = 8'd167;
b_mant0 = 8'd128; b_mant1 = 8'd133; b_mant2 = 8'd254; b_mant3 = 8'd70;
a_exp0 = 10'd897; a_exp1 = 10'd193; a_exp2 = 10'd279; a_exp3 = 10'd71;
b_exp0 = 10'd380; b_exp1 = 10'd467; b_exp2 = 10'd755; b_exp3 = 10'd925;
a_sign0 = 4'd10; a_sign1 = 4'd16; a_sign2 = 4'd13; a_sign3 = 4'd0;
b_sign0 = 4'd14; b_sign1 = 4'd12; b_sign2 = 4'd13; b_sign3 = 4'd16;
@(posedge clk_i);
a_mant0 = 8'd65; a_mant1 = 8'd167; a_mant2 = 8'd72; a_mant3 = 8'd253;
b_mant0 = 8'd100; b_mant1 = 8'd66; b_mant2 = 8'd189; b_mant3 = 8'd111;
a_exp0 = 10'd914; a_exp1 = 10'd803; a_exp2 = 10'd1023; a_exp3 = 10'd550;
b_exp0 = 10'd168; b_exp1 = 10'd835; b_exp2 = 10'd635; b_exp3 = 10'd207;
a_sign0 = 4'd2; a_sign1 = 4'd4; a_sign2 = 4'd8; a_sign3 = 4'd1;
b_sign0 = 4'd12; b_sign1 = 4'd2; b_sign2 = 4'd0; b_sign3 = 4'd5;
@(posedge clk_i);
shared_exps0 = 8'd122;
shared_exps1 = 8'd144;
a_mant0 = 8'd82; a_mant1 = 8'd97; a_mant2 = 8'd174; a_mant3 = 8'd242;
b_mant0 = 8'd218; b_mant1 = 8'd188; b_mant2 = 8'd87; b_mant3 = 8'd94;
a_exp0 = 10'd332; a_exp1 = 10'd766; a_exp2 = 10'd536; a_exp3 = 10'd257;
b_exp0 = 10'd544; b_exp1 = 10'd474; b_exp2 = 10'd632; b_exp3 = 10'd143;
a_sign0 = 4'd8; a_sign1 = 4'd11; a_sign2 = 4'd4; a_sign3 = 4'd4;
b_sign0 = 4'd2; b_sign1 = 4'd6; b_sign2 = 4'd4; b_sign3 = 4'd11;
@(posedge clk_i);
a_mant0 = 8'd28; a_mant1 = 8'd163; a_mant2 = 8'd125; a_mant3 = 8'd100;
b_mant0 = 8'd204; b_mant1 = 8'd219; b_mant2 = 8'd6; b_mant3 = 8'd118;
a_exp0 = 10'd792; a_exp1 = 10'd690; a_exp2 = 10'd888; a_exp3 = 10'd325;
b_exp0 = 10'd384; b_exp1 = 10'd757; b_exp2 = 10'd225; b_exp3 = 10'd307;
a_sign0 = 4'd7; a_sign1 = 4'd9; a_sign2 = 4'd11; a_sign3 = 4'd12;
b_sign0 = 4'd16; b_sign1 = 4'd15; b_sign2 = 4'd8; b_sign3 = 4'd5;
@(posedge clk_i);
a_mant0 = 8'd89; a_mant1 = 8'd182; a_mant2 = 8'd93; a_mant3 = 8'd188;
b_mant0 = 8'd128; b_mant1 = 8'd90; b_mant2 = 8'd220; b_mant3 = 8'd95;
a_exp0 = 10'd587; a_exp1 = 10'd291; a_exp2 = 10'd539; a_exp3 = 10'd842;
b_exp0 = 10'd40; b_exp1 = 10'd972; b_exp2 = 10'd376; b_exp3 = 10'd777;
a_sign0 = 4'd4; a_sign1 = 4'd8; a_sign2 = 4'd12; a_sign3 = 4'd12;
b_sign0 = 4'd12; b_sign1 = 4'd3; b_sign2 = 4'd7; b_sign3 = 4'd12;
@(posedge clk_i);
a_mant0 = 8'd90; a_mant1 = 8'd225; a_mant2 = 8'd244; a_mant3 = 8'd3;
b_mant0 = 8'd170; b_mant1 = 8'd4; b_mant2 = 8'd104; b_mant3 = 8'd12;
a_exp0 = 10'd453; a_exp1 = 10'd840; a_exp2 = 10'd339; a_exp3 = 10'd474;
b_exp0 = 10'd954; b_exp1 = 10'd207; b_exp2 = 10'd100; b_exp3 = 10'd348;
a_sign0 = 4'd3; a_sign1 = 4'd14; a_sign2 = 4'd13; a_sign3 = 4'd1;
b_sign0 = 4'd7; b_sign1 = 4'd16; b_sign2 = 4'd4; b_sign3 = 4'd0;
@(posedge clk_i);
a_mant0 = 8'd255; a_mant1 = 8'd0; a_mant2 = 8'd235; a_mant3 = 8'd188;
b_mant0 = 8'd181; b_mant1 = 8'd100; b_mant2 = 8'd76; b_mant3 = 8'd7;
a_exp0 = 10'd777; a_exp1 = 10'd439; a_exp2 = 10'd779; a_exp3 = 10'd684;
b_exp0 = 10'd143; b_exp1 = 10'd425; b_exp2 = 10'd249; b_exp3 = 10'd684;
a_sign0 = 4'd5; a_sign1 = 4'd6; a_sign2 = 4'd9; a_sign3 = 4'd7;
b_sign0 = 4'd15; b_sign1 = 4'd8; b_sign2 = 4'd14; b_sign3 = 4'd13;
@(posedge clk_i);
a_mant0 = 8'd241; a_mant1 = 8'd193; a_mant2 = 8'd14; a_mant3 = 8'd241;
b_mant0 = 8'd97; b_mant1 = 8'd199; b_mant2 = 8'd139; b_mant3 = 8'd231;
a_exp0 = 10'd1011; a_exp1 = 10'd630; a_exp2 = 10'd154; a_exp3 = 10'd141;
b_exp0 = 10'd804; b_exp1 = 10'd149; b_exp2 = 10'd76; b_exp3 = 10'd688;
a_sign0 = 4'd9; a_sign1 = 4'd5; a_sign2 = 4'd2; a_sign3 = 4'd16;
b_sign0 = 4'd8; b_sign1 = 4'd14; b_sign2 = 4'd5; b_sign3 = 4'd1;
@(posedge clk_i);
a_mant0 = 8'd98; a_mant1 = 8'd119; a_mant2 = 8'd180; a_mant3 = 8'd250;
b_mant0 = 8'd29; b_mant1 = 8'd180; b_mant2 = 8'd197; b_mant3 = 8'd108;
a_exp0 = 10'd836; a_exp1 = 10'd50; a_exp2 = 10'd863; a_exp3 = 10'd755;
b_exp0 = 10'd460; b_exp1 = 10'd357; b_exp2 = 10'd273; b_exp3 = 10'd955;
a_sign0 = 4'd11; a_sign1 = 4'd3; a_sign2 = 4'd4; a_sign3 = 4'd12;
b_sign0 = 4'd5; b_sign1 = 4'd13; b_sign2 = 4'd15; b_sign3 = 4'd5;
@(posedge clk_i);
a_mant0 = 8'd243; a_mant1 = 8'd145; a_mant2 = 8'd248; a_mant3 = 8'd87;
b_mant0 = 8'd138; b_mant1 = 8'd134; b_mant2 = 8'd221; b_mant3 = 8'd62;
a_exp0 = 10'd928; a_exp1 = 10'd493; a_exp2 = 10'd343; a_exp3 = 10'd262;
b_exp0 = 10'd19; b_exp1 = 10'd648; b_exp2 = 10'd760; b_exp3 = 10'd10;
a_sign0 = 4'd14; a_sign1 = 4'd12; a_sign2 = 4'd2; a_sign3 = 4'd15;
b_sign0 = 4'd16; b_sign1 = 4'd15; b_sign2 = 4'd6; b_sign3 = 4'd9;
@(posedge clk_i);
shared_exps0 = 8'd136;
shared_exps1 = 8'd156;
a_mant0 = 8'd35; a_mant1 = 8'd28; a_mant2 = 8'd15; a_mant3 = 8'd30;
b_mant0 = 8'd25; b_mant1 = 8'd14; b_mant2 = 8'd15; b_mant3 = 8'd152;
a_exp0 = 10'd810; a_exp1 = 10'd188; a_exp2 = 10'd57; a_exp3 = 10'd632;
b_exp0 = 10'd538; b_exp1 = 10'd226; b_exp2 = 10'd243; b_exp3 = 10'd960;
a_sign0 = 4'd10; a_sign1 = 4'd16; a_sign2 = 4'd1; a_sign3 = 4'd8;
b_sign0 = 4'd6; b_sign1 = 4'd16; b_sign2 = 4'd10; b_sign3 = 4'd1;
@(posedge clk_i);
a_mant0 = 8'd50; a_mant1 = 8'd197; a_mant2 = 8'd218; a_mant3 = 8'd203;
b_mant0 = 8'd27; b_mant1 = 8'd36; b_mant2 = 8'd105; b_mant3 = 8'd118;
a_exp0 = 10'd954; a_exp1 = 10'd378; a_exp2 = 10'd933; a_exp3 = 10'd586;
b_exp0 = 10'd325; b_exp1 = 10'd128; b_exp2 = 10'd552; b_exp3 = 10'd811;
a_sign0 = 4'd5; a_sign1 = 4'd3; a_sign2 = 4'd11; a_sign3 = 4'd4;
b_sign0 = 4'd12; b_sign1 = 4'd5; b_sign2 = 4'd6; b_sign3 = 4'd13;
@(posedge clk_i);
a_mant0 = 8'd49; a_mant1 = 8'd27; a_mant2 = 8'd95; a_mant3 = 8'd91;
b_mant0 = 8'd179; b_mant1 = 8'd199; b_mant2 = 8'd65; b_mant3 = 8'd95;
a_exp0 = 10'd230; a_exp1 = 10'd257; a_exp2 = 10'd783; a_exp3 = 10'd304;
b_exp0 = 10'd640; b_exp1 = 10'd175; b_exp2 = 10'd712; b_exp3 = 10'd784;
a_sign0 = 4'd5; a_sign1 = 4'd10; a_sign2 = 4'd7; a_sign3 = 4'd1;
b_sign0 = 4'd4; b_sign1 = 4'd8; b_sign2 = 4'd13; b_sign3 = 4'd10;
@(posedge clk_i);
a_mant0 = 8'd81; a_mant1 = 8'd67; a_mant2 = 8'd24; a_mant3 = 8'd34;
b_mant0 = 8'd201; b_mant1 = 8'd144; b_mant2 = 8'd134; b_mant3 = 8'd188;
a_exp0 = 10'd99; a_exp1 = 10'd955; a_exp2 = 10'd391; a_exp3 = 10'd76;
b_exp0 = 10'd979; b_exp1 = 10'd70; b_exp2 = 10'd756; b_exp3 = 10'd222;
a_sign0 = 4'd4; a_sign1 = 4'd14; a_sign2 = 4'd7; a_sign3 = 4'd11;
b_sign0 = 4'd2; b_sign1 = 4'd15; b_sign2 = 4'd10; b_sign3 = 4'd10;
@(posedge clk_i);
a_mant0 = 8'd127; a_mant1 = 8'd175; a_mant2 = 8'd64; a_mant3 = 8'd111;
b_mant0 = 8'd35; b_mant1 = 8'd77; b_mant2 = 8'd255; b_mant3 = 8'd74;
a_exp0 = 10'd663; a_exp1 = 10'd180; a_exp2 = 10'd433; a_exp3 = 10'd690;
b_exp0 = 10'd2; b_exp1 = 10'd276; b_exp2 = 10'd370; b_exp3 = 10'd908;
a_sign0 = 4'd15; a_sign1 = 4'd9; a_sign2 = 4'd6; a_sign3 = 4'd9;
b_sign0 = 4'd13; b_sign1 = 4'd0; b_sign2 = 4'd4; b_sign3 = 4'd12;
@(posedge clk_i);
a_mant0 = 8'd173; a_mant1 = 8'd42; a_mant2 = 8'd225; a_mant3 = 8'd208;
b_mant0 = 8'd139; b_mant1 = 8'd214; b_mant2 = 8'd169; b_mant3 = 8'd92;
a_exp0 = 10'd838; a_exp1 = 10'd880; a_exp2 = 10'd900; a_exp3 = 10'd228;
b_exp0 = 10'd542; b_exp1 = 10'd110; b_exp2 = 10'd568; b_exp3 = 10'd914;
a_sign0 = 4'd1; a_sign1 = 4'd13; a_sign2 = 4'd10; a_sign3 = 4'd0;
b_sign0 = 4'd12; b_sign1 = 4'd5; b_sign2 = 4'd10; b_sign3 = 4'd7;
@(posedge clk_i);
a_mant0 = 8'd54; a_mant1 = 8'd182; a_mant2 = 8'd106; a_mant3 = 8'd199;
b_mant0 = 8'd46; b_mant1 = 8'd87; b_mant2 = 8'd37; b_mant3 = 8'd203;
a_exp0 = 10'd871; a_exp1 = 10'd526; a_exp2 = 10'd886; a_exp3 = 10'd155;
b_exp0 = 10'd981; b_exp1 = 10'd870; b_exp2 = 10'd454; b_exp3 = 10'd321;
a_sign0 = 4'd8; a_sign1 = 4'd15; a_sign2 = 4'd0; a_sign3 = 4'd1;
b_sign0 = 4'd8; b_sign1 = 4'd4; b_sign2 = 4'd11; b_sign3 = 4'd9;
@(posedge clk_i);
a_mant0 = 8'd98; a_mant1 = 8'd122; a_mant2 = 8'd120; a_mant3 = 8'd146;
b_mant0 = 8'd247; b_mant1 = 8'd29; b_mant2 = 8'd26; b_mant3 = 8'd86;
a_exp0 = 10'd506; a_exp1 = 10'd351; a_exp2 = 10'd83; a_exp3 = 10'd711;
b_exp0 = 10'd128; b_exp1 = 10'd625; b_exp2 = 10'd380; b_exp3 = 10'd76;
a_sign0 = 4'd12; a_sign1 = 4'd11; a_sign2 = 4'd6; a_sign3 = 4'd3;
b_sign0 = 4'd10; b_sign1 = 4'd10; b_sign2 = 4'd10; b_sign3 = 4'd12;
@(posedge clk_i);
shared_exps0 = 8'd121;
shared_exps1 = 8'd139;
rstn = 0;
@(posedge clk_i);
rstn = 1;
a_mant0 = 8'd195; a_mant1 = 8'd41; a_mant2 = 8'd133; a_mant3 = 8'd166;
b_mant0 = 8'd173; b_mant1 = 8'd51; b_mant2 = 8'd0; b_mant3 = 8'd113;
a_exp0 = 10'd842; a_exp1 = 10'd200; a_exp2 = 10'd171; a_exp3 = 10'd160;
b_exp0 = 10'd628; b_exp1 = 10'd786; b_exp2 = 10'd61; b_exp3 = 10'd604;
a_sign0 = 4'd0; a_sign1 = 4'd3; a_sign2 = 4'd10; a_sign3 = 4'd0;
b_sign0 = 4'd0; b_sign1 = 4'd0; b_sign2 = 4'd16; b_sign3 = 4'd4;
@(posedge clk_i);
a_mant0 = 8'd41; a_mant1 = 8'd177; a_mant2 = 8'd56; a_mant3 = 8'd8;
b_mant0 = 8'd61; b_mant1 = 8'd49; b_mant2 = 8'd82; b_mant3 = 8'd119;
a_exp0 = 10'd920; a_exp1 = 10'd25; a_exp2 = 10'd29; a_exp3 = 10'd232;
b_exp0 = 10'd821; b_exp1 = 10'd273; b_exp2 = 10'd436; b_exp3 = 10'd164;
a_sign0 = 4'd12; a_sign1 = 4'd10; a_sign2 = 4'd15; a_sign3 = 4'd6;
b_sign0 = 4'd11; b_sign1 = 4'd3; b_sign2 = 4'd3; b_sign3 = 4'd9;
@(posedge clk_i);
a_mant0 = 8'd180; a_mant1 = 8'd181; a_mant2 = 8'd45; a_mant3 = 8'd126;
b_mant0 = 8'd20; b_mant1 = 8'd210; b_mant2 = 8'd129; b_mant3 = 8'd6;
a_exp0 = 10'd477; a_exp1 = 10'd352; a_exp2 = 10'd91; a_exp3 = 10'd312;
b_exp0 = 10'd468; b_exp1 = 10'd86; b_exp2 = 10'd218; b_exp3 = 10'd899;
a_sign0 = 4'd13; a_sign1 = 4'd16; a_sign2 = 4'd3; a_sign3 = 4'd15;
b_sign0 = 4'd9; b_sign1 = 4'd0; b_sign2 = 4'd4; b_sign3 = 4'd10;
@(posedge clk_i);
a_mant0 = 8'd254; a_mant1 = 8'd22; a_mant2 = 8'd223; a_mant3 = 8'd183;
b_mant0 = 8'd95; b_mant1 = 8'd96; b_mant2 = 8'd94; b_mant3 = 8'd81;
a_exp0 = 10'd75; a_exp1 = 10'd307; a_exp2 = 10'd33; a_exp3 = 10'd120;
b_exp0 = 10'd195; b_exp1 = 10'd1022; b_exp2 = 10'd915; b_exp3 = 10'd767;
a_sign0 = 4'd6; a_sign1 = 4'd0; a_sign2 = 4'd4; a_sign3 = 4'd11;
b_sign0 = 4'd10; b_sign1 = 4'd8; b_sign2 = 4'd2; b_sign3 = 4'd0;
@(posedge clk_i);
a_mant0 = 8'd174; a_mant1 = 8'd125; a_mant2 = 8'd141; a_mant3 = 8'd89;
b_mant0 = 8'd189; b_mant1 = 8'd121; b_mant2 = 8'd125; b_mant3 = 8'd211;
a_exp0 = 10'd771; a_exp1 = 10'd614; a_exp2 = 10'd116; a_exp3 = 10'd1003;
b_exp0 = 10'd928; b_exp1 = 10'd51; b_exp2 = 10'd879; b_exp3 = 10'd899;
a_sign0 = 4'd11; a_sign1 = 4'd10; a_sign2 = 4'd11; a_sign3 = 4'd10;
b_sign0 = 4'd5; b_sign1 = 4'd15; b_sign2 = 4'd4; b_sign3 = 4'd7;
@(posedge clk_i);
a_mant0 = 8'd104; a_mant1 = 8'd124; a_mant2 = 8'd24; a_mant3 = 8'd116;
b_mant0 = 8'd27; b_mant1 = 8'd130; b_mant2 = 8'd184; b_mant3 = 8'd113;
a_exp0 = 10'd548; a_exp1 = 10'd132; a_exp2 = 10'd992; a_exp3 = 10'd449;
b_exp0 = 10'd983; b_exp1 = 10'd991; b_exp2 = 10'd541; b_exp3 = 10'd584;
a_sign0 = 4'd0; a_sign1 = 4'd8; a_sign2 = 4'd4; a_sign3 = 4'd10;
b_sign0 = 4'd12; b_sign1 = 4'd7; b_sign2 = 4'd13; b_sign3 = 4'd8;
@(posedge clk_i);
a_mant0 = 8'd217; a_mant1 = 8'd124; a_mant2 = 8'd168; a_mant3 = 8'd84;
b_mant0 = 8'd41; b_mant1 = 8'd223; b_mant2 = 8'd77; b_mant3 = 8'd220;
a_exp0 = 10'd173; a_exp1 = 10'd607; a_exp2 = 10'd324; a_exp3 = 10'd962;
b_exp0 = 10'd1017; b_exp1 = 10'd387; b_exp2 = 10'd198; b_exp3 = 10'd572;
a_sign0 = 4'd12; a_sign1 = 4'd11; a_sign2 = 4'd12; a_sign3 = 4'd10;
b_sign0 = 4'd4; b_sign1 = 4'd14; b_sign2 = 4'd3; b_sign3 = 4'd9;
@(posedge clk_i);
shared_exps0 = 8'd154;
shared_exps1 = 8'd131;
a_mant0 = 8'd67; a_mant1 = 8'd199; a_mant2 = 8'd188; a_mant3 = 8'd199;
b_mant0 = 8'd92; b_mant1 = 8'd224; b_mant2 = 8'd176; b_mant3 = 8'd136;
a_exp0 = 10'd429; a_exp1 = 10'd544; a_exp2 = 10'd1022; a_exp3 = 10'd18;
b_exp0 = 10'd302; b_exp1 = 10'd452; b_exp2 = 10'd825; b_exp3 = 10'd263;
a_sign0 = 4'd12; a_sign1 = 4'd10; a_sign2 = 4'd13; a_sign3 = 4'd2;
b_sign0 = 4'd7; b_sign1 = 4'd1; b_sign2 = 4'd4; b_sign3 = 4'd12;
@(posedge clk_i);
a_mant0 = 8'd124; a_mant1 = 8'd234; a_mant2 = 8'd111; a_mant3 = 8'd138;
b_mant0 = 8'd103; b_mant1 = 8'd61; b_mant2 = 8'd131; b_mant3 = 8'd128;
a_exp0 = 10'd67; a_exp1 = 10'd822; a_exp2 = 10'd182; a_exp3 = 10'd556;
b_exp0 = 10'd511; b_exp1 = 10'd487; b_exp2 = 10'd415; b_exp3 = 10'd874;
a_sign0 = 4'd1; a_sign1 = 4'd15; a_sign2 = 4'd12; a_sign3 = 4'd16;
b_sign0 = 4'd16; b_sign1 = 4'd11; b_sign2 = 4'd0; b_sign3 = 4'd11;
@(posedge clk_i);
a_mant0 = 8'd156; a_mant1 = 8'd164; a_mant2 = 8'd176; a_mant3 = 8'd190;
b_mant0 = 8'd242; b_mant1 = 8'd62; b_mant2 = 8'd37; b_mant3 = 8'd167;
a_exp0 = 10'd177; a_exp1 = 10'd727; a_exp2 = 10'd729; a_exp3 = 10'd834;
b_exp0 = 10'd503; b_exp1 = 10'd320; b_exp2 = 10'd1014; b_exp3 = 10'd133;
a_sign0 = 4'd13; a_sign1 = 4'd4; a_sign2 = 4'd14; a_sign3 = 4'd15;
b_sign0 = 4'd5; b_sign1 = 4'd12; b_sign2 = 4'd4; b_sign3 = 4'd2;
@(posedge clk_i);
a_mant0 = 8'd226; a_mant1 = 8'd62; a_mant2 = 8'd59; a_mant3 = 8'd203;
b_mant0 = 8'd3; b_mant1 = 8'd175; b_mant2 = 8'd242; b_mant3 = 8'd230;
a_exp0 = 10'd471; a_exp1 = 10'd738; a_exp2 = 10'd1023; a_exp3 = 10'd477;
b_exp0 = 10'd650; b_exp1 = 10'd86; b_exp2 = 10'd864; b_exp3 = 10'd648;
a_sign0 = 4'd16; a_sign1 = 4'd11; a_sign2 = 4'd16; a_sign3 = 4'd7;
b_sign0 = 4'd14; b_sign1 = 4'd7; b_sign2 = 4'd6; b_sign3 = 4'd8;
@(posedge clk_i);
a_mant0 = 8'd117; a_mant1 = 8'd190; a_mant2 = 8'd74; a_mant3 = 8'd85;
b_mant0 = 8'd82; b_mant1 = 8'd186; b_mant2 = 8'd212; b_mant3 = 8'd0;
a_exp0 = 10'd484; a_exp1 = 10'd103; a_exp2 = 10'd703; a_exp3 = 10'd309;
b_exp0 = 10'd559; b_exp1 = 10'd961; b_exp2 = 10'd433; b_exp3 = 10'd929;
a_sign0 = 4'd4; a_sign1 = 4'd16; a_sign2 = 4'd1; a_sign3 = 4'd2;
b_sign0 = 4'd11; b_sign1 = 4'd5; b_sign2 = 4'd10; b_sign3 = 4'd6;
@(posedge clk_i);
a_mant0 = 8'd146; a_mant1 = 8'd180; a_mant2 = 8'd71; a_mant3 = 8'd11;
b_mant0 = 8'd105; b_mant1 = 8'd223; b_mant2 = 8'd5; b_mant3 = 8'd231;
a_exp0 = 10'd822; a_exp1 = 10'd983; a_exp2 = 10'd128; a_exp3 = 10'd706;
b_exp0 = 10'd872; b_exp1 = 10'd1012; b_exp2 = 10'd356; b_exp3 = 10'd414;
a_sign0 = 4'd15; a_sign1 = 4'd1; a_sign2 = 4'd8; a_sign3 = 4'd11;
b_sign0 = 4'd3; b_sign1 = 4'd10; b_sign2 = 4'd1; b_sign3 = 4'd4;
@(posedge clk_i);
a_mant0 = 8'd109; a_mant1 = 8'd102; a_mant2 = 8'd227; a_mant3 = 8'd30;
b_mant0 = 8'd43; b_mant1 = 8'd201; b_mant2 = 8'd101; b_mant3 = 8'd206;
a_exp0 = 10'd861; a_exp1 = 10'd861; a_exp2 = 10'd485; a_exp3 = 10'd549;
b_exp0 = 10'd416; b_exp1 = 10'd170; b_exp2 = 10'd917; b_exp3 = 10'd540;
a_sign0 = 4'd4; a_sign1 = 4'd11; a_sign2 = 4'd16; a_sign3 = 4'd5;
b_sign0 = 4'd15; b_sign1 = 4'd3; b_sign2 = 4'd9; b_sign3 = 4'd9;
@(posedge clk_i);
a_mant0 = 8'd73; a_mant1 = 8'd210; a_mant2 = 8'd90; a_mant3 = 8'd182;
b_mant0 = 8'd138; b_mant1 = 8'd140; b_mant2 = 8'd66; b_mant3 = 8'd230;
a_exp0 = 10'd780; a_exp1 = 10'd9; a_exp2 = 10'd319; a_exp3 = 10'd148;
b_exp0 = 10'd175; b_exp1 = 10'd707; b_exp2 = 10'd426; b_exp3 = 10'd603;
a_sign0 = 4'd4; a_sign1 = 4'd4; a_sign2 = 4'd0; a_sign3 = 4'd10;
b_sign0 = 4'd7; b_sign1 = 4'd10; b_sign2 = 4'd15; b_sign3 = 4'd13;
@(posedge clk_i);
shared_exps0 = 8'd122;
shared_exps1 = 8'd136;
a_mant0 = 8'd135; a_mant1 = 8'd155; a_mant2 = 8'd43; a_mant3 = 8'd20;
b_mant0 = 8'd133; b_mant1 = 8'd17; b_mant2 = 8'd229; b_mant3 = 8'd243;
a_exp0 = 10'd496; a_exp1 = 10'd403; a_exp2 = 10'd876; a_exp3 = 10'd916;
b_exp0 = 10'd555; b_exp1 = 10'd506; b_exp2 = 10'd1002; b_exp3 = 10'd995;
a_sign0 = 4'd13; a_sign1 = 4'd2; a_sign2 = 4'd12; a_sign3 = 4'd15;
b_sign0 = 4'd15; b_sign1 = 4'd15; b_sign2 = 4'd7; b_sign3 = 4'd13;
@(posedge clk_i);
a_mant0 = 8'd115; a_mant1 = 8'd52; a_mant2 = 8'd197; a_mant3 = 8'd55;
b_mant0 = 8'd209; b_mant1 = 8'd211; b_mant2 = 8'd133; b_mant3 = 8'd31;
a_exp0 = 10'd32; a_exp1 = 10'd346; a_exp2 = 10'd571; a_exp3 = 10'd289;
b_exp0 = 10'd256; b_exp1 = 10'd969; b_exp2 = 10'd203; b_exp3 = 10'd466;
a_sign0 = 4'd16; a_sign1 = 4'd2; a_sign2 = 4'd8; a_sign3 = 4'd5;
b_sign0 = 4'd12; b_sign1 = 4'd7; b_sign2 = 4'd6; b_sign3 = 4'd9;
@(posedge clk_i);
a_mant0 = 8'd250; a_mant1 = 8'd117; a_mant2 = 8'd54; a_mant3 = 8'd112;
b_mant0 = 8'd60; b_mant1 = 8'd218; b_mant2 = 8'd61; b_mant3 = 8'd146;
a_exp0 = 10'd213; a_exp1 = 10'd84; a_exp2 = 10'd1003; a_exp3 = 10'd810;
b_exp0 = 10'd756; b_exp1 = 10'd739; b_exp2 = 10'd947; b_exp3 = 10'd390;
a_sign0 = 4'd13; a_sign1 = 4'd10; a_sign2 = 4'd11; a_sign3 = 4'd1;
b_sign0 = 4'd1; b_sign1 = 4'd13; b_sign2 = 4'd13; b_sign3 = 4'd1;
@(posedge clk_i);
a_mant0 = 8'd230; a_mant1 = 8'd96; a_mant2 = 8'd229; a_mant3 = 8'd76;
b_mant0 = 8'd119; b_mant1 = 8'd168; b_mant2 = 8'd218; b_mant3 = 8'd126;
a_exp0 = 10'd518; a_exp1 = 10'd492; a_exp2 = 10'd926; a_exp3 = 10'd1004;
b_exp0 = 10'd415; b_exp1 = 10'd417; b_exp2 = 10'd821; b_exp3 = 10'd277;
a_sign0 = 4'd3; a_sign1 = 4'd1; a_sign2 = 4'd6; a_sign3 = 4'd7;
b_sign0 = 4'd10; b_sign1 = 4'd3; b_sign2 = 4'd2; b_sign3 = 4'd5;
@(posedge clk_i);
a_mant0 = 8'd212; a_mant1 = 8'd48; a_mant2 = 8'd90; a_mant3 = 8'd46;
b_mant0 = 8'd213; b_mant1 = 8'd206; b_mant2 = 8'd97; b_mant3 = 8'd236;
a_exp0 = 10'd102; a_exp1 = 10'd815; a_exp2 = 10'd567; a_exp3 = 10'd439;
b_exp0 = 10'd204; b_exp1 = 10'd108; b_exp2 = 10'd381; b_exp3 = 10'd459;
a_sign0 = 4'd4; a_sign1 = 4'd12; a_sign2 = 4'd13; a_sign3 = 4'd1;
b_sign0 = 4'd16; b_sign1 = 4'd12; b_sign2 = 4'd3; b_sign3 = 4'd4;
@(posedge clk_i);
a_mant0 = 8'd1; a_mant1 = 8'd202; a_mant2 = 8'd86; a_mant3 = 8'd49;
b_mant0 = 8'd222; b_mant1 = 8'd31; b_mant2 = 8'd72; b_mant3 = 8'd182;
a_exp0 = 10'd946; a_exp1 = 10'd280; a_exp2 = 10'd946; a_exp3 = 10'd933;
b_exp0 = 10'd86; b_exp1 = 10'd892; b_exp2 = 10'd732; b_exp3 = 10'd341;
a_sign0 = 4'd7; a_sign1 = 4'd0; a_sign2 = 4'd4; a_sign3 = 4'd11;
b_sign0 = 4'd16; b_sign1 = 4'd8; b_sign2 = 4'd12; b_sign3 = 4'd16;
@(posedge clk_i);
a_mant0 = 8'd91; a_mant1 = 8'd134; a_mant2 = 8'd150; a_mant3 = 8'd216;
b_mant0 = 8'd246; b_mant1 = 8'd133; b_mant2 = 8'd150; b_mant3 = 8'd22;
a_exp0 = 10'd259; a_exp1 = 10'd147; a_exp2 = 10'd731; a_exp3 = 10'd531;
b_exp0 = 10'd56; b_exp1 = 10'd598; b_exp2 = 10'd497; b_exp3 = 10'd791;
a_sign0 = 4'd10; a_sign1 = 4'd6; a_sign2 = 4'd6; a_sign3 = 4'd8;
b_sign0 = 4'd15; b_sign1 = 4'd0; b_sign2 = 4'd7; b_sign3 = 4'd5;
@(posedge clk_i);
a_mant0 = 8'd23; a_mant1 = 8'd177; a_mant2 = 8'd48; a_mant3 = 8'd107;
b_mant0 = 8'd182; b_mant1 = 8'd80; b_mant2 = 8'd22; b_mant3 = 8'd74;
a_exp0 = 10'd312; a_exp1 = 10'd695; a_exp2 = 10'd148; a_exp3 = 10'd424;
b_exp0 = 10'd22; b_exp1 = 10'd832; b_exp2 = 10'd260; b_exp3 = 10'd485;
a_sign0 = 4'd6; a_sign1 = 4'd3; a_sign2 = 4'd5; a_sign3 = 4'd4;
b_sign0 = 4'd8; b_sign1 = 4'd7; b_sign2 = 4'd11; b_sign3 = 4'd9;
@(posedge clk_i);
shared_exps0 = 8'd124;
shared_exps1 = 8'd112;
a_mant0 = 8'd172; a_mant1 = 8'd101; a_mant2 = 8'd179; a_mant3 = 8'd207;
b_mant0 = 8'd195; b_mant1 = 8'd205; b_mant2 = 8'd86; b_mant3 = 8'd62;
a_exp0 = 10'd56; a_exp1 = 10'd899; a_exp2 = 10'd171; a_exp3 = 10'd911;
b_exp0 = 10'd1008; b_exp1 = 10'd161; b_exp2 = 10'd598; b_exp3 = 10'd844;
a_sign0 = 4'd16; a_sign1 = 4'd8; a_sign2 = 4'd16; a_sign3 = 4'd13;
b_sign0 = 4'd11; b_sign1 = 4'd11; b_sign2 = 4'd14; b_sign3 = 4'd3;
@(posedge clk_i);
a_mant0 = 8'd19; a_mant1 = 8'd218; a_mant2 = 8'd72; a_mant3 = 8'd70;
b_mant0 = 8'd73; b_mant1 = 8'd116; b_mant2 = 8'd0; b_mant3 = 8'd234;
a_exp0 = 10'd746; a_exp1 = 10'd354; a_exp2 = 10'd386; a_exp3 = 10'd419;
b_exp0 = 10'd424; b_exp1 = 10'd856; b_exp2 = 10'd899; b_exp3 = 10'd60;
a_sign0 = 4'd15; a_sign1 = 4'd1; a_sign2 = 4'd2; a_sign3 = 4'd3;
b_sign0 = 4'd0; b_sign1 = 4'd12; b_sign2 = 4'd3; b_sign3 = 4'd16;
@(posedge clk_i);
a_mant0 = 8'd234; a_mant1 = 8'd228; a_mant2 = 8'd149; a_mant3 = 8'd82;
b_mant0 = 8'd155; b_mant1 = 8'd0; b_mant2 = 8'd23; b_mant3 = 8'd152;
a_exp0 = 10'd793; a_exp1 = 10'd172; a_exp2 = 10'd275; a_exp3 = 10'd595;
b_exp0 = 10'd312; b_exp1 = 10'd989; b_exp2 = 10'd180; b_exp3 = 10'd242;
a_sign0 = 4'd10; a_sign1 = 4'd14; a_sign2 = 4'd9; a_sign3 = 4'd4;
b_sign0 = 4'd3; b_sign1 = 4'd14; b_sign2 = 4'd5; b_sign3 = 4'd13;
@(posedge clk_i);
a_mant0 = 8'd24; a_mant1 = 8'd84; a_mant2 = 8'd200; a_mant3 = 8'd197;
b_mant0 = 8'd32; b_mant1 = 8'd86; b_mant2 = 8'd181; b_mant3 = 8'd23;
a_exp0 = 10'd243; a_exp1 = 10'd129; a_exp2 = 10'd1004; a_exp3 = 10'd940;
b_exp0 = 10'd237; b_exp1 = 10'd822; b_exp2 = 10'd272; b_exp3 = 10'd841;
a_sign0 = 4'd14; a_sign1 = 4'd13; a_sign2 = 4'd13; a_sign3 = 4'd5;
b_sign0 = 4'd13; b_sign1 = 4'd11; b_sign2 = 4'd3; b_sign3 = 4'd10;
@(posedge clk_i);
a_mant0 = 8'd139; a_mant1 = 8'd210; a_mant2 = 8'd61; a_mant3 = 8'd7;
b_mant0 = 8'd84; b_mant1 = 8'd161; b_mant2 = 8'd130; b_mant3 = 8'd112;
a_exp0 = 10'd637; a_exp1 = 10'd852; a_exp2 = 10'd698; a_exp3 = 10'd686;
b_exp0 = 10'd588; b_exp1 = 10'd576; b_exp2 = 10'd55; b_exp3 = 10'd982;
a_sign0 = 4'd15; a_sign1 = 4'd14; a_sign2 = 4'd9; a_sign3 = 4'd14;
b_sign0 = 4'd8; b_sign1 = 4'd1; b_sign2 = 4'd0; b_sign3 = 4'd9;
@(posedge clk_i);
a_mant0 = 8'd63; a_mant1 = 8'd43; a_mant2 = 8'd165; a_mant3 = 8'd138;
b_mant0 = 8'd222; b_mant1 = 8'd150; b_mant2 = 8'd10; b_mant3 = 8'd118;
a_exp0 = 10'd46; a_exp1 = 10'd1013; a_exp2 = 10'd661; a_exp3 = 10'd887;
b_exp0 = 10'd306; b_exp1 = 10'd626; b_exp2 = 10'd443; b_exp3 = 10'd406;
a_sign0 = 4'd12; a_sign1 = 4'd14; a_sign2 = 4'd13; a_sign3 = 4'd2;
b_sign0 = 4'd13; b_sign1 = 4'd10; b_sign2 = 4'd4; b_sign3 = 4'd2;
@(posedge clk_i);
a_mant0 = 8'd90; a_mant1 = 8'd2; a_mant2 = 8'd214; a_mant3 = 8'd208;
b_mant0 = 8'd186; b_mant1 = 8'd224; b_mant2 = 8'd5; b_mant3 = 8'd8;
a_exp0 = 10'd456; a_exp1 = 10'd99; a_exp2 = 10'd631; a_exp3 = 10'd713;
b_exp0 = 10'd866; b_exp1 = 10'd273; b_exp2 = 10'd732; b_exp3 = 10'd54;
a_sign0 = 4'd8; a_sign1 = 4'd3; a_sign2 = 4'd5; a_sign3 = 4'd2;
b_sign0 = 4'd16; b_sign1 = 4'd5; b_sign2 = 4'd2; b_sign3 = 4'd14;
@(posedge clk_i);
a_mant0 = 8'd128; a_mant1 = 8'd26; a_mant2 = 8'd225; a_mant3 = 8'd186;
b_mant0 = 8'd245; b_mant1 = 8'd124; b_mant2 = 8'd187; b_mant3 = 8'd179;
a_exp0 = 10'd955; a_exp1 = 10'd866; a_exp2 = 10'd148; a_exp3 = 10'd812;
b_exp0 = 10'd340; b_exp1 = 10'd950; b_exp2 = 10'd642; b_exp3 = 10'd411;
a_sign0 = 4'd15; a_sign1 = 4'd11; a_sign2 = 4'd4; a_sign3 = 4'd15;
b_sign0 = 4'd16; b_sign1 = 4'd3; b_sign2 = 4'd10; b_sign3 = 4'd8;
@(posedge clk_i);
shared_exps0 = 8'd138;
shared_exps1 = 8'd129;
rstn = 0;
@(posedge clk_i);
rstn = 1;
a_mant0 = 8'd168; a_mant1 = 8'd62; a_mant2 = 8'd36; a_mant3 = 8'd86;
b_mant0 = 8'd240; b_mant1 = 8'd66; b_mant2 = 8'd62; b_mant3 = 8'd247;
a_exp0 = 10'd365; a_exp1 = 10'd821; a_exp2 = 10'd776; a_exp3 = 10'd644;
b_exp0 = 10'd460; b_exp1 = 10'd685; b_exp2 = 10'd520; b_exp3 = 10'd148;
a_sign0 = 4'd4; a_sign1 = 4'd13; a_sign2 = 4'd5; a_sign3 = 4'd2;
b_sign0 = 4'd5; b_sign1 = 4'd16; b_sign2 = 4'd9; b_sign3 = 4'd10;
@(posedge clk_i);
a_mant0 = 8'd124; a_mant1 = 8'd173; a_mant2 = 8'd163; a_mant3 = 8'd100;
b_mant0 = 8'd193; b_mant1 = 8'd174; b_mant2 = 8'd138; b_mant3 = 8'd72;
a_exp0 = 10'd703; a_exp1 = 10'd757; a_exp2 = 10'd810; a_exp3 = 10'd563;
b_exp0 = 10'd656; b_exp1 = 10'd108; b_exp2 = 10'd964; b_exp3 = 10'd704;
a_sign0 = 4'd8; a_sign1 = 4'd4; a_sign2 = 4'd6; a_sign3 = 4'd14;
b_sign0 = 4'd1; b_sign1 = 4'd15; b_sign2 = 4'd15; b_sign3 = 4'd3;
@(posedge clk_i);
a_mant0 = 8'd64; a_mant1 = 8'd229; a_mant2 = 8'd110; a_mant3 = 8'd49;
b_mant0 = 8'd74; b_mant1 = 8'd147; b_mant2 = 8'd38; b_mant3 = 8'd161;
a_exp0 = 10'd42; a_exp1 = 10'd367; a_exp2 = 10'd712; a_exp3 = 10'd453;
b_exp0 = 10'd279; b_exp1 = 10'd105; b_exp2 = 10'd9; b_exp3 = 10'd681;
a_sign0 = 4'd3; a_sign1 = 4'd16; a_sign2 = 4'd3; a_sign3 = 4'd2;
b_sign0 = 4'd8; b_sign1 = 4'd9; b_sign2 = 4'd8; b_sign3 = 4'd11;
@(posedge clk_i);
a_mant0 = 8'd55; a_mant1 = 8'd6; a_mant2 = 8'd204; a_mant3 = 8'd117;
b_mant0 = 8'd109; b_mant1 = 8'd162; b_mant2 = 8'd245; b_mant3 = 8'd128;
a_exp0 = 10'd162; a_exp1 = 10'd106; a_exp2 = 10'd592; a_exp3 = 10'd383;
b_exp0 = 10'd916; b_exp1 = 10'd252; b_exp2 = 10'd170; b_exp3 = 10'd96;
a_sign0 = 4'd7; a_sign1 = 4'd11; a_sign2 = 4'd8; a_sign3 = 4'd6;
b_sign0 = 4'd12; b_sign1 = 4'd9; b_sign2 = 4'd12; b_sign3 = 4'd8;
@(posedge clk_i);
a_mant0 = 8'd67; a_mant1 = 8'd47; a_mant2 = 8'd43; a_mant3 = 8'd39;
b_mant0 = 8'd181; b_mant1 = 8'd238; b_mant2 = 8'd193; b_mant3 = 8'd231;
a_exp0 = 10'd989; a_exp1 = 10'd988; a_exp2 = 10'd532; a_exp3 = 10'd203;
b_exp0 = 10'd86; b_exp1 = 10'd504; b_exp2 = 10'd761; b_exp3 = 10'd776;
a_sign0 = 4'd12; a_sign1 = 4'd1; a_sign2 = 4'd9; a_sign3 = 4'd8;
b_sign0 = 4'd11; b_sign1 = 4'd16; b_sign2 = 4'd12; b_sign3 = 4'd0;
@(posedge clk_i);
a_mant0 = 8'd69; a_mant1 = 8'd253; a_mant2 = 8'd211; a_mant3 = 8'd129;
b_mant0 = 8'd137; b_mant1 = 8'd155; b_mant2 = 8'd102; b_mant3 = 8'd26;
a_exp0 = 10'd624; a_exp1 = 10'd787; a_exp2 = 10'd1008; a_exp3 = 10'd543;
b_exp0 = 10'd117; b_exp1 = 10'd966; b_exp2 = 10'd808; b_exp3 = 10'd691;
a_sign0 = 4'd5; a_sign1 = 4'd10; a_sign2 = 4'd5; a_sign3 = 4'd1;
b_sign0 = 4'd5; b_sign1 = 4'd0; b_sign2 = 4'd1; b_sign3 = 4'd1;
@(posedge clk_i);
a_mant0 = 8'd28; a_mant1 = 8'd188; a_mant2 = 8'd201; a_mant3 = 8'd253;
b_mant0 = 8'd6; b_mant1 = 8'd150; b_mant2 = 8'd194; b_mant3 = 8'd113;
a_exp0 = 10'd128; a_exp1 = 10'd726; a_exp2 = 10'd865; a_exp3 = 10'd246;
b_exp0 = 10'd653; b_exp1 = 10'd515; b_exp2 = 10'd350; b_exp3 = 10'd504;
a_sign0 = 4'd12; a_sign1 = 4'd10; a_sign2 = 4'd7; a_sign3 = 4'd11;
b_sign0 = 4'd1; b_sign1 = 4'd3; b_sign2 = 4'd0; b_sign3 = 4'd13;
@(posedge clk_i);
shared_exps0 = 8'd120;
shared_exps1 = 8'd108;
a_mant0 = 8'd134; a_mant1 = 8'd21; a_mant2 = 8'd122; a_mant3 = 8'd17;
b_mant0 = 8'd0; b_mant1 = 8'd96; b_mant2 = 8'd187; b_mant3 = 8'd146;
a_exp0 = 10'd253; a_exp1 = 10'd373; a_exp2 = 10'd245; a_exp3 = 10'd542;
b_exp0 = 10'd654; b_exp1 = 10'd266; b_exp2 = 10'd42; b_exp3 = 10'd96;
a_sign0 = 4'd8; a_sign1 = 4'd5; a_sign2 = 4'd8; a_sign3 = 4'd12;
b_sign0 = 4'd8; b_sign1 = 4'd6; b_sign2 = 4'd16; b_sign3 = 4'd4;
@(posedge clk_i);
a_mant0 = 8'd184; a_mant1 = 8'd180; a_mant2 = 8'd125; a_mant3 = 8'd87;
b_mant0 = 8'd131; b_mant1 = 8'd231; b_mant2 = 8'd6; b_mant3 = 8'd52;
a_exp0 = 10'd576; a_exp1 = 10'd196; a_exp2 = 10'd811; a_exp3 = 10'd897;
b_exp0 = 10'd319; b_exp1 = 10'd874; b_exp2 = 10'd728; b_exp3 = 10'd447;
a_sign0 = 4'd3; a_sign1 = 4'd5; a_sign2 = 4'd7; a_sign3 = 4'd14;
b_sign0 = 4'd3; b_sign1 = 4'd9; b_sign2 = 4'd12; b_sign3 = 4'd11;
@(posedge clk_i);
a_mant0 = 8'd28; a_mant1 = 8'd229; a_mant2 = 8'd228; a_mant3 = 8'd235;
b_mant0 = 8'd205; b_mant1 = 8'd118; b_mant2 = 8'd102; b_mant3 = 8'd123;
a_exp0 = 10'd233; a_exp1 = 10'd787; a_exp2 = 10'd967; a_exp3 = 10'd619;
b_exp0 = 10'd140; b_exp1 = 10'd241; b_exp2 = 10'd956; b_exp3 = 10'd738;
a_sign0 = 4'd16; a_sign1 = 4'd12; a_sign2 = 4'd6; a_sign3 = 4'd8;
b_sign0 = 4'd13; b_sign1 = 4'd11; b_sign2 = 4'd11; b_sign3 = 4'd1;
@(posedge clk_i);
a_mant0 = 8'd14; a_mant1 = 8'd155; a_mant2 = 8'd34; a_mant3 = 8'd152;
b_mant0 = 8'd253; b_mant1 = 8'd233; b_mant2 = 8'd57; b_mant3 = 8'd9;
a_exp0 = 10'd633; a_exp1 = 10'd1001; a_exp2 = 10'd943; a_exp3 = 10'd951;
b_exp0 = 10'd661; b_exp1 = 10'd490; b_exp2 = 10'd998; b_exp3 = 10'd746;
a_sign0 = 4'd0; a_sign1 = 4'd15; a_sign2 = 4'd3; a_sign3 = 4'd2;
b_sign0 = 4'd5; b_sign1 = 4'd9; b_sign2 = 4'd3; b_sign3 = 4'd15;
@(posedge clk_i);
a_mant0 = 8'd64; a_mant1 = 8'd32; a_mant2 = 8'd11; a_mant3 = 8'd255;
b_mant0 = 8'd71; b_mant1 = 8'd47; b_mant2 = 8'd197; b_mant3 = 8'd37;
a_exp0 = 10'd842; a_exp1 = 10'd388; a_exp2 = 10'd785; a_exp3 = 10'd935;
b_exp0 = 10'd501; b_exp1 = 10'd391; b_exp2 = 10'd569; b_exp3 = 10'd924;
a_sign0 = 4'd12; a_sign1 = 4'd6; a_sign2 = 4'd9; a_sign3 = 4'd4;
b_sign0 = 4'd11; b_sign1 = 4'd6; b_sign2 = 4'd11; b_sign3 = 4'd9;
@(posedge clk_i);
a_mant0 = 8'd227; a_mant1 = 8'd100; a_mant2 = 8'd48; a_mant3 = 8'd125;
b_mant0 = 8'd143; b_mant1 = 8'd66; b_mant2 = 8'd66; b_mant3 = 8'd195;
a_exp0 = 10'd13; a_exp1 = 10'd120; a_exp2 = 10'd928; a_exp3 = 10'd481;
b_exp0 = 10'd480; b_exp1 = 10'd62; b_exp2 = 10'd430; b_exp3 = 10'd941;
a_sign0 = 4'd9; a_sign1 = 4'd15; a_sign2 = 4'd2; a_sign3 = 4'd6;
b_sign0 = 4'd14; b_sign1 = 4'd12; b_sign2 = 4'd9; b_sign3 = 4'd14;
@(posedge clk_i);
a_mant0 = 8'd138; a_mant1 = 8'd10; a_mant2 = 8'd231; a_mant3 = 8'd119;
b_mant0 = 8'd83; b_mant1 = 8'd114; b_mant2 = 8'd188; b_mant3 = 8'd234;
a_exp0 = 10'd140; a_exp1 = 10'd39; a_exp2 = 10'd621; a_exp3 = 10'd1012;
b_exp0 = 10'd96; b_exp1 = 10'd820; b_exp2 = 10'd223; b_exp3 = 10'd639;
a_sign0 = 4'd8; a_sign1 = 4'd6; a_sign2 = 4'd8; a_sign3 = 4'd4;
b_sign0 = 4'd10; b_sign1 = 4'd3; b_sign2 = 4'd14; b_sign3 = 4'd6;
@(posedge clk_i);
a_mant0 = 8'd137; a_mant1 = 8'd31; a_mant2 = 8'd118; a_mant3 = 8'd106;
b_mant0 = 8'd239; b_mant1 = 8'd202; b_mant2 = 8'd32; b_mant3 = 8'd109;
a_exp0 = 10'd137; a_exp1 = 10'd714; a_exp2 = 10'd549; a_exp3 = 10'd35;
b_exp0 = 10'd763; b_exp1 = 10'd880; b_exp2 = 10'd584; b_exp3 = 10'd561;
a_sign0 = 4'd15; a_sign1 = 4'd8; a_sign2 = 4'd1; a_sign3 = 4'd13;
b_sign0 = 4'd0; b_sign1 = 4'd15; b_sign2 = 4'd10; b_sign3 = 4'd2;
@(posedge clk_i);
shared_exps0 = 8'd145;
shared_exps1 = 8'd139;
a_mant0 = 8'd77; a_mant1 = 8'd140; a_mant2 = 8'd51; a_mant3 = 8'd46;
b_mant0 = 8'd234; b_mant1 = 8'd209; b_mant2 = 8'd167; b_mant3 = 8'd206;
a_exp0 = 10'd13; a_exp1 = 10'd397; a_exp2 = 10'd64; a_exp3 = 10'd641;
b_exp0 = 10'd419; b_exp1 = 10'd767; b_exp2 = 10'd1023; b_exp3 = 10'd939;
a_sign0 = 4'd13; a_sign1 = 4'd12; a_sign2 = 4'd16; a_sign3 = 4'd3;
b_sign0 = 4'd0; b_sign1 = 4'd6; b_sign2 = 4'd6; b_sign3 = 4'd9;
@(posedge clk_i);
a_mant0 = 8'd255; a_mant1 = 8'd145; a_mant2 = 8'd170; a_mant3 = 8'd61;
b_mant0 = 8'd106; b_mant1 = 8'd142; b_mant2 = 8'd9; b_mant3 = 8'd145;
a_exp0 = 10'd209; a_exp1 = 10'd369; a_exp2 = 10'd792; a_exp3 = 10'd797;
b_exp0 = 10'd725; b_exp1 = 10'd792; b_exp2 = 10'd984; b_exp3 = 10'd768;
a_sign0 = 4'd5; a_sign1 = 4'd1; a_sign2 = 4'd1; a_sign3 = 4'd4;
b_sign0 = 4'd10; b_sign1 = 4'd1; b_sign2 = 4'd0; b_sign3 = 4'd7;
@(posedge clk_i);
a_mant0 = 8'd22; a_mant1 = 8'd104; a_mant2 = 8'd204; a_mant3 = 8'd255;
b_mant0 = 8'd79; b_mant1 = 8'd182; b_mant2 = 8'd187; b_mant3 = 8'd217;
a_exp0 = 10'd231; a_exp1 = 10'd942; a_exp2 = 10'd551; a_exp3 = 10'd442;
b_exp0 = 10'd257; b_exp1 = 10'd74; b_exp2 = 10'd707; b_exp3 = 10'd176;
a_sign0 = 4'd6; a_sign1 = 4'd4; a_sign2 = 4'd12; a_sign3 = 4'd8;
b_sign0 = 4'd9; b_sign1 = 4'd11; b_sign2 = 4'd6; b_sign3 = 4'd5;
@(posedge clk_i);
a_mant0 = 8'd65; a_mant1 = 8'd14; a_mant2 = 8'd242; a_mant3 = 8'd235;
b_mant0 = 8'd249; b_mant1 = 8'd210; b_mant2 = 8'd107; b_mant3 = 8'd97;
a_exp0 = 10'd483; a_exp1 = 10'd806; a_exp2 = 10'd385; a_exp3 = 10'd669;
b_exp0 = 10'd983; b_exp1 = 10'd994; b_exp2 = 10'd896; b_exp3 = 10'd268;
a_sign0 = 4'd2; a_sign1 = 4'd11; a_sign2 = 4'd6; a_sign3 = 4'd9;
b_sign0 = 4'd11; b_sign1 = 4'd7; b_sign2 = 4'd7; b_sign3 = 4'd2;
@(posedge clk_i);
a_mant0 = 8'd95; a_mant1 = 8'd210; a_mant2 = 8'd140; a_mant3 = 8'd172;
b_mant0 = 8'd162; b_mant1 = 8'd9; b_mant2 = 8'd238; b_mant3 = 8'd208;
a_exp0 = 10'd967; a_exp1 = 10'd934; a_exp2 = 10'd777; a_exp3 = 10'd547;
b_exp0 = 10'd876; b_exp1 = 10'd149; b_exp2 = 10'd443; b_exp3 = 10'd432;
a_sign0 = 4'd3; a_sign1 = 4'd6; a_sign2 = 4'd14; a_sign3 = 4'd4;
b_sign0 = 4'd9; b_sign1 = 4'd5; b_sign2 = 4'd1; b_sign3 = 4'd9;
@(posedge clk_i);
a_mant0 = 8'd4; a_mant1 = 8'd94; a_mant2 = 8'd65; a_mant3 = 8'd55;
b_mant0 = 8'd194; b_mant1 = 8'd149; b_mant2 = 8'd43; b_mant3 = 8'd222;
a_exp0 = 10'd490; a_exp1 = 10'd539; a_exp2 = 10'd882; a_exp3 = 10'd962;
b_exp0 = 10'd721; b_exp1 = 10'd310; b_exp2 = 10'd452; b_exp3 = 10'd332;
a_sign0 = 4'd2; a_sign1 = 4'd10; a_sign2 = 4'd3; a_sign3 = 4'd5;
b_sign0 = 4'd8; b_sign1 = 4'd6; b_sign2 = 4'd6; b_sign3 = 4'd3;
@(posedge clk_i);
a_mant0 = 8'd70; a_mant1 = 8'd160; a_mant2 = 8'd21; a_mant3 = 8'd139;
b_mant0 = 8'd201; b_mant1 = 8'd85; b_mant2 = 8'd36; b_mant3 = 8'd101;
a_exp0 = 10'd899; a_exp1 = 10'd659; a_exp2 = 10'd422; a_exp3 = 10'd238;
b_exp0 = 10'd920; b_exp1 = 10'd578; b_exp2 = 10'd461; b_exp3 = 10'd309;
a_sign0 = 4'd14; a_sign1 = 4'd15; a_sign2 = 4'd15; a_sign3 = 4'd13;
b_sign0 = 4'd6; b_sign1 = 4'd5; b_sign2 = 4'd3; b_sign3 = 4'd15;
@(posedge clk_i);
a_mant0 = 8'd208; a_mant1 = 8'd10; a_mant2 = 8'd157; a_mant3 = 8'd218;
b_mant0 = 8'd197; b_mant1 = 8'd86; b_mant2 = 8'd240; b_mant3 = 8'd69;
a_exp0 = 10'd417; a_exp1 = 10'd933; a_exp2 = 10'd298; a_exp3 = 10'd37;
b_exp0 = 10'd135; b_exp1 = 10'd512; b_exp2 = 10'd533; b_exp3 = 10'd547;
a_sign0 = 4'd16; a_sign1 = 4'd3; a_sign2 = 4'd15; a_sign3 = 4'd0;
b_sign0 = 4'd1; b_sign1 = 4'd5; b_sign2 = 4'd9; b_sign3 = 4'd6;
@(posedge clk_i);
shared_exps0 = 8'd164;
shared_exps1 = 8'd123;
a_mant0 = 8'd64; a_mant1 = 8'd8; a_mant2 = 8'd50; a_mant3 = 8'd138;
b_mant0 = 8'd85; b_mant1 = 8'd106; b_mant2 = 8'd108; b_mant3 = 8'd59;
a_exp0 = 10'd881; a_exp1 = 10'd794; a_exp2 = 10'd899; a_exp3 = 10'd687;
b_exp0 = 10'd593; b_exp1 = 10'd490; b_exp2 = 10'd893; b_exp3 = 10'd297;
a_sign0 = 4'd16; a_sign1 = 4'd9; a_sign2 = 4'd15; a_sign3 = 4'd4;
b_sign0 = 4'd5; b_sign1 = 4'd15; b_sign2 = 4'd11; b_sign3 = 4'd3;
@(posedge clk_i);
a_mant0 = 8'd107; a_mant1 = 8'd90; a_mant2 = 8'd155; a_mant3 = 8'd86;
b_mant0 = 8'd180; b_mant1 = 8'd252; b_mant2 = 8'd168; b_mant3 = 8'd127;
a_exp0 = 10'd710; a_exp1 = 10'd410; a_exp2 = 10'd202; a_exp3 = 10'd383;
b_exp0 = 10'd412; b_exp1 = 10'd789; b_exp2 = 10'd198; b_exp3 = 10'd134;
a_sign0 = 4'd8; a_sign1 = 4'd14; a_sign2 = 4'd16; a_sign3 = 4'd13;
b_sign0 = 4'd5; b_sign1 = 4'd13; b_sign2 = 4'd15; b_sign3 = 4'd7;
@(posedge clk_i);
a_mant0 = 8'd219; a_mant1 = 8'd28; a_mant2 = 8'd71; a_mant3 = 8'd245;
b_mant0 = 8'd166; b_mant1 = 8'd174; b_mant2 = 8'd148; b_mant3 = 8'd58;
a_exp0 = 10'd924; a_exp1 = 10'd818; a_exp2 = 10'd705; a_exp3 = 10'd12;
b_exp0 = 10'd482; b_exp1 = 10'd14; b_exp2 = 10'd746; b_exp3 = 10'd296;
a_sign0 = 4'd5; a_sign1 = 4'd5; a_sign2 = 4'd7; a_sign3 = 4'd10;
b_sign0 = 4'd13; b_sign1 = 4'd4; b_sign2 = 4'd9; b_sign3 = 4'd3;
@(posedge clk_i);
a_mant0 = 8'd191; a_mant1 = 8'd170; a_mant2 = 8'd14; a_mant3 = 8'd148;
b_mant0 = 8'd83; b_mant1 = 8'd183; b_mant2 = 8'd110; b_mant3 = 8'd195;
a_exp0 = 10'd733; a_exp1 = 10'd251; a_exp2 = 10'd76; a_exp3 = 10'd516;
b_exp0 = 10'd252; b_exp1 = 10'd54; b_exp2 = 10'd17; b_exp3 = 10'd532;
a_sign0 = 4'd13; a_sign1 = 4'd0; a_sign2 = 4'd4; a_sign3 = 4'd16;
b_sign0 = 4'd0; b_sign1 = 4'd3; b_sign2 = 4'd8; b_sign3 = 4'd5;
@(posedge clk_i);
a_mant0 = 8'd99; a_mant1 = 8'd18; a_mant2 = 8'd155; a_mant3 = 8'd47;
b_mant0 = 8'd59; b_mant1 = 8'd183; b_mant2 = 8'd250; b_mant3 = 8'd216;
a_exp0 = 10'd486; a_exp1 = 10'd992; a_exp2 = 10'd916; a_exp3 = 10'd297;
b_exp0 = 10'd851; b_exp1 = 10'd498; b_exp2 = 10'd328; b_exp3 = 10'd519;
a_sign0 = 4'd6; a_sign1 = 4'd10; a_sign2 = 4'd0; a_sign3 = 4'd15;
b_sign0 = 4'd15; b_sign1 = 4'd1; b_sign2 = 4'd10; b_sign3 = 4'd16;
@(posedge clk_i);
a_mant0 = 8'd189; a_mant1 = 8'd4; a_mant2 = 8'd45; a_mant3 = 8'd113;
b_mant0 = 8'd178; b_mant1 = 8'd14; b_mant2 = 8'd137; b_mant3 = 8'd29;
a_exp0 = 10'd819; a_exp1 = 10'd497; a_exp2 = 10'd181; a_exp3 = 10'd302;
b_exp0 = 10'd915; b_exp1 = 10'd192; b_exp2 = 10'd82; b_exp3 = 10'd28;
a_sign0 = 4'd3; a_sign1 = 4'd15; a_sign2 = 4'd6; a_sign3 = 4'd10;
b_sign0 = 4'd1; b_sign1 = 4'd0; b_sign2 = 4'd16; b_sign3 = 4'd11;
@(posedge clk_i);
a_mant0 = 8'd115; a_mant1 = 8'd76; a_mant2 = 8'd112; a_mant3 = 8'd114;
b_mant0 = 8'd108; b_mant1 = 8'd203; b_mant2 = 8'd46; b_mant3 = 8'd94;
a_exp0 = 10'd81; a_exp1 = 10'd645; a_exp2 = 10'd161; a_exp3 = 10'd599;
b_exp0 = 10'd123; b_exp1 = 10'd180; b_exp2 = 10'd940; b_exp3 = 10'd148;
a_sign0 = 4'd9; a_sign1 = 4'd2; a_sign2 = 4'd10; a_sign3 = 4'd0;
b_sign0 = 4'd11; b_sign1 = 4'd2; b_sign2 = 4'd9; b_sign3 = 4'd0;
@(posedge clk_i);
a_mant0 = 8'd137; a_mant1 = 8'd188; a_mant2 = 8'd179; a_mant3 = 8'd188;
b_mant0 = 8'd120; b_mant1 = 8'd150; b_mant2 = 8'd114; b_mant3 = 8'd145;
a_exp0 = 10'd321; a_exp1 = 10'd203; a_exp2 = 10'd490; a_exp3 = 10'd586;
b_exp0 = 10'd608; b_exp1 = 10'd667; b_exp2 = 10'd426; b_exp3 = 10'd292;
a_sign0 = 4'd2; a_sign1 = 4'd13; a_sign2 = 4'd0; a_sign3 = 4'd3;
b_sign0 = 4'd4; b_sign1 = 4'd0; b_sign2 = 4'd7; b_sign3 = 4'd7;
@(posedge clk_i);
shared_exps0 = 8'd104;
shared_exps1 = 8'd129;
rstn = 0;
@(posedge clk_i);
rstn = 1;
a_mant0 = 8'd160; a_mant1 = 8'd244; a_mant2 = 8'd252; a_mant3 = 8'd40;
b_mant0 = 8'd245; b_mant1 = 8'd106; b_mant2 = 8'd156; b_mant3 = 8'd71;
a_exp0 = 10'd431; a_exp1 = 10'd284; a_exp2 = 10'd705; a_exp3 = 10'd847;
b_exp0 = 10'd154; b_exp1 = 10'd872; b_exp2 = 10'd622; b_exp3 = 10'd923;
a_sign0 = 4'd9; a_sign1 = 4'd14; a_sign2 = 4'd4; a_sign3 = 4'd0;
b_sign0 = 4'd9; b_sign1 = 4'd4; b_sign2 = 4'd12; b_sign3 = 4'd2;
@(posedge clk_i);
a_mant0 = 8'd236; a_mant1 = 8'd34; a_mant2 = 8'd21; a_mant3 = 8'd10;
b_mant0 = 8'd113; b_mant1 = 8'd40; b_mant2 = 8'd223; b_mant3 = 8'd198;
a_exp0 = 10'd708; a_exp1 = 10'd720; a_exp2 = 10'd923; a_exp3 = 10'd861;
b_exp0 = 10'd491; b_exp1 = 10'd375; b_exp2 = 10'd824; b_exp3 = 10'd358;
a_sign0 = 4'd13; a_sign1 = 4'd9; a_sign2 = 4'd16; a_sign3 = 4'd12;
b_sign0 = 4'd8; b_sign1 = 4'd6; b_sign2 = 4'd6; b_sign3 = 4'd2;
@(posedge clk_i);
a_mant0 = 8'd242; a_mant1 = 8'd206; a_mant2 = 8'd100; a_mant3 = 8'd69;
b_mant0 = 8'd153; b_mant1 = 8'd203; b_mant2 = 8'd203; b_mant3 = 8'd238;
a_exp0 = 10'd469; a_exp1 = 10'd239; a_exp2 = 10'd604; a_exp3 = 10'd934;
b_exp0 = 10'd994; b_exp1 = 10'd651; b_exp2 = 10'd970; b_exp3 = 10'd611;
a_sign0 = 4'd0; a_sign1 = 4'd13; a_sign2 = 4'd0; a_sign3 = 4'd8;
b_sign0 = 4'd1; b_sign1 = 4'd1; b_sign2 = 4'd9; b_sign3 = 4'd8;
@(posedge clk_i);
a_mant0 = 8'd22; a_mant1 = 8'd230; a_mant2 = 8'd219; a_mant3 = 8'd60;
b_mant0 = 8'd114; b_mant1 = 8'd162; b_mant2 = 8'd3; b_mant3 = 8'd146;
a_exp0 = 10'd139; a_exp1 = 10'd716; a_exp2 = 10'd376; a_exp3 = 10'd753;
b_exp0 = 10'd584; b_exp1 = 10'd594; b_exp2 = 10'd580; b_exp3 = 10'd421;
a_sign0 = 4'd6; a_sign1 = 4'd0; a_sign2 = 4'd1; a_sign3 = 4'd4;
b_sign0 = 4'd13; b_sign1 = 4'd10; b_sign2 = 4'd3; b_sign3 = 4'd16;
@(posedge clk_i);
a_mant0 = 8'd79; a_mant1 = 8'd24; a_mant2 = 8'd50; a_mant3 = 8'd147;
b_mant0 = 8'd61; b_mant1 = 8'd249; b_mant2 = 8'd248; b_mant3 = 8'd186;
a_exp0 = 10'd605; a_exp1 = 10'd254; a_exp2 = 10'd637; a_exp3 = 10'd150;
b_exp0 = 10'd620; b_exp1 = 10'd122; b_exp2 = 10'd755; b_exp3 = 10'd179;
a_sign0 = 4'd7; a_sign1 = 4'd11; a_sign2 = 4'd2; a_sign3 = 4'd8;
b_sign0 = 4'd5; b_sign1 = 4'd2; b_sign2 = 4'd10; b_sign3 = 4'd10;
@(posedge clk_i);
a_mant0 = 8'd118; a_mant1 = 8'd139; a_mant2 = 8'd234; a_mant3 = 8'd55;
b_mant0 = 8'd11; b_mant1 = 8'd54; b_mant2 = 8'd116; b_mant3 = 8'd168;
a_exp0 = 10'd993; a_exp1 = 10'd844; a_exp2 = 10'd820; a_exp3 = 10'd17;
b_exp0 = 10'd648; b_exp1 = 10'd475; b_exp2 = 10'd864; b_exp3 = 10'd1004;
a_sign0 = 4'd8; a_sign1 = 4'd15; a_sign2 = 4'd7; a_sign3 = 4'd11;
b_sign0 = 4'd12; b_sign1 = 4'd15; b_sign2 = 4'd11; b_sign3 = 4'd9;
@(posedge clk_i);
a_mant0 = 8'd211; a_mant1 = 8'd252; a_mant2 = 8'd14; a_mant3 = 8'd141;
b_mant0 = 8'd105; b_mant1 = 8'd34; b_mant2 = 8'd163; b_mant3 = 8'd228;
a_exp0 = 10'd791; a_exp1 = 10'd914; a_exp2 = 10'd294; a_exp3 = 10'd299;
b_exp0 = 10'd343; b_exp1 = 10'd71; b_exp2 = 10'd988; b_exp3 = 10'd940;
a_sign0 = 4'd13; a_sign1 = 4'd9; a_sign2 = 4'd14; a_sign3 = 4'd8;
b_sign0 = 4'd12; b_sign1 = 4'd1; b_sign2 = 4'd15; b_sign3 = 4'd1;
@(posedge clk_i);
shared_exps0 = 8'd90;
shared_exps1 = 8'd149;
a_mant0 = 8'd55; a_mant1 = 8'd121; a_mant2 = 8'd223; a_mant3 = 8'd145;
b_mant0 = 8'd114; b_mant1 = 8'd135; b_mant2 = 8'd73; b_mant3 = 8'd135;
a_exp0 = 10'd388; a_exp1 = 10'd620; a_exp2 = 10'd662; a_exp3 = 10'd52;
b_exp0 = 10'd211; b_exp1 = 10'd356; b_exp2 = 10'd362; b_exp3 = 10'd179;
a_sign0 = 4'd16; a_sign1 = 4'd16; a_sign2 = 4'd12; a_sign3 = 4'd1;
b_sign0 = 4'd3; b_sign1 = 4'd5; b_sign2 = 4'd2; b_sign3 = 4'd6;
@(posedge clk_i);
a_mant0 = 8'd185; a_mant1 = 8'd0; a_mant2 = 8'd141; a_mant3 = 8'd109;
b_mant0 = 8'd229; b_mant1 = 8'd0; b_mant2 = 8'd153; b_mant3 = 8'd224;
a_exp0 = 10'd256; a_exp1 = 10'd318; a_exp2 = 10'd351; a_exp3 = 10'd673;
b_exp0 = 10'd515; b_exp1 = 10'd341; b_exp2 = 10'd64; b_exp3 = 10'd456;
a_sign0 = 4'd11; a_sign1 = 4'd1; a_sign2 = 4'd7; a_sign3 = 4'd7;
b_sign0 = 4'd3; b_sign1 = 4'd2; b_sign2 = 4'd8; b_sign3 = 4'd1;
@(posedge clk_i);
a_mant0 = 8'd5; a_mant1 = 8'd25; a_mant2 = 8'd149; a_mant3 = 8'd82;
b_mant0 = 8'd24; b_mant1 = 8'd85; b_mant2 = 8'd107; b_mant3 = 8'd200;
a_exp0 = 10'd506; a_exp1 = 10'd535; a_exp2 = 10'd414; a_exp3 = 10'd607;
b_exp0 = 10'd132; b_exp1 = 10'd932; b_exp2 = 10'd458; b_exp3 = 10'd797;
a_sign0 = 4'd11; a_sign1 = 4'd1; a_sign2 = 4'd9; a_sign3 = 4'd3;
b_sign0 = 4'd8; b_sign1 = 4'd4; b_sign2 = 4'd13; b_sign3 = 4'd9;
@(posedge clk_i);
a_mant0 = 8'd21; a_mant1 = 8'd119; a_mant2 = 8'd25; a_mant3 = 8'd45;
b_mant0 = 8'd86; b_mant1 = 8'd175; b_mant2 = 8'd110; b_mant3 = 8'd105;
a_exp0 = 10'd418; a_exp1 = 10'd115; a_exp2 = 10'd708; a_exp3 = 10'd69;
b_exp0 = 10'd587; b_exp1 = 10'd718; b_exp2 = 10'd246; b_exp3 = 10'd322;
a_sign0 = 4'd0; a_sign1 = 4'd5; a_sign2 = 4'd4; a_sign3 = 4'd9;
b_sign0 = 4'd15; b_sign1 = 4'd10; b_sign2 = 4'd2; b_sign3 = 4'd10;
@(posedge clk_i);
a_mant0 = 8'd181; a_mant1 = 8'd224; a_mant2 = 8'd165; a_mant3 = 8'd246;
b_mant0 = 8'd9; b_mant1 = 8'd201; b_mant2 = 8'd47; b_mant3 = 8'd88;
a_exp0 = 10'd989; a_exp1 = 10'd145; a_exp2 = 10'd480; a_exp3 = 10'd635;
b_exp0 = 10'd725; b_exp1 = 10'd975; b_exp2 = 10'd630; b_exp3 = 10'd940;
a_sign0 = 4'd10; a_sign1 = 4'd13; a_sign2 = 4'd13; a_sign3 = 4'd16;
b_sign0 = 4'd13; b_sign1 = 4'd9; b_sign2 = 4'd7; b_sign3 = 4'd11;
@(posedge clk_i);
a_mant0 = 8'd187; a_mant1 = 8'd223; a_mant2 = 8'd178; a_mant3 = 8'd208;
b_mant0 = 8'd146; b_mant1 = 8'd77; b_mant2 = 8'd198; b_mant3 = 8'd54;
a_exp0 = 10'd752; a_exp1 = 10'd565; a_exp2 = 10'd1016; a_exp3 = 10'd400;
b_exp0 = 10'd330; b_exp1 = 10'd122; b_exp2 = 10'd309; b_exp3 = 10'd799;
a_sign0 = 4'd8; a_sign1 = 4'd4; a_sign2 = 4'd15; a_sign3 = 4'd8;
b_sign0 = 4'd3; b_sign1 = 4'd5; b_sign2 = 4'd13; b_sign3 = 4'd9;
@(posedge clk_i);
a_mant0 = 8'd153; a_mant1 = 8'd91; a_mant2 = 8'd42; a_mant3 = 8'd109;
b_mant0 = 8'd23; b_mant1 = 8'd120; b_mant2 = 8'd78; b_mant3 = 8'd64;
a_exp0 = 10'd21; a_exp1 = 10'd93; a_exp2 = 10'd435; a_exp3 = 10'd517;
b_exp0 = 10'd367; b_exp1 = 10'd381; b_exp2 = 10'd88; b_exp3 = 10'd230;
a_sign0 = 4'd12; a_sign1 = 4'd6; a_sign2 = 4'd12; a_sign3 = 4'd8;
b_sign0 = 4'd0; b_sign1 = 4'd12; b_sign2 = 4'd5; b_sign3 = 4'd16;
@(posedge clk_i);
a_mant0 = 8'd69; a_mant1 = 8'd137; a_mant2 = 8'd235; a_mant3 = 8'd70;
b_mant0 = 8'd239; b_mant1 = 8'd112; b_mant2 = 8'd115; b_mant3 = 8'd204;
a_exp0 = 10'd636; a_exp1 = 10'd397; a_exp2 = 10'd304; a_exp3 = 10'd14;
b_exp0 = 10'd956; b_exp1 = 10'd156; b_exp2 = 10'd564; b_exp3 = 10'd197;
a_sign0 = 4'd2; a_sign1 = 4'd12; a_sign2 = 4'd4; a_sign3 = 4'd4;
b_sign0 = 4'd5; b_sign1 = 4'd2; b_sign2 = 4'd7; b_sign3 = 4'd5;
@(posedge clk_i);
shared_exps0 = 8'd108;
shared_exps1 = 8'd131;
a_mant0 = 8'd83; a_mant1 = 8'd158; a_mant2 = 8'd190; a_mant3 = 8'd172;
b_mant0 = 8'd246; b_mant1 = 8'd215; b_mant2 = 8'd88; b_mant3 = 8'd96;
a_exp0 = 10'd296; a_exp1 = 10'd866; a_exp2 = 10'd588; a_exp3 = 10'd7;
b_exp0 = 10'd887; b_exp1 = 10'd957; b_exp2 = 10'd183; b_exp3 = 10'd283;
a_sign0 = 4'd4; a_sign1 = 4'd12; a_sign2 = 4'd6; a_sign3 = 4'd13;
b_sign0 = 4'd6; b_sign1 = 4'd1; b_sign2 = 4'd5; b_sign3 = 4'd10;
@(posedge clk_i);
a_mant0 = 8'd49; a_mant1 = 8'd227; a_mant2 = 8'd135; a_mant3 = 8'd68;
b_mant0 = 8'd210; b_mant1 = 8'd180; b_mant2 = 8'd112; b_mant3 = 8'd182;
a_exp0 = 10'd753; a_exp1 = 10'd365; a_exp2 = 10'd299; a_exp3 = 10'd96;
b_exp0 = 10'd467; b_exp1 = 10'd1003; b_exp2 = 10'd977; b_exp3 = 10'd149;
a_sign0 = 4'd6; a_sign1 = 4'd11; a_sign2 = 4'd5; a_sign3 = 4'd10;
b_sign0 = 4'd12; b_sign1 = 4'd10; b_sign2 = 4'd5; b_sign3 = 4'd10;
@(posedge clk_i);
a_mant0 = 8'd217; a_mant1 = 8'd31; a_mant2 = 8'd244; a_mant3 = 8'd123;
b_mant0 = 8'd229; b_mant1 = 8'd213; b_mant2 = 8'd242; b_mant3 = 8'd247;
a_exp0 = 10'd2; a_exp1 = 10'd690; a_exp2 = 10'd373; a_exp3 = 10'd952;
b_exp0 = 10'd912; b_exp1 = 10'd700; b_exp2 = 10'd590; b_exp3 = 10'd852;
a_sign0 = 4'd0; a_sign1 = 4'd8; a_sign2 = 4'd4; a_sign3 = 4'd10;
b_sign0 = 4'd13; b_sign1 = 4'd7; b_sign2 = 4'd14; b_sign3 = 4'd0;
@(posedge clk_i);
a_mant0 = 8'd174; a_mant1 = 8'd73; a_mant2 = 8'd119; a_mant3 = 8'd247;
b_mant0 = 8'd189; b_mant1 = 8'd106; b_mant2 = 8'd125; b_mant3 = 8'd141;
a_exp0 = 10'd326; a_exp1 = 10'd980; a_exp2 = 10'd165; a_exp3 = 10'd914;
b_exp0 = 10'd327; b_exp1 = 10'd327; b_exp2 = 10'd378; b_exp3 = 10'd474;
a_sign0 = 4'd16; a_sign1 = 4'd10; a_sign2 = 4'd15; a_sign3 = 4'd0;
b_sign0 = 4'd0; b_sign1 = 4'd12; b_sign2 = 4'd1; b_sign3 = 4'd10;
@(posedge clk_i);
a_mant0 = 8'd27; a_mant1 = 8'd53; a_mant2 = 8'd179; a_mant3 = 8'd76;
b_mant0 = 8'd9; b_mant1 = 8'd156; b_mant2 = 8'd191; b_mant3 = 8'd237;
a_exp0 = 10'd51; a_exp1 = 10'd615; a_exp2 = 10'd466; a_exp3 = 10'd844;
b_exp0 = 10'd341; b_exp1 = 10'd751; b_exp2 = 10'd422; b_exp3 = 10'd480;
a_sign0 = 4'd5; a_sign1 = 4'd0; a_sign2 = 4'd7; a_sign3 = 4'd6;
b_sign0 = 4'd1; b_sign1 = 4'd7; b_sign2 = 4'd5; b_sign3 = 4'd9;
@(posedge clk_i);
a_mant0 = 8'd231; a_mant1 = 8'd60; a_mant2 = 8'd200; a_mant3 = 8'd19;
b_mant0 = 8'd57; b_mant1 = 8'd59; b_mant2 = 8'd254; b_mant3 = 8'd126;
a_exp0 = 10'd496; a_exp1 = 10'd302; a_exp2 = 10'd184; a_exp3 = 10'd571;
b_exp0 = 10'd662; b_exp1 = 10'd279; b_exp2 = 10'd84; b_exp3 = 10'd56;
a_sign0 = 4'd2; a_sign1 = 4'd12; a_sign2 = 4'd13; a_sign3 = 4'd14;
b_sign0 = 4'd6; b_sign1 = 4'd6; b_sign2 = 4'd9; b_sign3 = 4'd5;
@(posedge clk_i);
a_mant0 = 8'd76; a_mant1 = 8'd252; a_mant2 = 8'd86; a_mant3 = 8'd136;
b_mant0 = 8'd97; b_mant1 = 8'd234; b_mant2 = 8'd224; b_mant3 = 8'd14;
a_exp0 = 10'd613; a_exp1 = 10'd340; a_exp2 = 10'd251; a_exp3 = 10'd476;
b_exp0 = 10'd874; b_exp1 = 10'd243; b_exp2 = 10'd815; b_exp3 = 10'd742;
a_sign0 = 4'd13; a_sign1 = 4'd10; a_sign2 = 4'd15; a_sign3 = 4'd14;
b_sign0 = 4'd4; b_sign1 = 4'd15; b_sign2 = 4'd0; b_sign3 = 4'd6;
@(posedge clk_i);
a_mant0 = 8'd72; a_mant1 = 8'd146; a_mant2 = 8'd251; a_mant3 = 8'd93;
b_mant0 = 8'd58; b_mant1 = 8'd85; b_mant2 = 8'd120; b_mant3 = 8'd224;
a_exp0 = 10'd484; a_exp1 = 10'd218; a_exp2 = 10'd739; a_exp3 = 10'd159;
b_exp0 = 10'd49; b_exp1 = 10'd553; b_exp2 = 10'd207; b_exp3 = 10'd232;
a_sign0 = 4'd13; a_sign1 = 4'd15; a_sign2 = 4'd16; a_sign3 = 4'd7;
b_sign0 = 4'd15; b_sign1 = 4'd5; b_sign2 = 4'd9; b_sign3 = 4'd4;
@(posedge clk_i);
shared_exps0 = 8'd119;
shared_exps1 = 8'd127;
a_mant0 = 8'd193; a_mant1 = 8'd43; a_mant2 = 8'd152; a_mant3 = 8'd131;
b_mant0 = 8'd132; b_mant1 = 8'd80; b_mant2 = 8'd189; b_mant3 = 8'd111;
a_exp0 = 10'd616; a_exp1 = 10'd270; a_exp2 = 10'd933; a_exp3 = 10'd227;
b_exp0 = 10'd433; b_exp1 = 10'd815; b_exp2 = 10'd218; b_exp3 = 10'd164;
a_sign0 = 4'd12; a_sign1 = 4'd14; a_sign2 = 4'd16; a_sign3 = 4'd4;
b_sign0 = 4'd4; b_sign1 = 4'd11; b_sign2 = 4'd11; b_sign3 = 4'd5;
@(posedge clk_i);
a_mant0 = 8'd162; a_mant1 = 8'd197; a_mant2 = 8'd27; a_mant3 = 8'd213;
b_mant0 = 8'd48; b_mant1 = 8'd30; b_mant2 = 8'd9; b_mant3 = 8'd177;
a_exp0 = 10'd249; a_exp1 = 10'd762; a_exp2 = 10'd835; a_exp3 = 10'd693;
b_exp0 = 10'd432; b_exp1 = 10'd764; b_exp2 = 10'd942; b_exp3 = 10'd104;
a_sign0 = 4'd8; a_sign1 = 4'd7; a_sign2 = 4'd16; a_sign3 = 4'd1;
b_sign0 = 4'd5; b_sign1 = 4'd6; b_sign2 = 4'd13; b_sign3 = 4'd16;
@(posedge clk_i);
a_mant0 = 8'd170; a_mant1 = 8'd10; a_mant2 = 8'd94; a_mant3 = 8'd156;
b_mant0 = 8'd160; b_mant1 = 8'd197; b_mant2 = 8'd235; b_mant3 = 8'd80;
a_exp0 = 10'd251; a_exp1 = 10'd210; a_exp2 = 10'd532; a_exp3 = 10'd255;
b_exp0 = 10'd506; b_exp1 = 10'd498; b_exp2 = 10'd88; b_exp3 = 10'd230;
a_sign0 = 4'd15; a_sign1 = 4'd6; a_sign2 = 4'd5; a_sign3 = 4'd3;
b_sign0 = 4'd5; b_sign1 = 4'd4; b_sign2 = 4'd11; b_sign3 = 4'd8;
@(posedge clk_i);
a_mant0 = 8'd189; a_mant1 = 8'd109; a_mant2 = 8'd254; a_mant3 = 8'd50;
b_mant0 = 8'd191; b_mant1 = 8'd119; b_mant2 = 8'd89; b_mant3 = 8'd230;
a_exp0 = 10'd323; a_exp1 = 10'd302; a_exp2 = 10'd227; a_exp3 = 10'd893;
b_exp0 = 10'd497; b_exp1 = 10'd32; b_exp2 = 10'd263; b_exp3 = 10'd1019;
a_sign0 = 4'd2; a_sign1 = 4'd6; a_sign2 = 4'd14; a_sign3 = 4'd11;
b_sign0 = 4'd11; b_sign1 = 4'd1; b_sign2 = 4'd11; b_sign3 = 4'd14;
@(posedge clk_i);
a_mant0 = 8'd67; a_mant1 = 8'd145; a_mant2 = 8'd118; a_mant3 = 8'd69;
b_mant0 = 8'd56; b_mant1 = 8'd100; b_mant2 = 8'd52; b_mant3 = 8'd191;
a_exp0 = 10'd887; a_exp1 = 10'd263; a_exp2 = 10'd540; a_exp3 = 10'd319;
b_exp0 = 10'd525; b_exp1 = 10'd754; b_exp2 = 10'd326; b_exp3 = 10'd766;
a_sign0 = 4'd15; a_sign1 = 4'd12; a_sign2 = 4'd10; a_sign3 = 4'd6;
b_sign0 = 4'd12; b_sign1 = 4'd11; b_sign2 = 4'd3; b_sign3 = 4'd9;
@(posedge clk_i);
a_mant0 = 8'd147; a_mant1 = 8'd149; a_mant2 = 8'd57; a_mant3 = 8'd150;
b_mant0 = 8'd236; b_mant1 = 8'd30; b_mant2 = 8'd153; b_mant3 = 8'd208;
a_exp0 = 10'd958; a_exp1 = 10'd540; a_exp2 = 10'd348; a_exp3 = 10'd563;
b_exp0 = 10'd972; b_exp1 = 10'd342; b_exp2 = 10'd823; b_exp3 = 10'd290;
a_sign0 = 4'd15; a_sign1 = 4'd14; a_sign2 = 4'd4; a_sign3 = 4'd4;
b_sign0 = 4'd12; b_sign1 = 4'd13; b_sign2 = 4'd7; b_sign3 = 4'd7;
@(posedge clk_i);
a_mant0 = 8'd191; a_mant1 = 8'd107; a_mant2 = 8'd26; a_mant3 = 8'd199;
b_mant0 = 8'd174; b_mant1 = 8'd133; b_mant2 = 8'd221; b_mant3 = 8'd42;
a_exp0 = 10'd243; a_exp1 = 10'd1015; a_exp2 = 10'd885; a_exp3 = 10'd716;
b_exp0 = 10'd782; b_exp1 = 10'd336; b_exp2 = 10'd728; b_exp3 = 10'd415;
a_sign0 = 4'd2; a_sign1 = 4'd14; a_sign2 = 4'd12; a_sign3 = 4'd13;
b_sign0 = 4'd15; b_sign1 = 4'd11; b_sign2 = 4'd12; b_sign3 = 4'd5;
@(posedge clk_i);
a_mant0 = 8'd189; a_mant1 = 8'd85; a_mant2 = 8'd66; a_mant3 = 8'd1;
b_mant0 = 8'd128; b_mant1 = 8'd178; b_mant2 = 8'd97; b_mant3 = 8'd42;
a_exp0 = 10'd696; a_exp1 = 10'd128; a_exp2 = 10'd59; a_exp3 = 10'd151;
b_exp0 = 10'd940; b_exp1 = 10'd914; b_exp2 = 10'd370; b_exp3 = 10'd176;
a_sign0 = 4'd7; a_sign1 = 4'd11; a_sign2 = 4'd16; a_sign3 = 4'd3;
b_sign0 = 4'd12; b_sign1 = 4'd8; b_sign2 = 4'd5; b_sign3 = 4'd11;
@(posedge clk_i);
shared_exps0 = 8'd123;
shared_exps1 = 8'd129;
rstn = 0;
@(posedge clk_i);
rstn = 1;
a_mant0 = 8'd218; a_mant1 = 8'd74; a_mant2 = 8'd232; a_mant3 = 8'd87;
b_mant0 = 8'd114; b_mant1 = 8'd115; b_mant2 = 8'd215; b_mant3 = 8'd74;
a_exp0 = 10'd144; a_exp1 = 10'd817; a_exp2 = 10'd21; a_exp3 = 10'd12;
b_exp0 = 10'd890; b_exp1 = 10'd198; b_exp2 = 10'd545; b_exp3 = 10'd911;
a_sign0 = 4'd16; a_sign1 = 4'd9; a_sign2 = 4'd9; a_sign3 = 4'd11;
b_sign0 = 4'd3; b_sign1 = 4'd1; b_sign2 = 4'd2; b_sign3 = 4'd14;
@(posedge clk_i);
a_mant0 = 8'd96; a_mant1 = 8'd223; a_mant2 = 8'd53; a_mant3 = 8'd242;
b_mant0 = 8'd217; b_mant1 = 8'd182; b_mant2 = 8'd138; b_mant3 = 8'd209;
a_exp0 = 10'd127; a_exp1 = 10'd58; a_exp2 = 10'd786; a_exp3 = 10'd799;
b_exp0 = 10'd911; b_exp1 = 10'd408; b_exp2 = 10'd739; b_exp3 = 10'd687;
a_sign0 = 4'd3; a_sign1 = 4'd4; a_sign2 = 4'd2; a_sign3 = 4'd12;
b_sign0 = 4'd14; b_sign1 = 4'd12; b_sign2 = 4'd1; b_sign3 = 4'd10;
@(posedge clk_i);
a_mant0 = 8'd190; a_mant1 = 8'd50; a_mant2 = 8'd142; a_mant3 = 8'd89;
b_mant0 = 8'd132; b_mant1 = 8'd64; b_mant2 = 8'd13; b_mant3 = 8'd166;
a_exp0 = 10'd634; a_exp1 = 10'd161; a_exp2 = 10'd284; a_exp3 = 10'd402;
b_exp0 = 10'd862; b_exp1 = 10'd994; b_exp2 = 10'd466; b_exp3 = 10'd777;
a_sign0 = 4'd12; a_sign1 = 4'd12; a_sign2 = 4'd12; a_sign3 = 4'd14;
b_sign0 = 4'd3; b_sign1 = 4'd13; b_sign2 = 4'd7; b_sign3 = 4'd16;
@(posedge clk_i);
a_mant0 = 8'd13; a_mant1 = 8'd177; a_mant2 = 8'd42; a_mant3 = 8'd152;
b_mant0 = 8'd104; b_mant1 = 8'd199; b_mant2 = 8'd92; b_mant3 = 8'd136;
a_exp0 = 10'd259; a_exp1 = 10'd373; a_exp2 = 10'd1004; a_exp3 = 10'd269;
b_exp0 = 10'd105; b_exp1 = 10'd435; b_exp2 = 10'd382; b_exp3 = 10'd13;
a_sign0 = 4'd12; a_sign1 = 4'd3; a_sign2 = 4'd10; a_sign3 = 4'd0;
b_sign0 = 4'd8; b_sign1 = 4'd9; b_sign2 = 4'd16; b_sign3 = 4'd8;
@(posedge clk_i);
a_mant0 = 8'd215; a_mant1 = 8'd195; a_mant2 = 8'd195; a_mant3 = 8'd238;
b_mant0 = 8'd201; b_mant1 = 8'd192; b_mant2 = 8'd92; b_mant3 = 8'd40;
a_exp0 = 10'd720; a_exp1 = 10'd774; a_exp2 = 10'd109; a_exp3 = 10'd959;
b_exp0 = 10'd676; b_exp1 = 10'd109; b_exp2 = 10'd504; b_exp3 = 10'd222;
a_sign0 = 4'd3; a_sign1 = 4'd9; a_sign2 = 4'd12; a_sign3 = 4'd16;
b_sign0 = 4'd10; b_sign1 = 4'd5; b_sign2 = 4'd10; b_sign3 = 4'd3;
@(posedge clk_i);
a_mant0 = 8'd6; a_mant1 = 8'd130; a_mant2 = 8'd111; a_mant3 = 8'd158;
b_mant0 = 8'd197; b_mant1 = 8'd10; b_mant2 = 8'd137; b_mant3 = 8'd189;
a_exp0 = 10'd332; a_exp1 = 10'd374; a_exp2 = 10'd931; a_exp3 = 10'd116;
b_exp0 = 10'd340; b_exp1 = 10'd203; b_exp2 = 10'd337; b_exp3 = 10'd892;
a_sign0 = 4'd2; a_sign1 = 4'd14; a_sign2 = 4'd0; a_sign3 = 4'd0;
b_sign0 = 4'd5; b_sign1 = 4'd10; b_sign2 = 4'd16; b_sign3 = 4'd1;
@(posedge clk_i);
a_mant0 = 8'd214; a_mant1 = 8'd205; a_mant2 = 8'd165; a_mant3 = 8'd88;
b_mant0 = 8'd236; b_mant1 = 8'd141; b_mant2 = 8'd35; b_mant3 = 8'd200;
a_exp0 = 10'd59; a_exp1 = 10'd825; a_exp2 = 10'd1004; a_exp3 = 10'd909;
b_exp0 = 10'd617; b_exp1 = 10'd980; b_exp2 = 10'd24; b_exp3 = 10'd288;
a_sign0 = 4'd8; a_sign1 = 4'd11; a_sign2 = 4'd0; a_sign3 = 4'd2;
b_sign0 = 4'd10; b_sign1 = 4'd16; b_sign2 = 4'd10; b_sign3 = 4'd13;
@(posedge clk_i);
shared_exps0 = 8'd131;
shared_exps1 = 8'd126;
a_mant0 = 8'd21; a_mant1 = 8'd70; a_mant2 = 8'd50; a_mant3 = 8'd75;
b_mant0 = 8'd76; b_mant1 = 8'd116; b_mant2 = 8'd10; b_mant3 = 8'd68;
a_exp0 = 10'd877; a_exp1 = 10'd219; a_exp2 = 10'd695; a_exp3 = 10'd578;
b_exp0 = 10'd806; b_exp1 = 10'd82; b_exp2 = 10'd158; b_exp3 = 10'd446;
a_sign0 = 4'd11; a_sign1 = 4'd4; a_sign2 = 4'd0; a_sign3 = 4'd10;
b_sign0 = 4'd1; b_sign1 = 4'd3; b_sign2 = 4'd14; b_sign3 = 4'd10;
@(posedge clk_i);
a_mant0 = 8'd48; a_mant1 = 8'd199; a_mant2 = 8'd108; a_mant3 = 8'd251;
b_mant0 = 8'd241; b_mant1 = 8'd68; b_mant2 = 8'd18; b_mant3 = 8'd84;
a_exp0 = 10'd836; a_exp1 = 10'd878; a_exp2 = 10'd74; a_exp3 = 10'd194;
b_exp0 = 10'd522; b_exp1 = 10'd537; b_exp2 = 10'd795; b_exp3 = 10'd780;
a_sign0 = 4'd10; a_sign1 = 4'd16; a_sign2 = 4'd7; a_sign3 = 4'd2;
b_sign0 = 4'd0; b_sign1 = 4'd12; b_sign2 = 4'd9; b_sign3 = 4'd2;
@(posedge clk_i);
a_mant0 = 8'd73; a_mant1 = 8'd189; a_mant2 = 8'd10; a_mant3 = 8'd228;
b_mant0 = 8'd221; b_mant1 = 8'd138; b_mant2 = 8'd203; b_mant3 = 8'd244;
a_exp0 = 10'd909; a_exp1 = 10'd640; a_exp2 = 10'd788; a_exp3 = 10'd241;
b_exp0 = 10'd401; b_exp1 = 10'd859; b_exp2 = 10'd87; b_exp3 = 10'd946;
a_sign0 = 4'd8; a_sign1 = 4'd13; a_sign2 = 4'd15; a_sign3 = 4'd8;
b_sign0 = 4'd5; b_sign1 = 4'd0; b_sign2 = 4'd16; b_sign3 = 4'd7;
@(posedge clk_i);
a_mant0 = 8'd137; a_mant1 = 8'd102; a_mant2 = 8'd212; a_mant3 = 8'd66;
b_mant0 = 8'd115; b_mant1 = 8'd117; b_mant2 = 8'd65; b_mant3 = 8'd57;
a_exp0 = 10'd122; a_exp1 = 10'd372; a_exp2 = 10'd1020; a_exp3 = 10'd733;
b_exp0 = 10'd877; b_exp1 = 10'd710; b_exp2 = 10'd662; b_exp3 = 10'd273;
a_sign0 = 4'd11; a_sign1 = 4'd11; a_sign2 = 4'd12; a_sign3 = 4'd15;
b_sign0 = 4'd4; b_sign1 = 4'd11; b_sign2 = 4'd11; b_sign3 = 4'd1;
@(posedge clk_i);
a_mant0 = 8'd135; a_mant1 = 8'd34; a_mant2 = 8'd99; a_mant3 = 8'd199;
b_mant0 = 8'd157; b_mant1 = 8'd111; b_mant2 = 8'd40; b_mant3 = 8'd165;
a_exp0 = 10'd62; a_exp1 = 10'd562; a_exp2 = 10'd998; a_exp3 = 10'd520;
b_exp0 = 10'd249; b_exp1 = 10'd98; b_exp2 = 10'd121; b_exp3 = 10'd961;
a_sign0 = 4'd12; a_sign1 = 4'd12; a_sign2 = 4'd6; a_sign3 = 4'd2;
b_sign0 = 4'd12; b_sign1 = 4'd9; b_sign2 = 4'd12; b_sign3 = 4'd16;
@(posedge clk_i);
a_mant0 = 8'd180; a_mant1 = 8'd139; a_mant2 = 8'd34; a_mant3 = 8'd65;
b_mant0 = 8'd238; b_mant1 = 8'd96; b_mant2 = 8'd105; b_mant3 = 8'd43;
a_exp0 = 10'd466; a_exp1 = 10'd863; a_exp2 = 10'd915; a_exp3 = 10'd787;
b_exp0 = 10'd181; b_exp1 = 10'd9; b_exp2 = 10'd801; b_exp3 = 10'd161;
a_sign0 = 4'd8; a_sign1 = 4'd14; a_sign2 = 4'd10; a_sign3 = 4'd8;
b_sign0 = 4'd13; b_sign1 = 4'd6; b_sign2 = 4'd12; b_sign3 = 4'd5;
@(posedge clk_i);
a_mant0 = 8'd104; a_mant1 = 8'd47; a_mant2 = 8'd148; a_mant3 = 8'd44;
b_mant0 = 8'd8; b_mant1 = 8'd123; b_mant2 = 8'd105; b_mant3 = 8'd106;
a_exp0 = 10'd1006; a_exp1 = 10'd441; a_exp2 = 10'd959; a_exp3 = 10'd815;
b_exp0 = 10'd1003; b_exp1 = 10'd904; b_exp2 = 10'd973; b_exp3 = 10'd751;
a_sign0 = 4'd14; a_sign1 = 4'd16; a_sign2 = 4'd16; a_sign3 = 4'd12;
b_sign0 = 4'd15; b_sign1 = 4'd12; b_sign2 = 4'd8; b_sign3 = 4'd0;
@(posedge clk_i);
a_mant0 = 8'd62; a_mant1 = 8'd68; a_mant2 = 8'd62; a_mant3 = 8'd226;
b_mant0 = 8'd249; b_mant1 = 8'd173; b_mant2 = 8'd197; b_mant3 = 8'd188;
a_exp0 = 10'd189; a_exp1 = 10'd656; a_exp2 = 10'd619; a_exp3 = 10'd135;
b_exp0 = 10'd535; b_exp1 = 10'd372; b_exp2 = 10'd831; b_exp3 = 10'd967;
a_sign0 = 4'd8; a_sign1 = 4'd1; a_sign2 = 4'd3; a_sign3 = 4'd10;
b_sign0 = 4'd3; b_sign1 = 4'd2; b_sign2 = 4'd7; b_sign3 = 4'd4;
@(posedge clk_i);
shared_exps0 = 8'd145;
shared_exps1 = 8'd117;
a_mant0 = 8'd181; a_mant1 = 8'd142; a_mant2 = 8'd142; a_mant3 = 8'd47;
b_mant0 = 8'd174; b_mant1 = 8'd162; b_mant2 = 8'd172; b_mant3 = 8'd65;
a_exp0 = 10'd3; a_exp1 = 10'd425; a_exp2 = 10'd507; a_exp3 = 10'd963;
b_exp0 = 10'd649; b_exp1 = 10'd763; b_exp2 = 10'd263; b_exp3 = 10'd725;
a_sign0 = 4'd15; a_sign1 = 4'd0; a_sign2 = 4'd4; a_sign3 = 4'd6;
b_sign0 = 4'd0; b_sign1 = 4'd8; b_sign2 = 4'd16; b_sign3 = 4'd11;
@(posedge clk_i);
a_mant0 = 8'd23; a_mant1 = 8'd201; a_mant2 = 8'd8; a_mant3 = 8'd199;
b_mant0 = 8'd64; b_mant1 = 8'd67; b_mant2 = 8'd238; b_mant3 = 8'd234;
a_exp0 = 10'd397; a_exp1 = 10'd666; a_exp2 = 10'd504; a_exp3 = 10'd477;
b_exp0 = 10'd716; b_exp1 = 10'd810; b_exp2 = 10'd603; b_exp3 = 10'd648;
a_sign0 = 4'd2; a_sign1 = 4'd3; a_sign2 = 4'd11; a_sign3 = 4'd16;
b_sign0 = 4'd3; b_sign1 = 4'd4; b_sign2 = 4'd10; b_sign3 = 4'd15;
@(posedge clk_i);
a_mant0 = 8'd90; a_mant1 = 8'd8; a_mant2 = 8'd205; a_mant3 = 8'd230;
b_mant0 = 8'd253; b_mant1 = 8'd248; b_mant2 = 8'd158; b_mant3 = 8'd212;
a_exp0 = 10'd969; a_exp1 = 10'd565; a_exp2 = 10'd732; a_exp3 = 10'd200;
b_exp0 = 10'd933; b_exp1 = 10'd509; b_exp2 = 10'd166; b_exp3 = 10'd859;
a_sign0 = 4'd12; a_sign1 = 4'd13; a_sign2 = 4'd0; a_sign3 = 4'd12;
b_sign0 = 4'd16; b_sign1 = 4'd6; b_sign2 = 4'd0; b_sign3 = 4'd4;
@(posedge clk_i);
a_mant0 = 8'd21; a_mant1 = 8'd55; a_mant2 = 8'd90; a_mant3 = 8'd190;
b_mant0 = 8'd246; b_mant1 = 8'd47; b_mant2 = 8'd22; b_mant3 = 8'd81;
a_exp0 = 10'd609; a_exp1 = 10'd819; a_exp2 = 10'd579; a_exp3 = 10'd193;
b_exp0 = 10'd885; b_exp1 = 10'd850; b_exp2 = 10'd654; b_exp3 = 10'd148;
a_sign0 = 4'd2; a_sign1 = 4'd3; a_sign2 = 4'd9; a_sign3 = 4'd11;
b_sign0 = 4'd15; b_sign1 = 4'd5; b_sign2 = 4'd6; b_sign3 = 4'd3;
@(posedge clk_i);
a_mant0 = 8'd140; a_mant1 = 8'd203; a_mant2 = 8'd65; a_mant3 = 8'd180;
b_mant0 = 8'd255; b_mant1 = 8'd240; b_mant2 = 8'd30; b_mant3 = 8'd233;
a_exp0 = 10'd27; a_exp1 = 10'd586; a_exp2 = 10'd338; a_exp3 = 10'd511;
b_exp0 = 10'd979; b_exp1 = 10'd170; b_exp2 = 10'd999; b_exp3 = 10'd550;
a_sign0 = 4'd0; a_sign1 = 4'd13; a_sign2 = 4'd7; a_sign3 = 4'd8;
b_sign0 = 4'd16; b_sign1 = 4'd13; b_sign2 = 4'd11; b_sign3 = 4'd5;
@(posedge clk_i);
a_mant0 = 8'd67; a_mant1 = 8'd154; a_mant2 = 8'd63; a_mant3 = 8'd119;
b_mant0 = 8'd221; b_mant1 = 8'd29; b_mant2 = 8'd84; b_mant3 = 8'd176;
a_exp0 = 10'd18; a_exp1 = 10'd711; a_exp2 = 10'd657; a_exp3 = 10'd605;
b_exp0 = 10'd158; b_exp1 = 10'd442; b_exp2 = 10'd116; b_exp3 = 10'd976;
a_sign0 = 4'd15; a_sign1 = 4'd2; a_sign2 = 4'd14; a_sign3 = 4'd8;
b_sign0 = 4'd12; b_sign1 = 4'd11; b_sign2 = 4'd5; b_sign3 = 4'd4;
@(posedge clk_i);
a_mant0 = 8'd27; a_mant1 = 8'd23; a_mant2 = 8'd196; a_mant3 = 8'd154;
b_mant0 = 8'd12; b_mant1 = 8'd0; b_mant2 = 8'd102; b_mant3 = 8'd45;
a_exp0 = 10'd76; a_exp1 = 10'd435; a_exp2 = 10'd222; a_exp3 = 10'd521;
b_exp0 = 10'd245; b_exp1 = 10'd300; b_exp2 = 10'd132; b_exp3 = 10'd573;
a_sign0 = 4'd10; a_sign1 = 4'd11; a_sign2 = 4'd15; a_sign3 = 4'd16;
b_sign0 = 4'd15; b_sign1 = 4'd7; b_sign2 = 4'd0; b_sign3 = 4'd12;
@(posedge clk_i);
a_mant0 = 8'd135; a_mant1 = 8'd35; a_mant2 = 8'd79; a_mant3 = 8'd109;
b_mant0 = 8'd224; b_mant1 = 8'd216; b_mant2 = 8'd231; b_mant3 = 8'd179;
a_exp0 = 10'd213; a_exp1 = 10'd896; a_exp2 = 10'd167; a_exp3 = 10'd907;
b_exp0 = 10'd1010; b_exp1 = 10'd367; b_exp2 = 10'd250; b_exp3 = 10'd720;
a_sign0 = 4'd3; a_sign1 = 4'd15; a_sign2 = 4'd0; a_sign3 = 4'd1;
b_sign0 = 4'd0; b_sign1 = 4'd3; b_sign2 = 4'd12; b_sign3 = 4'd15;
@(posedge clk_i);
shared_exps0 = 8'd119;
shared_exps1 = 8'd90;
a_mant0 = 8'd204; a_mant1 = 8'd107; a_mant2 = 8'd17; a_mant3 = 8'd113;
b_mant0 = 8'd232; b_mant1 = 8'd216; b_mant2 = 8'd162; b_mant3 = 8'd158;
a_exp0 = 10'd596; a_exp1 = 10'd205; a_exp2 = 10'd819; a_exp3 = 10'd882;
b_exp0 = 10'd457; b_exp1 = 10'd407; b_exp2 = 10'd810; b_exp3 = 10'd1015;
a_sign0 = 4'd15; a_sign1 = 4'd6; a_sign2 = 4'd0; a_sign3 = 4'd8;
b_sign0 = 4'd6; b_sign1 = 4'd8; b_sign2 = 4'd1; b_sign3 = 4'd7;
@(posedge clk_i);
a_mant0 = 8'd191; a_mant1 = 8'd75; a_mant2 = 8'd187; a_mant3 = 8'd24;
b_mant0 = 8'd80; b_mant1 = 8'd22; b_mant2 = 8'd23; b_mant3 = 8'd62;
a_exp0 = 10'd471; a_exp1 = 10'd409; a_exp2 = 10'd612; a_exp3 = 10'd859;
b_exp0 = 10'd731; b_exp1 = 10'd172; b_exp2 = 10'd312; b_exp3 = 10'd742;
a_sign0 = 4'd13; a_sign1 = 4'd13; a_sign2 = 4'd0; a_sign3 = 4'd4;
b_sign0 = 4'd0; b_sign1 = 4'd5; b_sign2 = 4'd0; b_sign3 = 4'd11;
@(posedge clk_i);
a_mant0 = 8'd221; a_mant1 = 8'd116; a_mant2 = 8'd231; a_mant3 = 8'd94;
b_mant0 = 8'd98; b_mant1 = 8'd217; b_mant2 = 8'd159; b_mant3 = 8'd122;
a_exp0 = 10'd709; a_exp1 = 10'd788; a_exp2 = 10'd31; a_exp3 = 10'd431;
b_exp0 = 10'd936; b_exp1 = 10'd28; b_exp2 = 10'd961; b_exp3 = 10'd536;
a_sign0 = 4'd13; a_sign1 = 4'd16; a_sign2 = 4'd15; a_sign3 = 4'd2;
b_sign0 = 4'd1; b_sign1 = 4'd14; b_sign2 = 4'd7; b_sign3 = 4'd8;
@(posedge clk_i);
a_mant0 = 8'd206; a_mant1 = 8'd153; a_mant2 = 8'd186; a_mant3 = 8'd141;
b_mant0 = 8'd196; b_mant1 = 8'd179; b_mant2 = 8'd22; b_mant3 = 8'd144;
a_exp0 = 10'd272; a_exp1 = 10'd445; a_exp2 = 10'd5; a_exp3 = 10'd592;
b_exp0 = 10'd470; b_exp1 = 10'd880; b_exp2 = 10'd566; b_exp3 = 10'd658;
a_sign0 = 4'd11; a_sign1 = 4'd5; a_sign2 = 4'd14; a_sign3 = 4'd5;
b_sign0 = 4'd16; b_sign1 = 4'd5; b_sign2 = 4'd6; b_sign3 = 4'd10;
@(posedge clk_i);
a_mant0 = 8'd191; a_mant1 = 8'd216; a_mant2 = 8'd109; a_mant3 = 8'd169;
b_mant0 = 8'd188; b_mant1 = 8'd130; b_mant2 = 8'd158; b_mant3 = 8'd49;
a_exp0 = 10'd982; a_exp1 = 10'd359; a_exp2 = 10'd860; a_exp3 = 10'd134;
b_exp0 = 10'd954; b_exp1 = 10'd49; b_exp2 = 10'd280; b_exp3 = 10'd698;
a_sign0 = 4'd6; a_sign1 = 4'd1; a_sign2 = 4'd10; a_sign3 = 4'd11;
b_sign0 = 4'd10; b_sign1 = 4'd2; b_sign2 = 4'd7; b_sign3 = 4'd7;
@(posedge clk_i);
a_mant0 = 8'd173; a_mant1 = 8'd171; a_mant2 = 8'd67; a_mant3 = 8'd209;
b_mant0 = 8'd207; b_mant1 = 8'd2; b_mant2 = 8'd61; b_mant3 = 8'd34;
a_exp0 = 10'd211; a_exp1 = 10'd753; a_exp2 = 10'd672; a_exp3 = 10'd529;
b_exp0 = 10'd963; b_exp1 = 10'd53; b_exp2 = 10'd984; b_exp3 = 10'd588;
a_sign0 = 4'd2; a_sign1 = 4'd5; a_sign2 = 4'd10; a_sign3 = 4'd16;
b_sign0 = 4'd13; b_sign1 = 4'd5; b_sign2 = 4'd12; b_sign3 = 4'd13;
@(posedge clk_i);
a_mant0 = 8'd238; a_mant1 = 8'd14; a_mant2 = 8'd252; a_mant3 = 8'd131;
b_mant0 = 8'd80; b_mant1 = 8'd31; b_mant2 = 8'd80; b_mant3 = 8'd165;
a_exp0 = 10'd960; a_exp1 = 10'd818; a_exp2 = 10'd682; a_exp3 = 10'd714;
b_exp0 = 10'd353; b_exp1 = 10'd189; b_exp2 = 10'd535; b_exp3 = 10'd434;
a_sign0 = 4'd11; a_sign1 = 4'd16; a_sign2 = 4'd0; a_sign3 = 4'd14;
b_sign0 = 4'd11; b_sign1 = 4'd12; b_sign2 = 4'd6; b_sign3 = 4'd1;
@(posedge clk_i);
a_mant0 = 8'd144; a_mant1 = 8'd96; a_mant2 = 8'd35; a_mant3 = 8'd77;
b_mant0 = 8'd38; b_mant1 = 8'd78; b_mant2 = 8'd107; b_mant3 = 8'd122;
a_exp0 = 10'd755; a_exp1 = 10'd191; a_exp2 = 10'd403; a_exp3 = 10'd345;
b_exp0 = 10'd574; b_exp1 = 10'd919; b_exp2 = 10'd11; b_exp3 = 10'd359;
a_sign0 = 4'd4; a_sign1 = 4'd13; a_sign2 = 4'd14; a_sign3 = 4'd6;
b_sign0 = 4'd2; b_sign1 = 4'd0; b_sign2 = 4'd4; b_sign3 = 4'd0;
@(posedge clk_i);
shared_exps0 = 8'd111;
shared_exps1 = 8'd124;
rstn = 0;
@(posedge clk_i);
rstn = 1;
a_mant0 = 8'd97; a_mant1 = 8'd71; a_mant2 = 8'd137; a_mant3 = 8'd146;
b_mant0 = 8'd202; b_mant1 = 8'd207; b_mant2 = 8'd240; b_mant3 = 8'd28;
a_exp0 = 10'd728; a_exp1 = 10'd681; a_exp2 = 10'd637; a_exp3 = 10'd41;
b_exp0 = 10'd781; b_exp1 = 10'd550; b_exp2 = 10'd42; b_exp3 = 10'd772;
a_sign0 = 4'd7; a_sign1 = 4'd8; a_sign2 = 4'd9; a_sign3 = 4'd7;
b_sign0 = 4'd16; b_sign1 = 4'd1; b_sign2 = 4'd7; b_sign3 = 4'd3;
@(posedge clk_i);
a_mant0 = 8'd124; a_mant1 = 8'd15; a_mant2 = 8'd143; a_mant3 = 8'd218;
b_mant0 = 8'd230; b_mant1 = 8'd3; b_mant2 = 8'd224; b_mant3 = 8'd234;
a_exp0 = 10'd117; a_exp1 = 10'd927; a_exp2 = 10'd72; a_exp3 = 10'd364;
b_exp0 = 10'd858; b_exp1 = 10'd687; b_exp2 = 10'd583; b_exp3 = 10'd750;
a_sign0 = 4'd16; a_sign1 = 4'd12; a_sign2 = 4'd5; a_sign3 = 4'd7;
b_sign0 = 4'd0; b_sign1 = 4'd2; b_sign2 = 4'd7; b_sign3 = 4'd4;
@(posedge clk_i);
a_mant0 = 8'd81; a_mant1 = 8'd28; a_mant2 = 8'd179; a_mant3 = 8'd250;
b_mant0 = 8'd36; b_mant1 = 8'd178; b_mant2 = 8'd118; b_mant3 = 8'd132;
a_exp0 = 10'd23; a_exp1 = 10'd968; a_exp2 = 10'd779; a_exp3 = 10'd790;
b_exp0 = 10'd574; b_exp1 = 10'd552; b_exp2 = 10'd480; b_exp3 = 10'd759;
a_sign0 = 4'd16; a_sign1 = 4'd0; a_sign2 = 4'd0; a_sign3 = 4'd7;
b_sign0 = 4'd14; b_sign1 = 4'd1; b_sign2 = 4'd16; b_sign3 = 4'd6;
@(posedge clk_i);
a_mant0 = 8'd26; a_mant1 = 8'd48; a_mant2 = 8'd108; a_mant3 = 8'd125;
b_mant0 = 8'd240; b_mant1 = 8'd153; b_mant2 = 8'd112; b_mant3 = 8'd252;
a_exp0 = 10'd447; a_exp1 = 10'd151; a_exp2 = 10'd697; a_exp3 = 10'd340;
b_exp0 = 10'd527; b_exp1 = 10'd886; b_exp2 = 10'd271; b_exp3 = 10'd274;
a_sign0 = 4'd8; a_sign1 = 4'd12; a_sign2 = 4'd5; a_sign3 = 4'd5;
b_sign0 = 4'd4; b_sign1 = 4'd9; b_sign2 = 4'd14; b_sign3 = 4'd3;
@(posedge clk_i);
a_mant0 = 8'd41; a_mant1 = 8'd27; a_mant2 = 8'd240; a_mant3 = 8'd235;
b_mant0 = 8'd62; b_mant1 = 8'd98; b_mant2 = 8'd189; b_mant3 = 8'd9;
a_exp0 = 10'd806; a_exp1 = 10'd748; a_exp2 = 10'd1009; a_exp3 = 10'd914;
b_exp0 = 10'd303; b_exp1 = 10'd759; b_exp2 = 10'd661; b_exp3 = 10'd267;
a_sign0 = 4'd0; a_sign1 = 4'd4; a_sign2 = 4'd5; a_sign3 = 4'd1;
b_sign0 = 4'd15; b_sign1 = 4'd1; b_sign2 = 4'd6; b_sign3 = 4'd0;
@(posedge clk_i);
a_mant0 = 8'd91; a_mant1 = 8'd92; a_mant2 = 8'd125; a_mant3 = 8'd30;
b_mant0 = 8'd83; b_mant1 = 8'd111; b_mant2 = 8'd85; b_mant3 = 8'd25;
a_exp0 = 10'd823; a_exp1 = 10'd662; a_exp2 = 10'd589; a_exp3 = 10'd518;
b_exp0 = 10'd834; b_exp1 = 10'd507; b_exp2 = 10'd99; b_exp3 = 10'd658;
a_sign0 = 4'd14; a_sign1 = 4'd10; a_sign2 = 4'd0; a_sign3 = 4'd14;
b_sign0 = 4'd6; b_sign1 = 4'd14; b_sign2 = 4'd2; b_sign3 = 4'd15;
@(posedge clk_i);
a_mant0 = 8'd64; a_mant1 = 8'd119; a_mant2 = 8'd243; a_mant3 = 8'd222;
b_mant0 = 8'd230; b_mant1 = 8'd9; b_mant2 = 8'd125; b_mant3 = 8'd165;
a_exp0 = 10'd612; a_exp1 = 10'd868; a_exp2 = 10'd501; a_exp3 = 10'd103;
b_exp0 = 10'd93; b_exp1 = 10'd338; b_exp2 = 10'd490; b_exp3 = 10'd540;
a_sign0 = 4'd9; a_sign1 = 4'd16; a_sign2 = 4'd15; a_sign3 = 4'd10;
b_sign0 = 4'd14; b_sign1 = 4'd16; b_sign2 = 4'd3; b_sign3 = 4'd5;
@(posedge clk_i);
shared_exps0 = 8'd132;
shared_exps1 = 8'd158;
a_mant0 = 8'd64; a_mant1 = 8'd223; a_mant2 = 8'd178; a_mant3 = 8'd45;
b_mant0 = 8'd180; b_mant1 = 8'd61; b_mant2 = 8'd48; b_mant3 = 8'd55;
a_exp0 = 10'd143; a_exp1 = 10'd97; a_exp2 = 10'd24; a_exp3 = 10'd1019;
b_exp0 = 10'd12; b_exp1 = 10'd974; b_exp2 = 10'd397; b_exp3 = 10'd452;
a_sign0 = 4'd7; a_sign1 = 4'd5; a_sign2 = 4'd0; a_sign3 = 4'd2;
b_sign0 = 4'd1; b_sign1 = 4'd16; b_sign2 = 4'd12; b_sign3 = 4'd14;
@(posedge clk_i);
a_mant0 = 8'd51; a_mant1 = 8'd240; a_mant2 = 8'd146; a_mant3 = 8'd34;
b_mant0 = 8'd108; b_mant1 = 8'd51; b_mant2 = 8'd22; b_mant3 = 8'd111;
a_exp0 = 10'd237; a_exp1 = 10'd721; a_exp2 = 10'd650; a_exp3 = 10'd590;
b_exp0 = 10'd819; b_exp1 = 10'd696; b_exp2 = 10'd778; b_exp3 = 10'd593;
a_sign0 = 4'd7; a_sign1 = 4'd12; a_sign2 = 4'd3; a_sign3 = 4'd4;
b_sign0 = 4'd8; b_sign1 = 4'd10; b_sign2 = 4'd6; b_sign3 = 4'd2;
@(posedge clk_i);
a_mant0 = 8'd77; a_mant1 = 8'd130; a_mant2 = 8'd212; a_mant3 = 8'd62;
b_mant0 = 8'd36; b_mant1 = 8'd6; b_mant2 = 8'd175; b_mant3 = 8'd250;
a_exp0 = 10'd747; a_exp1 = 10'd472; a_exp2 = 10'd288; a_exp3 = 10'd631;
b_exp0 = 10'd628; b_exp1 = 10'd7; b_exp2 = 10'd960; b_exp3 = 10'd324;
a_sign0 = 4'd3; a_sign1 = 4'd14; a_sign2 = 4'd15; a_sign3 = 4'd10;
b_sign0 = 4'd7; b_sign1 = 4'd12; b_sign2 = 4'd5; b_sign3 = 4'd8;
@(posedge clk_i);
a_mant0 = 8'd209; a_mant1 = 8'd162; a_mant2 = 8'd131; a_mant3 = 8'd227;
b_mant0 = 8'd76; b_mant1 = 8'd176; b_mant2 = 8'd65; b_mant3 = 8'd62;
a_exp0 = 10'd521; a_exp1 = 10'd888; a_exp2 = 10'd332; a_exp3 = 10'd92;
b_exp0 = 10'd473; b_exp1 = 10'd391; b_exp2 = 10'd549; b_exp3 = 10'd496;
a_sign0 = 4'd6; a_sign1 = 4'd6; a_sign2 = 4'd6; a_sign3 = 4'd10;
b_sign0 = 4'd16; b_sign1 = 4'd11; b_sign2 = 4'd12; b_sign3 = 4'd6;
@(posedge clk_i);
a_mant0 = 8'd112; a_mant1 = 8'd22; a_mant2 = 8'd32; a_mant3 = 8'd18;
b_mant0 = 8'd239; b_mant1 = 8'd184; b_mant2 = 8'd48; b_mant3 = 8'd2;
a_exp0 = 10'd486; a_exp1 = 10'd314; a_exp2 = 10'd582; a_exp3 = 10'd47;
b_exp0 = 10'd637; b_exp1 = 10'd602; b_exp2 = 10'd365; b_exp3 = 10'd930;
a_sign0 = 4'd16; a_sign1 = 4'd8; a_sign2 = 4'd15; a_sign3 = 4'd10;
b_sign0 = 4'd0; b_sign1 = 4'd2; b_sign2 = 4'd9; b_sign3 = 4'd8;
@(posedge clk_i);
a_mant0 = 8'd24; a_mant1 = 8'd188; a_mant2 = 8'd33; a_mant3 = 8'd139;
b_mant0 = 8'd98; b_mant1 = 8'd60; b_mant2 = 8'd223; b_mant3 = 8'd23;
a_exp0 = 10'd135; a_exp1 = 10'd780; a_exp2 = 10'd258; a_exp3 = 10'd160;
b_exp0 = 10'd242; b_exp1 = 10'd540; b_exp2 = 10'd119; b_exp3 = 10'd17;
a_sign0 = 4'd15; a_sign1 = 4'd14; a_sign2 = 4'd0; a_sign3 = 4'd0;
b_sign0 = 4'd1; b_sign1 = 4'd16; b_sign2 = 4'd11; b_sign3 = 4'd6;
@(posedge clk_i);
a_mant0 = 8'd162; a_mant1 = 8'd83; a_mant2 = 8'd172; a_mant3 = 8'd56;
b_mant0 = 8'd103; b_mant1 = 8'd118; b_mant2 = 8'd119; b_mant3 = 8'd63;
a_exp0 = 10'd604; a_exp1 = 10'd541; a_exp2 = 10'd353; a_exp3 = 10'd340;
b_exp0 = 10'd40; b_exp1 = 10'd562; b_exp2 = 10'd571; b_exp3 = 10'd664;
a_sign0 = 4'd15; a_sign1 = 4'd14; a_sign2 = 4'd14; a_sign3 = 4'd14;
b_sign0 = 4'd0; b_sign1 = 4'd2; b_sign2 = 4'd7; b_sign3 = 4'd7;
@(posedge clk_i);
a_mant0 = 8'd146; a_mant1 = 8'd84; a_mant2 = 8'd37; a_mant3 = 8'd179;
b_mant0 = 8'd173; b_mant1 = 8'd98; b_mant2 = 8'd219; b_mant3 = 8'd32;
a_exp0 = 10'd94; a_exp1 = 10'd799; a_exp2 = 10'd724; a_exp3 = 10'd369;
b_exp0 = 10'd117; b_exp1 = 10'd1003; b_exp2 = 10'd309; b_exp3 = 10'd592;
a_sign0 = 4'd7; a_sign1 = 4'd6; a_sign2 = 4'd16; a_sign3 = 4'd1;
b_sign0 = 4'd1; b_sign1 = 4'd3; b_sign2 = 4'd15; b_sign3 = 4'd8;
@(posedge clk_i);
shared_exps0 = 8'd147;
shared_exps1 = 8'd138;
a_mant0 = 8'd17; a_mant1 = 8'd132; a_mant2 = 8'd178; a_mant3 = 8'd32;
b_mant0 = 8'd210; b_mant1 = 8'd122; b_mant2 = 8'd200; b_mant3 = 8'd49;
a_exp0 = 10'd199; a_exp1 = 10'd385; a_exp2 = 10'd971; a_exp3 = 10'd885;
b_exp0 = 10'd10; b_exp1 = 10'd874; b_exp2 = 10'd904; b_exp3 = 10'd745;
a_sign0 = 4'd9; a_sign1 = 4'd0; a_sign2 = 4'd9; a_sign3 = 4'd13;
b_sign0 = 4'd4; b_sign1 = 4'd2; b_sign2 = 4'd10; b_sign3 = 4'd11;
@(posedge clk_i);
a_mant0 = 8'd131; a_mant1 = 8'd241; a_mant2 = 8'd93; a_mant3 = 8'd196;
b_mant0 = 8'd201; b_mant1 = 8'd144; b_mant2 = 8'd165; b_mant3 = 8'd206;
a_exp0 = 10'd518; a_exp1 = 10'd135; a_exp2 = 10'd985; a_exp3 = 10'd578;
b_exp0 = 10'd683; b_exp1 = 10'd445; b_exp2 = 10'd193; b_exp3 = 10'd867;
a_sign0 = 4'd0; a_sign1 = 4'd8; a_sign2 = 4'd5; a_sign3 = 4'd7;
b_sign0 = 4'd0; b_sign1 = 4'd11; b_sign2 = 4'd1; b_sign3 = 4'd0;
@(posedge clk_i);
a_mant0 = 8'd171; a_mant1 = 8'd236; a_mant2 = 8'd209; a_mant3 = 8'd37;
b_mant0 = 8'd95; b_mant1 = 8'd238; b_mant2 = 8'd14; b_mant3 = 8'd9;
a_exp0 = 10'd977; a_exp1 = 10'd435; a_exp2 = 10'd925; a_exp3 = 10'd40;
b_exp0 = 10'd619; b_exp1 = 10'd40; b_exp2 = 10'd277; b_exp3 = 10'd726;
a_sign0 = 4'd12; a_sign1 = 4'd13; a_sign2 = 4'd1; a_sign3 = 4'd0;
b_sign0 = 4'd9; b_sign1 = 4'd2; b_sign2 = 4'd2; b_sign3 = 4'd2;
@(posedge clk_i);
a_mant0 = 8'd48; a_mant1 = 8'd244; a_mant2 = 8'd181; a_mant3 = 8'd178;
b_mant0 = 8'd142; b_mant1 = 8'd42; b_mant2 = 8'd232; b_mant3 = 8'd34;
a_exp0 = 10'd965; a_exp1 = 10'd969; a_exp2 = 10'd124; a_exp3 = 10'd752;
b_exp0 = 10'd990; b_exp1 = 10'd527; b_exp2 = 10'd487; b_exp3 = 10'd25;
a_sign0 = 4'd13; a_sign1 = 4'd11; a_sign2 = 4'd5; a_sign3 = 4'd10;
b_sign0 = 4'd4; b_sign1 = 4'd10; b_sign2 = 4'd2; b_sign3 = 4'd13;
@(posedge clk_i);
a_mant0 = 8'd31; a_mant1 = 8'd108; a_mant2 = 8'd55; a_mant3 = 8'd96;
b_mant0 = 8'd39; b_mant1 = 8'd159; b_mant2 = 8'd165; b_mant3 = 8'd47;
a_exp0 = 10'd925; a_exp1 = 10'd284; a_exp2 = 10'd30; a_exp3 = 10'd736;
b_exp0 = 10'd350; b_exp1 = 10'd857; b_exp2 = 10'd517; b_exp3 = 10'd489;
a_sign0 = 4'd15; a_sign1 = 4'd3; a_sign2 = 4'd5; a_sign3 = 4'd15;
b_sign0 = 4'd4; b_sign1 = 4'd16; b_sign2 = 4'd5; b_sign3 = 4'd1;
@(posedge clk_i);
a_mant0 = 8'd72; a_mant1 = 8'd14; a_mant2 = 8'd96; a_mant3 = 8'd131;
b_mant0 = 8'd63; b_mant1 = 8'd6; b_mant2 = 8'd75; b_mant3 = 8'd104;
a_exp0 = 10'd350; a_exp1 = 10'd908; a_exp2 = 10'd16; a_exp3 = 10'd758;
b_exp0 = 10'd867; b_exp1 = 10'd118; b_exp2 = 10'd90; b_exp3 = 10'd454;
a_sign0 = 4'd5; a_sign1 = 4'd7; a_sign2 = 4'd13; a_sign3 = 4'd6;
b_sign0 = 4'd0; b_sign1 = 4'd2; b_sign2 = 4'd2; b_sign3 = 4'd1;
@(posedge clk_i);
a_mant0 = 8'd138; a_mant1 = 8'd235; a_mant2 = 8'd212; a_mant3 = 8'd25;
b_mant0 = 8'd47; b_mant1 = 8'd37; b_mant2 = 8'd141; b_mant3 = 8'd66;
a_exp0 = 10'd875; a_exp1 = 10'd928; a_exp2 = 10'd889; a_exp3 = 10'd331;
b_exp0 = 10'd913; b_exp1 = 10'd515; b_exp2 = 10'd20; b_exp3 = 10'd929;
a_sign0 = 4'd12; a_sign1 = 4'd2; a_sign2 = 4'd4; a_sign3 = 4'd0;
b_sign0 = 4'd3; b_sign1 = 4'd11; b_sign2 = 4'd15; b_sign3 = 4'd7;
@(posedge clk_i);
a_mant0 = 8'd120; a_mant1 = 8'd40; a_mant2 = 8'd187; a_mant3 = 8'd204;
b_mant0 = 8'd234; b_mant1 = 8'd121; b_mant2 = 8'd101; b_mant3 = 8'd83;
a_exp0 = 10'd846; a_exp1 = 10'd70; a_exp2 = 10'd813; a_exp3 = 10'd656;
b_exp0 = 10'd409; b_exp1 = 10'd531; b_exp2 = 10'd755; b_exp3 = 10'd740;
a_sign0 = 4'd10; a_sign1 = 4'd16; a_sign2 = 4'd0; a_sign3 = 4'd1;
b_sign0 = 4'd9; b_sign1 = 4'd6; b_sign2 = 4'd2; b_sign3 = 4'd3;
@(posedge clk_i);
shared_exps0 = 8'd125;
shared_exps1 = 8'd147;
a_mant0 = 8'd118; a_mant1 = 8'd100; a_mant2 = 8'd224; a_mant3 = 8'd217;
b_mant0 = 8'd1; b_mant1 = 8'd229; b_mant2 = 8'd186; b_mant3 = 8'd252;
a_exp0 = 10'd593; a_exp1 = 10'd727; a_exp2 = 10'd310; a_exp3 = 10'd30;
b_exp0 = 10'd256; b_exp1 = 10'd951; b_exp2 = 10'd780; b_exp3 = 10'd179;
a_sign0 = 4'd7; a_sign1 = 4'd9; a_sign2 = 4'd2; a_sign3 = 4'd13;
b_sign0 = 4'd4; b_sign1 = 4'd9; b_sign2 = 4'd12; b_sign3 = 4'd11;
@(posedge clk_i);
a_mant0 = 8'd163; a_mant1 = 8'd141; a_mant2 = 8'd217; a_mant3 = 8'd204;
b_mant0 = 8'd71; b_mant1 = 8'd212; b_mant2 = 8'd239; b_mant3 = 8'd215;
a_exp0 = 10'd504; a_exp1 = 10'd245; a_exp2 = 10'd258; a_exp3 = 10'd75;
b_exp0 = 10'd820; b_exp1 = 10'd594; b_exp2 = 10'd505; b_exp3 = 10'd256;
a_sign0 = 4'd9; a_sign1 = 4'd5; a_sign2 = 4'd16; a_sign3 = 4'd13;
b_sign0 = 4'd6; b_sign1 = 4'd1; b_sign2 = 4'd2; b_sign3 = 4'd2;
@(posedge clk_i);
a_mant0 = 8'd44; a_mant1 = 8'd12; a_mant2 = 8'd79; a_mant3 = 8'd238;
b_mant0 = 8'd1; b_mant1 = 8'd124; b_mant2 = 8'd233; b_mant3 = 8'd77;
a_exp0 = 10'd24; a_exp1 = 10'd830; a_exp2 = 10'd999; a_exp3 = 10'd455;
b_exp0 = 10'd495; b_exp1 = 10'd215; b_exp2 = 10'd969; b_exp3 = 10'd983;
a_sign0 = 4'd5; a_sign1 = 4'd6; a_sign2 = 4'd9; a_sign3 = 4'd7;
b_sign0 = 4'd8; b_sign1 = 4'd9; b_sign2 = 4'd9; b_sign3 = 4'd7;
@(posedge clk_i);
a_mant0 = 8'd161; a_mant1 = 8'd218; a_mant2 = 8'd56; a_mant3 = 8'd76;
b_mant0 = 8'd238; b_mant1 = 8'd209; b_mant2 = 8'd80; b_mant3 = 8'd163;
a_exp0 = 10'd220; a_exp1 = 10'd132; a_exp2 = 10'd969; a_exp3 = 10'd242;
b_exp0 = 10'd113; b_exp1 = 10'd15; b_exp2 = 10'd9; b_exp3 = 10'd96;
a_sign0 = 4'd8; a_sign1 = 4'd14; a_sign2 = 4'd12; a_sign3 = 4'd11;
b_sign0 = 4'd9; b_sign1 = 4'd3; b_sign2 = 4'd9; b_sign3 = 4'd4;
@(posedge clk_i);
a_mant0 = 8'd162; a_mant1 = 8'd55; a_mant2 = 8'd92; a_mant3 = 8'd216;
b_mant0 = 8'd251; b_mant1 = 8'd235; b_mant2 = 8'd86; b_mant3 = 8'd35;
a_exp0 = 10'd344; a_exp1 = 10'd371; a_exp2 = 10'd836; a_exp3 = 10'd44;
b_exp0 = 10'd961; b_exp1 = 10'd242; b_exp2 = 10'd471; b_exp3 = 10'd314;
a_sign0 = 4'd2; a_sign1 = 4'd9; a_sign2 = 4'd8; a_sign3 = 4'd13;
b_sign0 = 4'd1; b_sign1 = 4'd2; b_sign2 = 4'd4; b_sign3 = 4'd5;
@(posedge clk_i);
a_mant0 = 8'd192; a_mant1 = 8'd216; a_mant2 = 8'd172; a_mant3 = 8'd9;
b_mant0 = 8'd215; b_mant1 = 8'd72; b_mant2 = 8'd117; b_mant3 = 8'd142;
a_exp0 = 10'd667; a_exp1 = 10'd614; a_exp2 = 10'd604; a_exp3 = 10'd449;
b_exp0 = 10'd437; b_exp1 = 10'd671; b_exp2 = 10'd340; b_exp3 = 10'd834;
a_sign0 = 4'd5; a_sign1 = 4'd8; a_sign2 = 4'd2; a_sign3 = 4'd9;
b_sign0 = 4'd13; b_sign1 = 4'd4; b_sign2 = 4'd5; b_sign3 = 4'd4;
@(posedge clk_i);
a_mant0 = 8'd151; a_mant1 = 8'd143; a_mant2 = 8'd185; a_mant3 = 8'd1;
b_mant0 = 8'd213; b_mant1 = 8'd21; b_mant2 = 8'd66; b_mant3 = 8'd245;
a_exp0 = 10'd829; a_exp1 = 10'd850; a_exp2 = 10'd921; a_exp3 = 10'd1012;
b_exp0 = 10'd887; b_exp1 = 10'd731; b_exp2 = 10'd801; b_exp3 = 10'd588;
a_sign0 = 4'd15; a_sign1 = 4'd6; a_sign2 = 4'd11; a_sign3 = 4'd6;
b_sign0 = 4'd5; b_sign1 = 4'd16; b_sign2 = 4'd12; b_sign3 = 4'd12;
@(posedge clk_i);
a_mant0 = 8'd254; a_mant1 = 8'd205; a_mant2 = 8'd59; a_mant3 = 8'd15;
b_mant0 = 8'd245; b_mant1 = 8'd61; b_mant2 = 8'd76; b_mant3 = 8'd107;
a_exp0 = 10'd541; a_exp1 = 10'd713; a_exp2 = 10'd174; a_exp3 = 10'd563;
b_exp0 = 10'd654; b_exp1 = 10'd834; b_exp2 = 10'd590; b_exp3 = 10'd596;
a_sign0 = 4'd5; a_sign1 = 4'd0; a_sign2 = 4'd8; a_sign3 = 4'd0;
b_sign0 = 4'd12; b_sign1 = 4'd13; b_sign2 = 4'd12; b_sign3 = 4'd16;
@(posedge clk_i);
shared_exps0 = 8'd133;
shared_exps1 = 8'd146;
rstn = 0;
@(posedge clk_i);
rstn = 1;
a_mant0 = 8'd139; a_mant1 = 8'd234; a_mant2 = 8'd44; a_mant3 = 8'd84;
b_mant0 = 8'd185; b_mant1 = 8'd234; b_mant2 = 8'd75; b_mant3 = 8'd168;
a_exp0 = 10'd99; a_exp1 = 10'd967; a_exp2 = 10'd354; a_exp3 = 10'd560;
b_exp0 = 10'd797; b_exp1 = 10'd804; b_exp2 = 10'd576; b_exp3 = 10'd222;
a_sign0 = 4'd15; a_sign1 = 4'd7; a_sign2 = 4'd16; a_sign3 = 4'd13;
b_sign0 = 4'd11; b_sign1 = 4'd12; b_sign2 = 4'd4; b_sign3 = 4'd14;
@(posedge clk_i);
a_mant0 = 8'd5; a_mant1 = 8'd75; a_mant2 = 8'd59; a_mant3 = 8'd69;
b_mant0 = 8'd242; b_mant1 = 8'd95; b_mant2 = 8'd142; b_mant3 = 8'd130;
a_exp0 = 10'd53; a_exp1 = 10'd951; a_exp2 = 10'd644; a_exp3 = 10'd150;
b_exp0 = 10'd913; b_exp1 = 10'd507; b_exp2 = 10'd259; b_exp3 = 10'd302;
a_sign0 = 4'd0; a_sign1 = 4'd9; a_sign2 = 4'd8; a_sign3 = 4'd10;
b_sign0 = 4'd1; b_sign1 = 4'd0; b_sign2 = 4'd1; b_sign3 = 4'd15;
@(posedge clk_i);
a_mant0 = 8'd191; a_mant1 = 8'd236; a_mant2 = 8'd252; a_mant3 = 8'd88;
b_mant0 = 8'd191; b_mant1 = 8'd243; b_mant2 = 8'd253; b_mant3 = 8'd152;
a_exp0 = 10'd858; a_exp1 = 10'd804; a_exp2 = 10'd501; a_exp3 = 10'd26;
b_exp0 = 10'd98; b_exp1 = 10'd223; b_exp2 = 10'd355; b_exp3 = 10'd420;
a_sign0 = 4'd11; a_sign1 = 4'd8; a_sign2 = 4'd4; a_sign3 = 4'd4;
b_sign0 = 4'd13; b_sign1 = 4'd2; b_sign2 = 4'd9; b_sign3 = 4'd9;
@(posedge clk_i);
a_mant0 = 8'd27; a_mant1 = 8'd94; a_mant2 = 8'd140; a_mant3 = 8'd114;
b_mant0 = 8'd8; b_mant1 = 8'd91; b_mant2 = 8'd102; b_mant3 = 8'd151;
a_exp0 = 10'd197; a_exp1 = 10'd60; a_exp2 = 10'd211; a_exp3 = 10'd346;
b_exp0 = 10'd857; b_exp1 = 10'd866; b_exp2 = 10'd57; b_exp3 = 10'd770;
a_sign0 = 4'd5; a_sign1 = 4'd1; a_sign2 = 4'd2; a_sign3 = 4'd0;
b_sign0 = 4'd0; b_sign1 = 4'd16; b_sign2 = 4'd0; b_sign3 = 4'd11;
@(posedge clk_i);
a_mant0 = 8'd201; a_mant1 = 8'd132; a_mant2 = 8'd251; a_mant3 = 8'd175;
b_mant0 = 8'd82; b_mant1 = 8'd151; b_mant2 = 8'd195; b_mant3 = 8'd109;
a_exp0 = 10'd103; a_exp1 = 10'd731; a_exp2 = 10'd769; a_exp3 = 10'd472;
b_exp0 = 10'd624; b_exp1 = 10'd7; b_exp2 = 10'd552; b_exp3 = 10'd82;
a_sign0 = 4'd15; a_sign1 = 4'd2; a_sign2 = 4'd4; a_sign3 = 4'd13;
b_sign0 = 4'd13; b_sign1 = 4'd0; b_sign2 = 4'd16; b_sign3 = 4'd5;
@(posedge clk_i);
a_mant0 = 8'd86; a_mant1 = 8'd237; a_mant2 = 8'd88; a_mant3 = 8'd97;
b_mant0 = 8'd22; b_mant1 = 8'd20; b_mant2 = 8'd176; b_mant3 = 8'd68;
a_exp0 = 10'd880; a_exp1 = 10'd793; a_exp2 = 10'd87; a_exp3 = 10'd383;
b_exp0 = 10'd535; b_exp1 = 10'd333; b_exp2 = 10'd320; b_exp3 = 10'd416;
a_sign0 = 4'd9; a_sign1 = 4'd15; a_sign2 = 4'd12; a_sign3 = 4'd13;
b_sign0 = 4'd0; b_sign1 = 4'd7; b_sign2 = 4'd5; b_sign3 = 4'd16;
@(posedge clk_i);
a_mant0 = 8'd203; a_mant1 = 8'd157; a_mant2 = 8'd202; a_mant3 = 8'd143;
b_mant0 = 8'd48; b_mant1 = 8'd171; b_mant2 = 8'd205; b_mant3 = 8'd179;
a_exp0 = 10'd89; a_exp1 = 10'd214; a_exp2 = 10'd120; a_exp3 = 10'd661;
b_exp0 = 10'd469; b_exp1 = 10'd133; b_exp2 = 10'd347; b_exp3 = 10'd828;
a_sign0 = 4'd8; a_sign1 = 4'd11; a_sign2 = 4'd10; a_sign3 = 4'd0;
b_sign0 = 4'd5; b_sign1 = 4'd16; b_sign2 = 4'd3; b_sign3 = 4'd3;
@(posedge clk_i);
shared_exps0 = 8'd116;
shared_exps1 = 8'd137;
a_mant0 = 8'd164; a_mant1 = 8'd8; a_mant2 = 8'd49; a_mant3 = 8'd70;
b_mant0 = 8'd34; b_mant1 = 8'd133; b_mant2 = 8'd211; b_mant3 = 8'd81;
a_exp0 = 10'd751; a_exp1 = 10'd582; a_exp2 = 10'd357; a_exp3 = 10'd946;
b_exp0 = 10'd278; b_exp1 = 10'd894; b_exp2 = 10'd437; b_exp3 = 10'd513;
a_sign0 = 4'd10; a_sign1 = 4'd2; a_sign2 = 4'd4; a_sign3 = 4'd13;
b_sign0 = 4'd3; b_sign1 = 4'd6; b_sign2 = 4'd3; b_sign3 = 4'd15;
@(posedge clk_i);
a_mant0 = 8'd65; a_mant1 = 8'd140; a_mant2 = 8'd112; a_mant3 = 8'd246;
b_mant0 = 8'd204; b_mant1 = 8'd48; b_mant2 = 8'd237; b_mant3 = 8'd111;
a_exp0 = 10'd808; a_exp1 = 10'd919; a_exp2 = 10'd632; a_exp3 = 10'd957;
b_exp0 = 10'd925; b_exp1 = 10'd830; b_exp2 = 10'd14; b_exp3 = 10'd109;
a_sign0 = 4'd0; a_sign1 = 4'd12; a_sign2 = 4'd6; a_sign3 = 4'd13;
b_sign0 = 4'd14; b_sign1 = 4'd3; b_sign2 = 4'd5; b_sign3 = 4'd13;
@(posedge clk_i);
a_mant0 = 8'd188; a_mant1 = 8'd191; a_mant2 = 8'd70; a_mant3 = 8'd157;
b_mant0 = 8'd72; b_mant1 = 8'd14; b_mant2 = 8'd132; b_mant3 = 8'd149;
a_exp0 = 10'd71; a_exp1 = 10'd466; a_exp2 = 10'd500; a_exp3 = 10'd603;
b_exp0 = 10'd643; b_exp1 = 10'd783; b_exp2 = 10'd274; b_exp3 = 10'd330;
a_sign0 = 4'd0; a_sign1 = 4'd14; a_sign2 = 4'd3; a_sign3 = 4'd13;
b_sign0 = 4'd14; b_sign1 = 4'd9; b_sign2 = 4'd12; b_sign3 = 4'd15;
@(posedge clk_i);
a_mant0 = 8'd206; a_mant1 = 8'd111; a_mant2 = 8'd187; a_mant3 = 8'd77;
b_mant0 = 8'd134; b_mant1 = 8'd21; b_mant2 = 8'd188; b_mant3 = 8'd228;
a_exp0 = 10'd336; a_exp1 = 10'd556; a_exp2 = 10'd862; a_exp3 = 10'd232;
b_exp0 = 10'd930; b_exp1 = 10'd75; b_exp2 = 10'd424; b_exp3 = 10'd286;
a_sign0 = 4'd2; a_sign1 = 4'd7; a_sign2 = 4'd3; a_sign3 = 4'd8;
b_sign0 = 4'd6; b_sign1 = 4'd12; b_sign2 = 4'd6; b_sign3 = 4'd6;
@(posedge clk_i);
a_mant0 = 8'd179; a_mant1 = 8'd61; a_mant2 = 8'd147; a_mant3 = 8'd129;
b_mant0 = 8'd193; b_mant1 = 8'd242; b_mant2 = 8'd120; b_mant3 = 8'd38;
a_exp0 = 10'd164; a_exp1 = 10'd651; a_exp2 = 10'd473; a_exp3 = 10'd968;
b_exp0 = 10'd194; b_exp1 = 10'd888; b_exp2 = 10'd1014; b_exp3 = 10'd887;
a_sign0 = 4'd2; a_sign1 = 4'd4; a_sign2 = 4'd9; a_sign3 = 4'd16;
b_sign0 = 4'd7; b_sign1 = 4'd7; b_sign2 = 4'd15; b_sign3 = 4'd8;
@(posedge clk_i);
a_mant0 = 8'd40; a_mant1 = 8'd246; a_mant2 = 8'd53; a_mant3 = 8'd92;
b_mant0 = 8'd132; b_mant1 = 8'd19; b_mant2 = 8'd14; b_mant3 = 8'd92;
a_exp0 = 10'd560; a_exp1 = 10'd812; a_exp2 = 10'd469; a_exp3 = 10'd826;
b_exp0 = 10'd386; b_exp1 = 10'd765; b_exp2 = 10'd612; b_exp3 = 10'd265;
a_sign0 = 4'd14; a_sign1 = 4'd16; a_sign2 = 4'd8; a_sign3 = 4'd13;
b_sign0 = 4'd4; b_sign1 = 4'd5; b_sign2 = 4'd10; b_sign3 = 4'd5;
@(posedge clk_i);
a_mant0 = 8'd249; a_mant1 = 8'd188; a_mant2 = 8'd174; a_mant3 = 8'd23;
b_mant0 = 8'd197; b_mant1 = 8'd215; b_mant2 = 8'd241; b_mant3 = 8'd77;
a_exp0 = 10'd1003; a_exp1 = 10'd130; a_exp2 = 10'd443; a_exp3 = 10'd654;
b_exp0 = 10'd592; b_exp1 = 10'd648; b_exp2 = 10'd676; b_exp3 = 10'd969;
a_sign0 = 4'd10; a_sign1 = 4'd10; a_sign2 = 4'd2; a_sign3 = 4'd12;
b_sign0 = 4'd13; b_sign1 = 4'd4; b_sign2 = 4'd2; b_sign3 = 4'd0;
@(posedge clk_i);
a_mant0 = 8'd205; a_mant1 = 8'd232; a_mant2 = 8'd27; a_mant3 = 8'd86;
b_mant0 = 8'd55; b_mant1 = 8'd52; b_mant2 = 8'd76; b_mant3 = 8'd95;
a_exp0 = 10'd890; a_exp1 = 10'd353; a_exp2 = 10'd712; a_exp3 = 10'd728;
b_exp0 = 10'd995; b_exp1 = 10'd719; b_exp2 = 10'd578; b_exp3 = 10'd896;
a_sign0 = 4'd0; a_sign1 = 4'd7; a_sign2 = 4'd1; a_sign3 = 4'd8;
b_sign0 = 4'd0; b_sign1 = 4'd1; b_sign2 = 4'd6; b_sign3 = 4'd14;
@(posedge clk_i);
shared_exps0 = 8'd122;
shared_exps1 = 8'd118;
a_mant0 = 8'd81; a_mant1 = 8'd220; a_mant2 = 8'd245; a_mant3 = 8'd136;
b_mant0 = 8'd109; b_mant1 = 8'd197; b_mant2 = 8'd60; b_mant3 = 8'd53;
a_exp0 = 10'd644; a_exp1 = 10'd891; a_exp2 = 10'd994; a_exp3 = 10'd157;
b_exp0 = 10'd54; b_exp1 = 10'd148; b_exp2 = 10'd959; b_exp3 = 10'd572;
a_sign0 = 4'd15; a_sign1 = 4'd1; a_sign2 = 4'd13; a_sign3 = 4'd3;
b_sign0 = 4'd9; b_sign1 = 4'd8; b_sign2 = 4'd5; b_sign3 = 4'd3;
@(posedge clk_i);
a_mant0 = 8'd181; a_mant1 = 8'd55; a_mant2 = 8'd122; a_mant3 = 8'd255;
b_mant0 = 8'd128; b_mant1 = 8'd176; b_mant2 = 8'd124; b_mant3 = 8'd140;
a_exp0 = 10'd236; a_exp1 = 10'd7; a_exp2 = 10'd346; a_exp3 = 10'd240;
b_exp0 = 10'd319; b_exp1 = 10'd1003; b_exp2 = 10'd137; b_exp3 = 10'd568;
a_sign0 = 4'd6; a_sign1 = 4'd13; a_sign2 = 4'd6; a_sign3 = 4'd7;
b_sign0 = 4'd0; b_sign1 = 4'd0; b_sign2 = 4'd12; b_sign3 = 4'd14;
@(posedge clk_i);
a_mant0 = 8'd228; a_mant1 = 8'd107; a_mant2 = 8'd79; a_mant3 = 8'd59;
b_mant0 = 8'd194; b_mant1 = 8'd112; b_mant2 = 8'd185; b_mant3 = 8'd51;
a_exp0 = 10'd917; a_exp1 = 10'd140; a_exp2 = 10'd782; a_exp3 = 10'd971;
b_exp0 = 10'd411; b_exp1 = 10'd591; b_exp2 = 10'd482; b_exp3 = 10'd870;
a_sign0 = 4'd1; a_sign1 = 4'd10; a_sign2 = 4'd8; a_sign3 = 4'd10;
b_sign0 = 4'd2; b_sign1 = 4'd16; b_sign2 = 4'd0; b_sign3 = 4'd9;
@(posedge clk_i);
a_mant0 = 8'd225; a_mant1 = 8'd180; a_mant2 = 8'd151; a_mant3 = 8'd113;
b_mant0 = 8'd105; b_mant1 = 8'd225; b_mant2 = 8'd196; b_mant3 = 8'd132;
a_exp0 = 10'd747; a_exp1 = 10'd630; a_exp2 = 10'd456; a_exp3 = 10'd772;
b_exp0 = 10'd473; b_exp1 = 10'd291; b_exp2 = 10'd911; b_exp3 = 10'd540;
a_sign0 = 4'd10; a_sign1 = 4'd3; a_sign2 = 4'd7; a_sign3 = 4'd2;
b_sign0 = 4'd14; b_sign1 = 4'd11; b_sign2 = 4'd16; b_sign3 = 4'd8;
@(posedge clk_i);
a_mant0 = 8'd121; a_mant1 = 8'd97; a_mant2 = 8'd197; a_mant3 = 8'd72;
b_mant0 = 8'd8; b_mant1 = 8'd115; b_mant2 = 8'd77; b_mant3 = 8'd23;
a_exp0 = 10'd854; a_exp1 = 10'd516; a_exp2 = 10'd645; a_exp3 = 10'd484;
b_exp0 = 10'd244; b_exp1 = 10'd494; b_exp2 = 10'd472; b_exp3 = 10'd151;
a_sign0 = 4'd8; a_sign1 = 4'd7; a_sign2 = 4'd0; a_sign3 = 4'd4;
b_sign0 = 4'd0; b_sign1 = 4'd6; b_sign2 = 4'd13; b_sign3 = 4'd4;
@(posedge clk_i);
a_mant0 = 8'd125; a_mant1 = 8'd167; a_mant2 = 8'd39; a_mant3 = 8'd14;
b_mant0 = 8'd227; b_mant1 = 8'd222; b_mant2 = 8'd96; b_mant3 = 8'd74;
a_exp0 = 10'd542; a_exp1 = 10'd912; a_exp2 = 10'd971; a_exp3 = 10'd726;
b_exp0 = 10'd254; b_exp1 = 10'd1020; b_exp2 = 10'd166; b_exp3 = 10'd553;
a_sign0 = 4'd6; a_sign1 = 4'd7; a_sign2 = 4'd16; a_sign3 = 4'd14;
b_sign0 = 4'd6; b_sign1 = 4'd1; b_sign2 = 4'd3; b_sign3 = 4'd13;
@(posedge clk_i);
a_mant0 = 8'd221; a_mant1 = 8'd163; a_mant2 = 8'd26; a_mant3 = 8'd196;
b_mant0 = 8'd96; b_mant1 = 8'd154; b_mant2 = 8'd169; b_mant3 = 8'd149;
a_exp0 = 10'd529; a_exp1 = 10'd370; a_exp2 = 10'd2; a_exp3 = 10'd726;
b_exp0 = 10'd126; b_exp1 = 10'd9; b_exp2 = 10'd361; b_exp3 = 10'd39;
a_sign0 = 4'd13; a_sign1 = 4'd15; a_sign2 = 4'd8; a_sign3 = 4'd11;
b_sign0 = 4'd11; b_sign1 = 4'd11; b_sign2 = 4'd6; b_sign3 = 4'd16;
@(posedge clk_i);
a_mant0 = 8'd253; a_mant1 = 8'd27; a_mant2 = 8'd101; a_mant3 = 8'd12;
b_mant0 = 8'd64; b_mant1 = 8'd153; b_mant2 = 8'd196; b_mant3 = 8'd178;
a_exp0 = 10'd434; a_exp1 = 10'd120; a_exp2 = 10'd446; a_exp3 = 10'd860;
b_exp0 = 10'd146; b_exp1 = 10'd390; b_exp2 = 10'd524; b_exp3 = 10'd128;
a_sign0 = 4'd4; a_sign1 = 4'd11; a_sign2 = 4'd10; a_sign3 = 4'd10;
b_sign0 = 4'd14; b_sign1 = 4'd8; b_sign2 = 4'd12; b_sign3 = 4'd7;
@(posedge clk_i);
shared_exps0 = 8'd111;
shared_exps1 = 8'd136;
a_mant0 = 8'd100; a_mant1 = 8'd224; a_mant2 = 8'd79; a_mant3 = 8'd95;
b_mant0 = 8'd244; b_mant1 = 8'd136; b_mant2 = 8'd32; b_mant3 = 8'd44;
a_exp0 = 10'd911; a_exp1 = 10'd291; a_exp2 = 10'd833; a_exp3 = 10'd60;
b_exp0 = 10'd348; b_exp1 = 10'd7; b_exp2 = 10'd24; b_exp3 = 10'd208;
a_sign0 = 4'd5; a_sign1 = 4'd2; a_sign2 = 4'd7; a_sign3 = 4'd12;
b_sign0 = 4'd2; b_sign1 = 4'd7; b_sign2 = 4'd9; b_sign3 = 4'd10;
@(posedge clk_i);
a_mant0 = 8'd24; a_mant1 = 8'd180; a_mant2 = 8'd95; a_mant3 = 8'd77;
b_mant0 = 8'd46; b_mant1 = 8'd34; b_mant2 = 8'd252; b_mant3 = 8'd216;
a_exp0 = 10'd92; a_exp1 = 10'd900; a_exp2 = 10'd973; a_exp3 = 10'd35;
b_exp0 = 10'd452; b_exp1 = 10'd752; b_exp2 = 10'd954; b_exp3 = 10'd715;
a_sign0 = 4'd8; a_sign1 = 4'd3; a_sign2 = 4'd2; a_sign3 = 4'd14;
b_sign0 = 4'd15; b_sign1 = 4'd13; b_sign2 = 4'd16; b_sign3 = 4'd6;
@(posedge clk_i);
a_mant0 = 8'd163; a_mant1 = 8'd85; a_mant2 = 8'd196; a_mant3 = 8'd13;
b_mant0 = 8'd223; b_mant1 = 8'd241; b_mant2 = 8'd125; b_mant3 = 8'd114;
a_exp0 = 10'd12; a_exp1 = 10'd427; a_exp2 = 10'd79; a_exp3 = 10'd666;
b_exp0 = 10'd822; b_exp1 = 10'd277; b_exp2 = 10'd360; b_exp3 = 10'd582;
a_sign0 = 4'd12; a_sign1 = 4'd4; a_sign2 = 4'd9; a_sign3 = 4'd15;
b_sign0 = 4'd9; b_sign1 = 4'd2; b_sign2 = 4'd12; b_sign3 = 4'd9;
@(posedge clk_i);
a_mant0 = 8'd84; a_mant1 = 8'd46; a_mant2 = 8'd205; a_mant3 = 8'd165;
b_mant0 = 8'd13; b_mant1 = 8'd116; b_mant2 = 8'd157; b_mant3 = 8'd140;
a_exp0 = 10'd448; a_exp1 = 10'd752; a_exp2 = 10'd31; a_exp3 = 10'd141;
b_exp0 = 10'd5; b_exp1 = 10'd904; b_exp2 = 10'd123; b_exp3 = 10'd292;
a_sign0 = 4'd2; a_sign1 = 4'd16; a_sign2 = 4'd16; a_sign3 = 4'd10;
b_sign0 = 4'd4; b_sign1 = 4'd8; b_sign2 = 4'd6; b_sign3 = 4'd9;
@(posedge clk_i);
a_mant0 = 8'd96; a_mant1 = 8'd12; a_mant2 = 8'd25; a_mant3 = 8'd141;
b_mant0 = 8'd72; b_mant1 = 8'd190; b_mant2 = 8'd133; b_mant3 = 8'd178;
a_exp0 = 10'd14; a_exp1 = 10'd906; a_exp2 = 10'd377; a_exp3 = 10'd151;
b_exp0 = 10'd926; b_exp1 = 10'd462; b_exp2 = 10'd220; b_exp3 = 10'd773;
a_sign0 = 4'd10; a_sign1 = 4'd11; a_sign2 = 4'd6; a_sign3 = 4'd9;
b_sign0 = 4'd6; b_sign1 = 4'd12; b_sign2 = 4'd1; b_sign3 = 4'd14;
@(posedge clk_i);
a_mant0 = 8'd22; a_mant1 = 8'd77; a_mant2 = 8'd207; a_mant3 = 8'd208;
b_mant0 = 8'd234; b_mant1 = 8'd18; b_mant2 = 8'd231; b_mant3 = 8'd202;
a_exp0 = 10'd115; a_exp1 = 10'd292; a_exp2 = 10'd549; a_exp3 = 10'd571;
b_exp0 = 10'd196; b_exp1 = 10'd455; b_exp2 = 10'd333; b_exp3 = 10'd376;
a_sign0 = 4'd10; a_sign1 = 4'd0; a_sign2 = 4'd5; a_sign3 = 4'd9;
b_sign0 = 4'd2; b_sign1 = 4'd1; b_sign2 = 4'd9; b_sign3 = 4'd2;
@(posedge clk_i);
a_mant0 = 8'd28; a_mant1 = 8'd126; a_mant2 = 8'd37; a_mant3 = 8'd49;
b_mant0 = 8'd84; b_mant1 = 8'd52; b_mant2 = 8'd50; b_mant3 = 8'd232;
a_exp0 = 10'd589; a_exp1 = 10'd496; a_exp2 = 10'd468; a_exp3 = 10'd880;
b_exp0 = 10'd718; b_exp1 = 10'd836; b_exp2 = 10'd28; b_exp3 = 10'd864;
a_sign0 = 4'd8; a_sign1 = 4'd8; a_sign2 = 4'd15; a_sign3 = 4'd1;
b_sign0 = 4'd1; b_sign1 = 4'd9; b_sign2 = 4'd10; b_sign3 = 4'd15;
@(posedge clk_i);
a_mant0 = 8'd99; a_mant1 = 8'd210; a_mant2 = 8'd255; a_mant3 = 8'd0;
b_mant0 = 8'd37; b_mant1 = 8'd248; b_mant2 = 8'd186; b_mant3 = 8'd97;
a_exp0 = 10'd717; a_exp1 = 10'd995; a_exp2 = 10'd53; a_exp3 = 10'd515;
b_exp0 = 10'd536; b_exp1 = 10'd983; b_exp2 = 10'd31; b_exp3 = 10'd326;
a_sign0 = 4'd16; a_sign1 = 4'd0; a_sign2 = 4'd6; a_sign3 = 4'd9;
b_sign0 = 4'd16; b_sign1 = 4'd1; b_sign2 = 4'd1; b_sign3 = 4'd12;
@(posedge clk_i);
shared_exps0 = 8'd112;
shared_exps1 = 8'd127;
rstn = 0;
@(posedge clk_i);
rstn = 1;
a_mant0 = 8'd155; a_mant1 = 8'd3; a_mant2 = 8'd4; a_mant3 = 8'd94;
b_mant0 = 8'd231; b_mant1 = 8'd2; b_mant2 = 8'd246; b_mant3 = 8'd228;
a_exp0 = 10'd520; a_exp1 = 10'd399; a_exp2 = 10'd25; a_exp3 = 10'd709;
b_exp0 = 10'd186; b_exp1 = 10'd332; b_exp2 = 10'd254; b_exp3 = 10'd105;
a_sign0 = 4'd10; a_sign1 = 4'd11; a_sign2 = 4'd6; a_sign3 = 4'd11;
b_sign0 = 4'd8; b_sign1 = 4'd7; b_sign2 = 4'd3; b_sign3 = 4'd8;
@(posedge clk_i);
a_mant0 = 8'd32; a_mant1 = 8'd32; a_mant2 = 8'd104; a_mant3 = 8'd239;
b_mant0 = 8'd151; b_mant1 = 8'd225; b_mant2 = 8'd106; b_mant3 = 8'd1;
a_exp0 = 10'd985; a_exp1 = 10'd906; a_exp2 = 10'd587; a_exp3 = 10'd494;
b_exp0 = 10'd238; b_exp1 = 10'd1020; b_exp2 = 10'd173; b_exp3 = 10'd872;
a_sign0 = 4'd16; a_sign1 = 4'd0; a_sign2 = 4'd6; a_sign3 = 4'd15;
b_sign0 = 4'd3; b_sign1 = 4'd15; b_sign2 = 4'd14; b_sign3 = 4'd6;
@(posedge clk_i);
a_mant0 = 8'd255; a_mant1 = 8'd250; a_mant2 = 8'd33; a_mant3 = 8'd109;
b_mant0 = 8'd5; b_mant1 = 8'd199; b_mant2 = 8'd247; b_mant3 = 8'd76;
a_exp0 = 10'd699; a_exp1 = 10'd592; a_exp2 = 10'd592; a_exp3 = 10'd389;
b_exp0 = 10'd986; b_exp1 = 10'd414; b_exp2 = 10'd893; b_exp3 = 10'd484;
a_sign0 = 4'd8; a_sign1 = 4'd1; a_sign2 = 4'd1; a_sign3 = 4'd5;
b_sign0 = 4'd1; b_sign1 = 4'd8; b_sign2 = 4'd3; b_sign3 = 4'd9;
@(posedge clk_i);
a_mant0 = 8'd39; a_mant1 = 8'd146; a_mant2 = 8'd8; a_mant3 = 8'd213;
b_mant0 = 8'd212; b_mant1 = 8'd69; b_mant2 = 8'd135; b_mant3 = 8'd252;
a_exp0 = 10'd242; a_exp1 = 10'd233; a_exp2 = 10'd228; a_exp3 = 10'd411;
b_exp0 = 10'd405; b_exp1 = 10'd216; b_exp2 = 10'd601; b_exp3 = 10'd720;
a_sign0 = 4'd6; a_sign1 = 4'd8; a_sign2 = 4'd0; a_sign3 = 4'd16;
b_sign0 = 4'd9; b_sign1 = 4'd8; b_sign2 = 4'd6; b_sign3 = 4'd2;
@(posedge clk_i);
a_mant0 = 8'd129; a_mant1 = 8'd71; a_mant2 = 8'd213; a_mant3 = 8'd219;
b_mant0 = 8'd229; b_mant1 = 8'd54; b_mant2 = 8'd224; b_mant3 = 8'd243;
a_exp0 = 10'd50; a_exp1 = 10'd160; a_exp2 = 10'd148; a_exp3 = 10'd191;
b_exp0 = 10'd90; b_exp1 = 10'd685; b_exp2 = 10'd997; b_exp3 = 10'd737;
a_sign0 = 4'd15; a_sign1 = 4'd16; a_sign2 = 4'd6; a_sign3 = 4'd13;
b_sign0 = 4'd3; b_sign1 = 4'd8; b_sign2 = 4'd12; b_sign3 = 4'd6;
@(posedge clk_i);
a_mant0 = 8'd29; a_mant1 = 8'd159; a_mant2 = 8'd59; a_mant3 = 8'd85;
b_mant0 = 8'd233; b_mant1 = 8'd105; b_mant2 = 8'd45; b_mant3 = 8'd207;
a_exp0 = 10'd367; a_exp1 = 10'd777; a_exp2 = 10'd625; a_exp3 = 10'd129;
b_exp0 = 10'd839; b_exp1 = 10'd764; b_exp2 = 10'd600; b_exp3 = 10'd664;
a_sign0 = 4'd8; a_sign1 = 4'd13; a_sign2 = 4'd11; a_sign3 = 4'd15;
b_sign0 = 4'd6; b_sign1 = 4'd14; b_sign2 = 4'd7; b_sign3 = 4'd15;
@(posedge clk_i);
a_mant0 = 8'd170; a_mant1 = 8'd204; a_mant2 = 8'd67; a_mant3 = 8'd211;
b_mant0 = 8'd135; b_mant1 = 8'd164; b_mant2 = 8'd179; b_mant3 = 8'd33;
a_exp0 = 10'd442; a_exp1 = 10'd43; a_exp2 = 10'd181; a_exp3 = 10'd446;
b_exp0 = 10'd392; b_exp1 = 10'd176; b_exp2 = 10'd843; b_exp3 = 10'd435;
a_sign0 = 4'd4; a_sign1 = 4'd5; a_sign2 = 4'd15; a_sign3 = 4'd12;
b_sign0 = 4'd9; b_sign1 = 4'd1; b_sign2 = 4'd10; b_sign3 = 4'd1;
@(posedge clk_i);
shared_exps0 = 8'd143;
shared_exps1 = 8'd127;
a_mant0 = 8'd190; a_mant1 = 8'd244; a_mant2 = 8'd90; a_mant3 = 8'd76;
b_mant0 = 8'd216; b_mant1 = 8'd183; b_mant2 = 8'd122; b_mant3 = 8'd167;
a_exp0 = 10'd824; a_exp1 = 10'd144; a_exp2 = 10'd708; a_exp3 = 10'd477;
b_exp0 = 10'd608; b_exp1 = 10'd824; b_exp2 = 10'd453; b_exp3 = 10'd81;
a_sign0 = 4'd8; a_sign1 = 4'd3; a_sign2 = 4'd2; a_sign3 = 4'd8;
b_sign0 = 4'd10; b_sign1 = 4'd9; b_sign2 = 4'd3; b_sign3 = 4'd5;
@(posedge clk_i);
a_mant0 = 8'd208; a_mant1 = 8'd209; a_mant2 = 8'd109; a_mant3 = 8'd176;
b_mant0 = 8'd70; b_mant1 = 8'd241; b_mant2 = 8'd32; b_mant3 = 8'd199;
a_exp0 = 10'd314; a_exp1 = 10'd870; a_exp2 = 10'd219; a_exp3 = 10'd970;
b_exp0 = 10'd824; b_exp1 = 10'd189; b_exp2 = 10'd566; b_exp3 = 10'd869;
a_sign0 = 4'd12; a_sign1 = 4'd6; a_sign2 = 4'd14; a_sign3 = 4'd8;
b_sign0 = 4'd5; b_sign1 = 4'd14; b_sign2 = 4'd1; b_sign3 = 4'd12;
@(posedge clk_i);
a_mant0 = 8'd134; a_mant1 = 8'd54; a_mant2 = 8'd156; a_mant3 = 8'd254;
b_mant0 = 8'd136; b_mant1 = 8'd36; b_mant2 = 8'd149; b_mant3 = 8'd8;
a_exp0 = 10'd263; a_exp1 = 10'd489; a_exp2 = 10'd866; a_exp3 = 10'd193;
b_exp0 = 10'd735; b_exp1 = 10'd261; b_exp2 = 10'd479; b_exp3 = 10'd802;
a_sign0 = 4'd16; a_sign1 = 4'd3; a_sign2 = 4'd15; a_sign3 = 4'd0;
b_sign0 = 4'd4; b_sign1 = 4'd1; b_sign2 = 4'd4; b_sign3 = 4'd1;
@(posedge clk_i);
a_mant0 = 8'd188; a_mant1 = 8'd137; a_mant2 = 8'd36; a_mant3 = 8'd206;
b_mant0 = 8'd75; b_mant1 = 8'd94; b_mant2 = 8'd196; b_mant3 = 8'd158;
a_exp0 = 10'd272; a_exp1 = 10'd997; a_exp2 = 10'd273; a_exp3 = 10'd334;
b_exp0 = 10'd889; b_exp1 = 10'd407; b_exp2 = 10'd876; b_exp3 = 10'd0;
a_sign0 = 4'd4; a_sign1 = 4'd4; a_sign2 = 4'd9; a_sign3 = 4'd10;
b_sign0 = 4'd11; b_sign1 = 4'd3; b_sign2 = 4'd11; b_sign3 = 4'd5;
@(posedge clk_i);
a_mant0 = 8'd241; a_mant1 = 8'd233; a_mant2 = 8'd203; a_mant3 = 8'd55;
b_mant0 = 8'd130; b_mant1 = 8'd230; b_mant2 = 8'd214; b_mant3 = 8'd122;
a_exp0 = 10'd641; a_exp1 = 10'd62; a_exp2 = 10'd931; a_exp3 = 10'd231;
b_exp0 = 10'd70; b_exp1 = 10'd0; b_exp2 = 10'd916; b_exp3 = 10'd348;
a_sign0 = 4'd7; a_sign1 = 4'd8; a_sign2 = 4'd2; a_sign3 = 4'd2;
b_sign0 = 4'd8; b_sign1 = 4'd7; b_sign2 = 4'd1; b_sign3 = 4'd1;
@(posedge clk_i);
a_mant0 = 8'd66; a_mant1 = 8'd226; a_mant2 = 8'd30; a_mant3 = 8'd201;
b_mant0 = 8'd209; b_mant1 = 8'd183; b_mant2 = 8'd68; b_mant3 = 8'd103;
a_exp0 = 10'd735; a_exp1 = 10'd748; a_exp2 = 10'd837; a_exp3 = 10'd57;
b_exp0 = 10'd287; b_exp1 = 10'd64; b_exp2 = 10'd54; b_exp3 = 10'd525;
a_sign0 = 4'd5; a_sign1 = 4'd4; a_sign2 = 4'd14; a_sign3 = 4'd0;
b_sign0 = 4'd9; b_sign1 = 4'd3; b_sign2 = 4'd12; b_sign3 = 4'd3;
@(posedge clk_i);
a_mant0 = 8'd3; a_mant1 = 8'd185; a_mant2 = 8'd1; a_mant3 = 8'd30;
b_mant0 = 8'd221; b_mant1 = 8'd233; b_mant2 = 8'd138; b_mant3 = 8'd246;
a_exp0 = 10'd671; a_exp1 = 10'd354; a_exp2 = 10'd57; a_exp3 = 10'd381;
b_exp0 = 10'd424; b_exp1 = 10'd805; b_exp2 = 10'd38; b_exp3 = 10'd685;
a_sign0 = 4'd11; a_sign1 = 4'd1; a_sign2 = 4'd0; a_sign3 = 4'd10;
b_sign0 = 4'd10; b_sign1 = 4'd7; b_sign2 = 4'd16; b_sign3 = 4'd14;
@(posedge clk_i);
a_mant0 = 8'd151; a_mant1 = 8'd141; a_mant2 = 8'd207; a_mant3 = 8'd186;
b_mant0 = 8'd41; b_mant1 = 8'd133; b_mant2 = 8'd165; b_mant3 = 8'd246;
a_exp0 = 10'd39; a_exp1 = 10'd108; a_exp2 = 10'd624; a_exp3 = 10'd874;
b_exp0 = 10'd302; b_exp1 = 10'd97; b_exp2 = 10'd103; b_exp3 = 10'd185;
a_sign0 = 4'd3; a_sign1 = 4'd16; a_sign2 = 4'd4; a_sign3 = 4'd9;
b_sign0 = 4'd8; b_sign1 = 4'd7; b_sign2 = 4'd10; b_sign3 = 4'd13;
@(posedge clk_i);
shared_exps0 = 8'd82;
shared_exps1 = 8'd140;
a_mant0 = 8'd231; a_mant1 = 8'd161; a_mant2 = 8'd71; a_mant3 = 8'd243;
b_mant0 = 8'd217; b_mant1 = 8'd163; b_mant2 = 8'd215; b_mant3 = 8'd75;
a_exp0 = 10'd121; a_exp1 = 10'd973; a_exp2 = 10'd117; a_exp3 = 10'd295;
b_exp0 = 10'd315; b_exp1 = 10'd720; b_exp2 = 10'd269; b_exp3 = 10'd654;
a_sign0 = 4'd10; a_sign1 = 4'd6; a_sign2 = 4'd1; a_sign3 = 4'd3;
b_sign0 = 4'd6; b_sign1 = 4'd13; b_sign2 = 4'd6; b_sign3 = 4'd9;
@(posedge clk_i);
a_mant0 = 8'd11; a_mant1 = 8'd91; a_mant2 = 8'd229; a_mant3 = 8'd126;
b_mant0 = 8'd208; b_mant1 = 8'd201; b_mant2 = 8'd167; b_mant3 = 8'd0;
a_exp0 = 10'd327; a_exp1 = 10'd131; a_exp2 = 10'd727; a_exp3 = 10'd692;
b_exp0 = 10'd622; b_exp1 = 10'd27; b_exp2 = 10'd411; b_exp3 = 10'd246;
a_sign0 = 4'd3; a_sign1 = 4'd7; a_sign2 = 4'd8; a_sign3 = 4'd0;
b_sign0 = 4'd3; b_sign1 = 4'd12; b_sign2 = 4'd2; b_sign3 = 4'd0;
@(posedge clk_i);
a_mant0 = 8'd64; a_mant1 = 8'd124; a_mant2 = 8'd207; a_mant3 = 8'd128;
b_mant0 = 8'd66; b_mant1 = 8'd38; b_mant2 = 8'd207; b_mant3 = 8'd238;
a_exp0 = 10'd245; a_exp1 = 10'd719; a_exp2 = 10'd442; a_exp3 = 10'd350;
b_exp0 = 10'd821; b_exp1 = 10'd510; b_exp2 = 10'd266; b_exp3 = 10'd57;
a_sign0 = 4'd8; a_sign1 = 4'd13; a_sign2 = 4'd8; a_sign3 = 4'd14;
b_sign0 = 4'd2; b_sign1 = 4'd3; b_sign2 = 4'd3; b_sign3 = 4'd5;
@(posedge clk_i);
a_mant0 = 8'd167; a_mant1 = 8'd204; a_mant2 = 8'd61; a_mant3 = 8'd107;
b_mant0 = 8'd88; b_mant1 = 8'd38; b_mant2 = 8'd57; b_mant3 = 8'd67;
a_exp0 = 10'd272; a_exp1 = 10'd711; a_exp2 = 10'd237; a_exp3 = 10'd243;
b_exp0 = 10'd86; b_exp1 = 10'd494; b_exp2 = 10'd899; b_exp3 = 10'd646;
a_sign0 = 4'd7; a_sign1 = 4'd0; a_sign2 = 4'd12; a_sign3 = 4'd11;
b_sign0 = 4'd1; b_sign1 = 4'd16; b_sign2 = 4'd11; b_sign3 = 4'd14;
@(posedge clk_i);
a_mant0 = 8'd174; a_mant1 = 8'd237; a_mant2 = 8'd85; a_mant3 = 8'd176;
b_mant0 = 8'd216; b_mant1 = 8'd238; b_mant2 = 8'd198; b_mant3 = 8'd103;
a_exp0 = 10'd482; a_exp1 = 10'd330; a_exp2 = 10'd979; a_exp3 = 10'd479;
b_exp0 = 10'd975; b_exp1 = 10'd641; b_exp2 = 10'd191; b_exp3 = 10'd323;
a_sign0 = 4'd7; a_sign1 = 4'd12; a_sign2 = 4'd16; a_sign3 = 4'd1;
b_sign0 = 4'd8; b_sign1 = 4'd4; b_sign2 = 4'd1; b_sign3 = 4'd16;
@(posedge clk_i);
a_mant0 = 8'd222; a_mant1 = 8'd165; a_mant2 = 8'd170; a_mant3 = 8'd74;
b_mant0 = 8'd51; b_mant1 = 8'd237; b_mant2 = 8'd230; b_mant3 = 8'd181;
a_exp0 = 10'd795; a_exp1 = 10'd596; a_exp2 = 10'd71; a_exp3 = 10'd177;
b_exp0 = 10'd917; b_exp1 = 10'd156; b_exp2 = 10'd980; b_exp3 = 10'd123;
a_sign0 = 4'd8; a_sign1 = 4'd5; a_sign2 = 4'd13; a_sign3 = 4'd0;
b_sign0 = 4'd2; b_sign1 = 4'd13; b_sign2 = 4'd13; b_sign3 = 4'd8;
@(posedge clk_i);
a_mant0 = 8'd49; a_mant1 = 8'd41; a_mant2 = 8'd169; a_mant3 = 8'd84;
b_mant0 = 8'd130; b_mant1 = 8'd26; b_mant2 = 8'd2; b_mant3 = 8'd214;
a_exp0 = 10'd287; a_exp1 = 10'd697; a_exp2 = 10'd960; a_exp3 = 10'd1005;
b_exp0 = 10'd798; b_exp1 = 10'd650; b_exp2 = 10'd587; b_exp3 = 10'd74;
a_sign0 = 4'd2; a_sign1 = 4'd16; a_sign2 = 4'd8; a_sign3 = 4'd4;
b_sign0 = 4'd15; b_sign1 = 4'd15; b_sign2 = 4'd10; b_sign3 = 4'd7;
@(posedge clk_i);
a_mant0 = 8'd17; a_mant1 = 8'd99; a_mant2 = 8'd193; a_mant3 = 8'd254;
b_mant0 = 8'd111; b_mant1 = 8'd30; b_mant2 = 8'd207; b_mant3 = 8'd143;
a_exp0 = 10'd878; a_exp1 = 10'd652; a_exp2 = 10'd696; a_exp3 = 10'd141;
b_exp0 = 10'd526; b_exp1 = 10'd918; b_exp2 = 10'd242; b_exp3 = 10'd256;
a_sign0 = 4'd10; a_sign1 = 4'd0; a_sign2 = 4'd10; a_sign3 = 4'd3;
b_sign0 = 4'd11; b_sign1 = 4'd14; b_sign2 = 4'd8; b_sign3 = 4'd13;
@(posedge clk_i);
shared_exps0 = 8'd151;
shared_exps1 = 8'd122;
a_mant0 = 8'd67; a_mant1 = 8'd89; a_mant2 = 8'd19; a_mant3 = 8'd59;
b_mant0 = 8'd89; b_mant1 = 8'd11; b_mant2 = 8'd174; b_mant3 = 8'd44;
a_exp0 = 10'd523; a_exp1 = 10'd893; a_exp2 = 10'd616; a_exp3 = 10'd48;
b_exp0 = 10'd363; b_exp1 = 10'd547; b_exp2 = 10'd300; b_exp3 = 10'd343;
a_sign0 = 4'd1; a_sign1 = 4'd3; a_sign2 = 4'd11; a_sign3 = 4'd7;
b_sign0 = 4'd1; b_sign1 = 4'd3; b_sign2 = 4'd12; b_sign3 = 4'd15;
@(posedge clk_i);
a_mant0 = 8'd252; a_mant1 = 8'd191; a_mant2 = 8'd124; a_mant3 = 8'd69;
b_mant0 = 8'd162; b_mant1 = 8'd160; b_mant2 = 8'd238; b_mant3 = 8'd36;
a_exp0 = 10'd686; a_exp1 = 10'd40; a_exp2 = 10'd982; a_exp3 = 10'd645;
b_exp0 = 10'd451; b_exp1 = 10'd38; b_exp2 = 10'd238; b_exp3 = 10'd974;
a_sign0 = 4'd12; a_sign1 = 4'd13; a_sign2 = 4'd10; a_sign3 = 4'd8;
b_sign0 = 4'd9; b_sign1 = 4'd11; b_sign2 = 4'd4; b_sign3 = 4'd8;
@(posedge clk_i);
a_mant0 = 8'd22; a_mant1 = 8'd142; a_mant2 = 8'd217; a_mant3 = 8'd56;
b_mant0 = 8'd0; b_mant1 = 8'd4; b_mant2 = 8'd169; b_mant3 = 8'd129;
a_exp0 = 10'd942; a_exp1 = 10'd157; a_exp2 = 10'd467; a_exp3 = 10'd95;
b_exp0 = 10'd321; b_exp1 = 10'd558; b_exp2 = 10'd690; b_exp3 = 10'd964;
a_sign0 = 4'd15; a_sign1 = 4'd12; a_sign2 = 4'd10; a_sign3 = 4'd12;
b_sign0 = 4'd16; b_sign1 = 4'd13; b_sign2 = 4'd16; b_sign3 = 4'd3;
@(posedge clk_i);
a_mant0 = 8'd91; a_mant1 = 8'd119; a_mant2 = 8'd153; a_mant3 = 8'd135;
b_mant0 = 8'd238; b_mant1 = 8'd113; b_mant2 = 8'd32; b_mant3 = 8'd204;
a_exp0 = 10'd489; a_exp1 = 10'd456; a_exp2 = 10'd602; a_exp3 = 10'd194;
b_exp0 = 10'd563; b_exp1 = 10'd381; b_exp2 = 10'd428; b_exp3 = 10'd1008;
a_sign0 = 4'd15; a_sign1 = 4'd8; a_sign2 = 4'd7; a_sign3 = 4'd12;
b_sign0 = 4'd12; b_sign1 = 4'd16; b_sign2 = 4'd10; b_sign3 = 4'd14;
@(posedge clk_i);
a_mant0 = 8'd30; a_mant1 = 8'd21; a_mant2 = 8'd193; a_mant3 = 8'd77;
b_mant0 = 8'd158; b_mant1 = 8'd131; b_mant2 = 8'd162; b_mant3 = 8'd251;
a_exp0 = 10'd11; a_exp1 = 10'd525; a_exp2 = 10'd508; a_exp3 = 10'd697;
b_exp0 = 10'd946; b_exp1 = 10'd335; b_exp2 = 10'd600; b_exp3 = 10'd975;
a_sign0 = 4'd12; a_sign1 = 4'd8; a_sign2 = 4'd1; a_sign3 = 4'd9;
b_sign0 = 4'd2; b_sign1 = 4'd13; b_sign2 = 4'd2; b_sign3 = 4'd10;
@(posedge clk_i);
a_mant0 = 8'd130; a_mant1 = 8'd99; a_mant2 = 8'd60; a_mant3 = 8'd176;
b_mant0 = 8'd14; b_mant1 = 8'd124; b_mant2 = 8'd238; b_mant3 = 8'd19;
a_exp0 = 10'd333; a_exp1 = 10'd421; a_exp2 = 10'd761; a_exp3 = 10'd520;
b_exp0 = 10'd251; b_exp1 = 10'd810; b_exp2 = 10'd482; b_exp3 = 10'd575;
a_sign0 = 4'd15; a_sign1 = 4'd13; a_sign2 = 4'd8; a_sign3 = 4'd14;
b_sign0 = 4'd2; b_sign1 = 4'd5; b_sign2 = 4'd2; b_sign3 = 4'd12;
@(posedge clk_i);
a_mant0 = 8'd79; a_mant1 = 8'd242; a_mant2 = 8'd176; a_mant3 = 8'd204;
b_mant0 = 8'd168; b_mant1 = 8'd47; b_mant2 = 8'd87; b_mant3 = 8'd33;
a_exp0 = 10'd170; a_exp1 = 10'd667; a_exp2 = 10'd499; a_exp3 = 10'd410;
b_exp0 = 10'd307; b_exp1 = 10'd80; b_exp2 = 10'd699; b_exp3 = 10'd505;
a_sign0 = 4'd2; a_sign1 = 4'd8; a_sign2 = 4'd11; a_sign3 = 4'd15;
b_sign0 = 4'd2; b_sign1 = 4'd15; b_sign2 = 4'd16; b_sign3 = 4'd13;
@(posedge clk_i);
a_mant0 = 8'd55; a_mant1 = 8'd56; a_mant2 = 8'd206; a_mant3 = 8'd240;
b_mant0 = 8'd79; b_mant1 = 8'd10; b_mant2 = 8'd178; b_mant3 = 8'd211;
a_exp0 = 10'd245; a_exp1 = 10'd699; a_exp2 = 10'd419; a_exp3 = 10'd584;
b_exp0 = 10'd521; b_exp1 = 10'd67; b_exp2 = 10'd242; b_exp3 = 10'd714;
a_sign0 = 4'd2; a_sign1 = 4'd12; a_sign2 = 4'd15; a_sign3 = 4'd2;
b_sign0 = 4'd2; b_sign1 = 4'd3; b_sign2 = 4'd3; b_sign3 = 4'd2;
@(posedge clk_i);
shared_exps0 = 8'd129;
shared_exps1 = 8'd154;
rstn = 0;
@(posedge clk_i);
rstn = 1;
a_mant0 = 8'd91; a_mant1 = 8'd43; a_mant2 = 8'd111; a_mant3 = 8'd156;
b_mant0 = 8'd213; b_mant1 = 8'd100; b_mant2 = 8'd207; b_mant3 = 8'd9;
a_exp0 = 10'd609; a_exp1 = 10'd947; a_exp2 = 10'd195; a_exp3 = 10'd59;
b_exp0 = 10'd978; b_exp1 = 10'd799; b_exp2 = 10'd215; b_exp3 = 10'd479;
a_sign0 = 4'd3; a_sign1 = 4'd8; a_sign2 = 4'd7; a_sign3 = 4'd13;
b_sign0 = 4'd6; b_sign1 = 4'd14; b_sign2 = 4'd0; b_sign3 = 4'd3;
@(posedge clk_i);
a_mant0 = 8'd95; a_mant1 = 8'd86; a_mant2 = 8'd134; a_mant3 = 8'd20;
b_mant0 = 8'd155; b_mant1 = 8'd47; b_mant2 = 8'd241; b_mant3 = 8'd150;
a_exp0 = 10'd746; a_exp1 = 10'd293; a_exp2 = 10'd815; a_exp3 = 10'd344;
b_exp0 = 10'd40; b_exp1 = 10'd661; b_exp2 = 10'd821; b_exp3 = 10'd572;
a_sign0 = 4'd14; a_sign1 = 4'd7; a_sign2 = 4'd14; a_sign3 = 4'd16;
b_sign0 = 4'd7; b_sign1 = 4'd6; b_sign2 = 4'd13; b_sign3 = 4'd1;
@(posedge clk_i);
a_mant0 = 8'd67; a_mant1 = 8'd79; a_mant2 = 8'd100; a_mant3 = 8'd241;
b_mant0 = 8'd103; b_mant1 = 8'd78; b_mant2 = 8'd20; b_mant3 = 8'd88;
a_exp0 = 10'd400; a_exp1 = 10'd991; a_exp2 = 10'd860; a_exp3 = 10'd456;
b_exp0 = 10'd422; b_exp1 = 10'd602; b_exp2 = 10'd969; b_exp3 = 10'd761;
a_sign0 = 4'd0; a_sign1 = 4'd4; a_sign2 = 4'd16; a_sign3 = 4'd13;
b_sign0 = 4'd1; b_sign1 = 4'd6; b_sign2 = 4'd0; b_sign3 = 4'd7;
@(posedge clk_i);
a_mant0 = 8'd189; a_mant1 = 8'd16; a_mant2 = 8'd139; a_mant3 = 8'd179;
b_mant0 = 8'd88; b_mant1 = 8'd197; b_mant2 = 8'd230; b_mant3 = 8'd229;
a_exp0 = 10'd224; a_exp1 = 10'd497; a_exp2 = 10'd255; a_exp3 = 10'd500;
b_exp0 = 10'd498; b_exp1 = 10'd39; b_exp2 = 10'd82; b_exp3 = 10'd381;
a_sign0 = 4'd3; a_sign1 = 4'd8; a_sign2 = 4'd12; a_sign3 = 4'd13;
b_sign0 = 4'd0; b_sign1 = 4'd7; b_sign2 = 4'd9; b_sign3 = 4'd15;
@(posedge clk_i);
a_mant0 = 8'd179; a_mant1 = 8'd236; a_mant2 = 8'd225; a_mant3 = 8'd253;
b_mant0 = 8'd153; b_mant1 = 8'd33; b_mant2 = 8'd159; b_mant3 = 8'd224;
a_exp0 = 10'd968; a_exp1 = 10'd25; a_exp2 = 10'd359; a_exp3 = 10'd67;
b_exp0 = 10'd609; b_exp1 = 10'd756; b_exp2 = 10'd801; b_exp3 = 10'd79;
a_sign0 = 4'd5; a_sign1 = 4'd6; a_sign2 = 4'd3; a_sign3 = 4'd11;
b_sign0 = 4'd14; b_sign1 = 4'd12; b_sign2 = 4'd2; b_sign3 = 4'd11;
@(posedge clk_i);
a_mant0 = 8'd9; a_mant1 = 8'd207; a_mant2 = 8'd240; a_mant3 = 8'd127;
b_mant0 = 8'd30; b_mant1 = 8'd132; b_mant2 = 8'd214; b_mant3 = 8'd169;
a_exp0 = 10'd648; a_exp1 = 10'd694; a_exp2 = 10'd896; a_exp3 = 10'd75;
b_exp0 = 10'd1003; b_exp1 = 10'd716; b_exp2 = 10'd337; b_exp3 = 10'd224;
a_sign0 = 4'd6; a_sign1 = 4'd5; a_sign2 = 4'd5; a_sign3 = 4'd0;
b_sign0 = 4'd10; b_sign1 = 4'd9; b_sign2 = 4'd3; b_sign3 = 4'd11;
@(posedge clk_i);
a_mant0 = 8'd236; a_mant1 = 8'd197; a_mant2 = 8'd176; a_mant3 = 8'd32;
b_mant0 = 8'd38; b_mant1 = 8'd160; b_mant2 = 8'd108; b_mant3 = 8'd248;
a_exp0 = 10'd758; a_exp1 = 10'd998; a_exp2 = 10'd684; a_exp3 = 10'd787;
b_exp0 = 10'd532; b_exp1 = 10'd685; b_exp2 = 10'd499; b_exp3 = 10'd927;
a_sign0 = 4'd9; a_sign1 = 4'd1; a_sign2 = 4'd15; a_sign3 = 4'd12;
b_sign0 = 4'd13; b_sign1 = 4'd7; b_sign2 = 4'd6; b_sign3 = 4'd11;
@(posedge clk_i);
shared_exps0 = 8'd149;
shared_exps1 = 8'd154;
a_mant0 = 8'd81; a_mant1 = 8'd163; a_mant2 = 8'd43; a_mant3 = 8'd180;
b_mant0 = 8'd26; b_mant1 = 8'd25; b_mant2 = 8'd68; b_mant3 = 8'd18;
a_exp0 = 10'd586; a_exp1 = 10'd569; a_exp2 = 10'd149; a_exp3 = 10'd203;
b_exp0 = 10'd677; b_exp1 = 10'd52; b_exp2 = 10'd782; b_exp3 = 10'd795;
a_sign0 = 4'd12; a_sign1 = 4'd9; a_sign2 = 4'd3; a_sign3 = 4'd16;
b_sign0 = 4'd3; b_sign1 = 4'd6; b_sign2 = 4'd12; b_sign3 = 4'd16;
@(posedge clk_i);
a_mant0 = 8'd97; a_mant1 = 8'd86; a_mant2 = 8'd41; a_mant3 = 8'd160;
b_mant0 = 8'd118; b_mant1 = 8'd4; b_mant2 = 8'd177; b_mant3 = 8'd75;
a_exp0 = 10'd64; a_exp1 = 10'd740; a_exp2 = 10'd282; a_exp3 = 10'd250;
b_exp0 = 10'd627; b_exp1 = 10'd830; b_exp2 = 10'd747; b_exp3 = 10'd323;
a_sign0 = 4'd0; a_sign1 = 4'd4; a_sign2 = 4'd10; a_sign3 = 4'd14;
b_sign0 = 4'd12; b_sign1 = 4'd11; b_sign2 = 4'd9; b_sign3 = 4'd0;
@(posedge clk_i);
a_mant0 = 8'd186; a_mant1 = 8'd105; a_mant2 = 8'd139; a_mant3 = 8'd63;
b_mant0 = 8'd149; b_mant1 = 8'd102; b_mant2 = 8'd57; b_mant3 = 8'd180;
a_exp0 = 10'd629; a_exp1 = 10'd417; a_exp2 = 10'd178; a_exp3 = 10'd87;
b_exp0 = 10'd1001; b_exp1 = 10'd562; b_exp2 = 10'd613; b_exp3 = 10'd795;
a_sign0 = 4'd6; a_sign1 = 4'd0; a_sign2 = 4'd14; a_sign3 = 4'd13;
b_sign0 = 4'd5; b_sign1 = 4'd12; b_sign2 = 4'd13; b_sign3 = 4'd5;
@(posedge clk_i);
a_mant0 = 8'd206; a_mant1 = 8'd110; a_mant2 = 8'd9; a_mant3 = 8'd125;
b_mant0 = 8'd37; b_mant1 = 8'd41; b_mant2 = 8'd61; b_mant3 = 8'd20;
a_exp0 = 10'd135; a_exp1 = 10'd890; a_exp2 = 10'd38; a_exp3 = 10'd798;
b_exp0 = 10'd497; b_exp1 = 10'd1021; b_exp2 = 10'd974; b_exp3 = 10'd669;
a_sign0 = 4'd5; a_sign1 = 4'd15; a_sign2 = 4'd8; a_sign3 = 4'd12;
b_sign0 = 4'd10; b_sign1 = 4'd2; b_sign2 = 4'd14; b_sign3 = 4'd15;
@(posedge clk_i);
a_mant0 = 8'd208; a_mant1 = 8'd142; a_mant2 = 8'd37; a_mant3 = 8'd21;
b_mant0 = 8'd10; b_mant1 = 8'd130; b_mant2 = 8'd135; b_mant3 = 8'd92;
a_exp0 = 10'd472; a_exp1 = 10'd571; a_exp2 = 10'd357; a_exp3 = 10'd696;
b_exp0 = 10'd96; b_exp1 = 10'd876; b_exp2 = 10'd37; b_exp3 = 10'd657;
a_sign0 = 4'd6; a_sign1 = 4'd4; a_sign2 = 4'd12; a_sign3 = 4'd15;
b_sign0 = 4'd9; b_sign1 = 4'd7; b_sign2 = 4'd2; b_sign3 = 4'd6;
@(posedge clk_i);
a_mant0 = 8'd192; a_mant1 = 8'd249; a_mant2 = 8'd100; a_mant3 = 8'd153;
b_mant0 = 8'd172; b_mant1 = 8'd6; b_mant2 = 8'd76; b_mant3 = 8'd58;
a_exp0 = 10'd463; a_exp1 = 10'd89; a_exp2 = 10'd140; a_exp3 = 10'd756;
b_exp0 = 10'd224; b_exp1 = 10'd107; b_exp2 = 10'd444; b_exp3 = 10'd933;
a_sign0 = 4'd6; a_sign1 = 4'd0; a_sign2 = 4'd13; a_sign3 = 4'd5;
b_sign0 = 4'd3; b_sign1 = 4'd14; b_sign2 = 4'd16; b_sign3 = 4'd7;
@(posedge clk_i);
a_mant0 = 8'd227; a_mant1 = 8'd39; a_mant2 = 8'd112; a_mant3 = 8'd224;
b_mant0 = 8'd242; b_mant1 = 8'd101; b_mant2 = 8'd244; b_mant3 = 8'd87;
a_exp0 = 10'd203; a_exp1 = 10'd309; a_exp2 = 10'd760; a_exp3 = 10'd47;
b_exp0 = 10'd654; b_exp1 = 10'd22; b_exp2 = 10'd703; b_exp3 = 10'd817;
a_sign0 = 4'd1; a_sign1 = 4'd5; a_sign2 = 4'd10; a_sign3 = 4'd8;
b_sign0 = 4'd10; b_sign1 = 4'd8; b_sign2 = 4'd4; b_sign3 = 4'd4;
@(posedge clk_i);
a_mant0 = 8'd55; a_mant1 = 8'd50; a_mant2 = 8'd117; a_mant3 = 8'd136;
b_mant0 = 8'd155; b_mant1 = 8'd175; b_mant2 = 8'd134; b_mant3 = 8'd15;
a_exp0 = 10'd128; a_exp1 = 10'd994; a_exp2 = 10'd617; a_exp3 = 10'd451;
b_exp0 = 10'd384; b_exp1 = 10'd494; b_exp2 = 10'd852; b_exp3 = 10'd893;
a_sign0 = 4'd6; a_sign1 = 4'd11; a_sign2 = 4'd3; a_sign3 = 4'd11;
b_sign0 = 4'd5; b_sign1 = 4'd10; b_sign2 = 4'd2; b_sign3 = 4'd2;
@(posedge clk_i);
shared_exps0 = 8'd93;
shared_exps1 = 8'd144;
a_mant0 = 8'd173; a_mant1 = 8'd121; a_mant2 = 8'd10; a_mant3 = 8'd211;
b_mant0 = 8'd73; b_mant1 = 8'd88; b_mant2 = 8'd51; b_mant3 = 8'd84;
a_exp0 = 10'd806; a_exp1 = 10'd490; a_exp2 = 10'd949; a_exp3 = 10'd861;
b_exp0 = 10'd1010; b_exp1 = 10'd462; b_exp2 = 10'd69; b_exp3 = 10'd734;
a_sign0 = 4'd16; a_sign1 = 4'd1; a_sign2 = 4'd13; a_sign3 = 4'd10;
b_sign0 = 4'd14; b_sign1 = 4'd11; b_sign2 = 4'd10; b_sign3 = 4'd4;
@(posedge clk_i);
a_mant0 = 8'd175; a_mant1 = 8'd100; a_mant2 = 8'd191; a_mant3 = 8'd63;
b_mant0 = 8'd24; b_mant1 = 8'd61; b_mant2 = 8'd19; b_mant3 = 8'd96;
a_exp0 = 10'd318; a_exp1 = 10'd511; a_exp2 = 10'd278; a_exp3 = 10'd317;
b_exp0 = 10'd641; b_exp1 = 10'd821; b_exp2 = 10'd177; b_exp3 = 10'd957;
a_sign0 = 4'd9; a_sign1 = 4'd7; a_sign2 = 4'd0; a_sign3 = 4'd5;
b_sign0 = 4'd12; b_sign1 = 4'd5; b_sign2 = 4'd10; b_sign3 = 4'd0;
@(posedge clk_i);
a_mant0 = 8'd86; a_mant1 = 8'd153; a_mant2 = 8'd4; a_mant3 = 8'd179;
b_mant0 = 8'd228; b_mant1 = 8'd100; b_mant2 = 8'd158; b_mant3 = 8'd172;
a_exp0 = 10'd810; a_exp1 = 10'd772; a_exp2 = 10'd642; a_exp3 = 10'd1000;
b_exp0 = 10'd225; b_exp1 = 10'd593; b_exp2 = 10'd973; b_exp3 = 10'd840;
a_sign0 = 4'd14; a_sign1 = 4'd5; a_sign2 = 4'd14; a_sign3 = 4'd3;
b_sign0 = 4'd1; b_sign1 = 4'd4; b_sign2 = 4'd11; b_sign3 = 4'd2;
@(posedge clk_i);
a_mant0 = 8'd153; a_mant1 = 8'd150; a_mant2 = 8'd197; a_mant3 = 8'd38;
b_mant0 = 8'd194; b_mant1 = 8'd29; b_mant2 = 8'd156; b_mant3 = 8'd252;
a_exp0 = 10'd600; a_exp1 = 10'd443; a_exp2 = 10'd545; a_exp3 = 10'd12;
b_exp0 = 10'd567; b_exp1 = 10'd610; b_exp2 = 10'd552; b_exp3 = 10'd828;
a_sign0 = 4'd16; a_sign1 = 4'd12; a_sign2 = 4'd16; a_sign3 = 4'd5;
b_sign0 = 4'd11; b_sign1 = 4'd10; b_sign2 = 4'd13; b_sign3 = 4'd13;
@(posedge clk_i);
a_mant0 = 8'd233; a_mant1 = 8'd195; a_mant2 = 8'd63; a_mant3 = 8'd199;
b_mant0 = 8'd167; b_mant1 = 8'd46; b_mant2 = 8'd163; b_mant3 = 8'd122;
a_exp0 = 10'd315; a_exp1 = 10'd493; a_exp2 = 10'd899; a_exp3 = 10'd22;
b_exp0 = 10'd689; b_exp1 = 10'd179; b_exp2 = 10'd669; b_exp3 = 10'd137;
a_sign0 = 4'd4; a_sign1 = 4'd3; a_sign2 = 4'd2; a_sign3 = 4'd8;
b_sign0 = 4'd1; b_sign1 = 4'd12; b_sign2 = 4'd13; b_sign3 = 4'd1;
@(posedge clk_i);
a_mant0 = 8'd247; a_mant1 = 8'd180; a_mant2 = 8'd228; a_mant3 = 8'd240;
b_mant0 = 8'd123; b_mant1 = 8'd159; b_mant2 = 8'd1; b_mant3 = 8'd243;
a_exp0 = 10'd144; a_exp1 = 10'd861; a_exp2 = 10'd368; a_exp3 = 10'd88;
b_exp0 = 10'd423; b_exp1 = 10'd662; b_exp2 = 10'd459; b_exp3 = 10'd382;
a_sign0 = 4'd6; a_sign1 = 4'd13; a_sign2 = 4'd4; a_sign3 = 4'd14;
b_sign0 = 4'd10; b_sign1 = 4'd11; b_sign2 = 4'd8; b_sign3 = 4'd6;
@(posedge clk_i);
a_mant0 = 8'd179; a_mant1 = 8'd11; a_mant2 = 8'd235; a_mant3 = 8'd53;
b_mant0 = 8'd205; b_mant1 = 8'd67; b_mant2 = 8'd231; b_mant3 = 8'd190;
a_exp0 = 10'd233; a_exp1 = 10'd251; a_exp2 = 10'd1009; a_exp3 = 10'd679;
b_exp0 = 10'd214; b_exp1 = 10'd936; b_exp2 = 10'd535; b_exp3 = 10'd850;
a_sign0 = 4'd15; a_sign1 = 4'd4; a_sign2 = 4'd0; a_sign3 = 4'd16;
b_sign0 = 4'd10; b_sign1 = 4'd10; b_sign2 = 4'd8; b_sign3 = 4'd15;
@(posedge clk_i);
a_mant0 = 8'd60; a_mant1 = 8'd149; a_mant2 = 8'd26; a_mant3 = 8'd4;
b_mant0 = 8'd92; b_mant1 = 8'd157; b_mant2 = 8'd122; b_mant3 = 8'd22;
a_exp0 = 10'd179; a_exp1 = 10'd17; a_exp2 = 10'd953; a_exp3 = 10'd705;
b_exp0 = 10'd92; b_exp1 = 10'd0; b_exp2 = 10'd1002; b_exp3 = 10'd183;
a_sign0 = 4'd3; a_sign1 = 4'd12; a_sign2 = 4'd11; a_sign3 = 4'd8;
b_sign0 = 4'd8; b_sign1 = 4'd1; b_sign2 = 4'd7; b_sign3 = 4'd11;
@(posedge clk_i);
shared_exps0 = 8'd105;
shared_exps1 = 8'd104;
a_mant0 = 8'd218; a_mant1 = 8'd210; a_mant2 = 8'd142; a_mant3 = 8'd68;
b_mant0 = 8'd4; b_mant1 = 8'd184; b_mant2 = 8'd190; b_mant3 = 8'd248;
a_exp0 = 10'd765; a_exp1 = 10'd900; a_exp2 = 10'd803; a_exp3 = 10'd478;
b_exp0 = 10'd95; b_exp1 = 10'd258; b_exp2 = 10'd20; b_exp3 = 10'd500;
a_sign0 = 4'd13; a_sign1 = 4'd2; a_sign2 = 4'd8; a_sign3 = 4'd12;
b_sign0 = 4'd11; b_sign1 = 4'd1; b_sign2 = 4'd14; b_sign3 = 4'd16;
@(posedge clk_i);
a_mant0 = 8'd183; a_mant1 = 8'd182; a_mant2 = 8'd185; a_mant3 = 8'd129;
b_mant0 = 8'd109; b_mant1 = 8'd74; b_mant2 = 8'd156; b_mant3 = 8'd23;
a_exp0 = 10'd398; a_exp1 = 10'd493; a_exp2 = 10'd955; a_exp3 = 10'd981;
b_exp0 = 10'd709; b_exp1 = 10'd62; b_exp2 = 10'd888; b_exp3 = 10'd561;
a_sign0 = 4'd13; a_sign1 = 4'd8; a_sign2 = 4'd6; a_sign3 = 4'd13;
b_sign0 = 4'd12; b_sign1 = 4'd4; b_sign2 = 4'd14; b_sign3 = 4'd5;
@(posedge clk_i);
a_mant0 = 8'd11; a_mant1 = 8'd74; a_mant2 = 8'd226; a_mant3 = 8'd171;
b_mant0 = 8'd67; b_mant1 = 8'd143; b_mant2 = 8'd21; b_mant3 = 8'd252;
a_exp0 = 10'd691; a_exp1 = 10'd862; a_exp2 = 10'd764; a_exp3 = 10'd235;
b_exp0 = 10'd454; b_exp1 = 10'd508; b_exp2 = 10'd325; b_exp3 = 10'd383;
a_sign0 = 4'd5; a_sign1 = 4'd8; a_sign2 = 4'd3; a_sign3 = 4'd2;
b_sign0 = 4'd16; b_sign1 = 4'd3; b_sign2 = 4'd12; b_sign3 = 4'd15;
@(posedge clk_i);
a_mant0 = 8'd42; a_mant1 = 8'd122; a_mant2 = 8'd23; a_mant3 = 8'd105;
b_mant0 = 8'd57; b_mant1 = 8'd72; b_mant2 = 8'd238; b_mant3 = 8'd237;
a_exp0 = 10'd439; a_exp1 = 10'd23; a_exp2 = 10'd473; a_exp3 = 10'd411;
b_exp0 = 10'd385; b_exp1 = 10'd419; b_exp2 = 10'd670; b_exp3 = 10'd662;
a_sign0 = 4'd15; a_sign1 = 4'd3; a_sign2 = 4'd9; a_sign3 = 4'd2;
b_sign0 = 4'd6; b_sign1 = 4'd4; b_sign2 = 4'd16; b_sign3 = 4'd2;
@(posedge clk_i);
a_mant0 = 8'd203; a_mant1 = 8'd210; a_mant2 = 8'd153; a_mant3 = 8'd37;
b_mant0 = 8'd141; b_mant1 = 8'd169; b_mant2 = 8'd246; b_mant3 = 8'd12;
a_exp0 = 10'd148; a_exp1 = 10'd806; a_exp2 = 10'd668; a_exp3 = 10'd830;
b_exp0 = 10'd48; b_exp1 = 10'd733; b_exp2 = 10'd702; b_exp3 = 10'd1022;
a_sign0 = 4'd12; a_sign1 = 4'd11; a_sign2 = 4'd0; a_sign3 = 4'd5;
b_sign0 = 4'd9; b_sign1 = 4'd10; b_sign2 = 4'd16; b_sign3 = 4'd14;
@(posedge clk_i);
a_mant0 = 8'd120; a_mant1 = 8'd166; a_mant2 = 8'd245; a_mant3 = 8'd29;
b_mant0 = 8'd23; b_mant1 = 8'd192; b_mant2 = 8'd96; b_mant3 = 8'd23;
a_exp0 = 10'd167; a_exp1 = 10'd694; a_exp2 = 10'd122; a_exp3 = 10'd592;
b_exp0 = 10'd497; b_exp1 = 10'd452; b_exp2 = 10'd71; b_exp3 = 10'd832;
a_sign0 = 4'd7; a_sign1 = 4'd0; a_sign2 = 4'd16; a_sign3 = 4'd4;
b_sign0 = 4'd4; b_sign1 = 4'd0; b_sign2 = 4'd10; b_sign3 = 4'd14;
@(posedge clk_i);
a_mant0 = 8'd138; a_mant1 = 8'd203; a_mant2 = 8'd141; a_mant3 = 8'd230;
b_mant0 = 8'd99; b_mant1 = 8'd159; b_mant2 = 8'd138; b_mant3 = 8'd140;
a_exp0 = 10'd456; a_exp1 = 10'd380; a_exp2 = 10'd961; a_exp3 = 10'd722;
b_exp0 = 10'd64; b_exp1 = 10'd182; b_exp2 = 10'd460; b_exp3 = 10'd89;
a_sign0 = 4'd12; a_sign1 = 4'd3; a_sign2 = 4'd13; a_sign3 = 4'd5;
b_sign0 = 4'd12; b_sign1 = 4'd16; b_sign2 = 4'd2; b_sign3 = 4'd7;
@(posedge clk_i);
a_mant0 = 8'd23; a_mant1 = 8'd31; a_mant2 = 8'd115; a_mant3 = 8'd219;
b_mant0 = 8'd151; b_mant1 = 8'd26; b_mant2 = 8'd187; b_mant3 = 8'd50;
a_exp0 = 10'd275; a_exp1 = 10'd513; a_exp2 = 10'd536; a_exp3 = 10'd69;
b_exp0 = 10'd286; b_exp1 = 10'd535; b_exp2 = 10'd0; b_exp3 = 10'd334;
a_sign0 = 4'd4; a_sign1 = 4'd14; a_sign2 = 4'd1; a_sign3 = 4'd10;
b_sign0 = 4'd3; b_sign1 = 4'd6; b_sign2 = 4'd8; b_sign3 = 4'd9;
@(posedge clk_i);
shared_exps0 = 8'd148;
shared_exps1 = 8'd111;
rstn = 0;
@(posedge clk_i);
rstn = 1;
a_mant0 = 8'd100; a_mant1 = 8'd243; a_mant2 = 8'd67; a_mant3 = 8'd217;
b_mant0 = 8'd160; b_mant1 = 8'd252; b_mant2 = 8'd121; b_mant3 = 8'd117;
a_exp0 = 10'd398; a_exp1 = 10'd965; a_exp2 = 10'd473; a_exp3 = 10'd960;
b_exp0 = 10'd604; b_exp1 = 10'd856; b_exp2 = 10'd408; b_exp3 = 10'd178;
a_sign0 = 4'd6; a_sign1 = 4'd13; a_sign2 = 4'd16; a_sign3 = 4'd6;
b_sign0 = 4'd15; b_sign1 = 4'd5; b_sign2 = 4'd5; b_sign3 = 4'd1;
@(posedge clk_i);
a_mant0 = 8'd170; a_mant1 = 8'd236; a_mant2 = 8'd206; a_mant3 = 8'd245;
b_mant0 = 8'd166; b_mant1 = 8'd237; b_mant2 = 8'd208; b_mant3 = 8'd85;
a_exp0 = 10'd256; a_exp1 = 10'd336; a_exp2 = 10'd382; a_exp3 = 10'd276;
b_exp0 = 10'd810; b_exp1 = 10'd10; b_exp2 = 10'd839; b_exp3 = 10'd237;
a_sign0 = 4'd6; a_sign1 = 4'd9; a_sign2 = 4'd13; a_sign3 = 4'd11;
b_sign0 = 4'd4; b_sign1 = 4'd8; b_sign2 = 4'd14; b_sign3 = 4'd8;
@(posedge clk_i);
a_mant0 = 8'd94; a_mant1 = 8'd138; a_mant2 = 8'd182; a_mant3 = 8'd73;
b_mant0 = 8'd142; b_mant1 = 8'd27; b_mant2 = 8'd131; b_mant3 = 8'd65;
a_exp0 = 10'd228; a_exp1 = 10'd716; a_exp2 = 10'd464; a_exp3 = 10'd42;
b_exp0 = 10'd409; b_exp1 = 10'd354; b_exp2 = 10'd496; b_exp3 = 10'd614;
a_sign0 = 4'd3; a_sign1 = 4'd14; a_sign2 = 4'd15; a_sign3 = 4'd12;
b_sign0 = 4'd1; b_sign1 = 4'd10; b_sign2 = 4'd11; b_sign3 = 4'd9;
@(posedge clk_i);
a_mant0 = 8'd112; a_mant1 = 8'd230; a_mant2 = 8'd180; a_mant3 = 8'd19;
b_mant0 = 8'd62; b_mant1 = 8'd85; b_mant2 = 8'd165; b_mant3 = 8'd22;
a_exp0 = 10'd799; a_exp1 = 10'd169; a_exp2 = 10'd4; a_exp3 = 10'd858;
b_exp0 = 10'd454; b_exp1 = 10'd418; b_exp2 = 10'd704; b_exp3 = 10'd547;
a_sign0 = 4'd9; a_sign1 = 4'd6; a_sign2 = 4'd6; a_sign3 = 4'd9;
b_sign0 = 4'd4; b_sign1 = 4'd8; b_sign2 = 4'd2; b_sign3 = 4'd10;
@(posedge clk_i);
a_mant0 = 8'd246; a_mant1 = 8'd66; a_mant2 = 8'd139; a_mant3 = 8'd162;
b_mant0 = 8'd201; b_mant1 = 8'd67; b_mant2 = 8'd16; b_mant3 = 8'd190;
a_exp0 = 10'd867; a_exp1 = 10'd499; a_exp2 = 10'd248; a_exp3 = 10'd333;
b_exp0 = 10'd331; b_exp1 = 10'd452; b_exp2 = 10'd331; b_exp3 = 10'd811;
a_sign0 = 4'd0; a_sign1 = 4'd9; a_sign2 = 4'd7; a_sign3 = 4'd12;
b_sign0 = 4'd12; b_sign1 = 4'd12; b_sign2 = 4'd9; b_sign3 = 4'd10;
@(posedge clk_i);
a_mant0 = 8'd244; a_mant1 = 8'd134; a_mant2 = 8'd101; a_mant3 = 8'd97;
b_mant0 = 8'd18; b_mant1 = 8'd150; b_mant2 = 8'd158; b_mant3 = 8'd85;
a_exp0 = 10'd765; a_exp1 = 10'd190; a_exp2 = 10'd816; a_exp3 = 10'd962;
b_exp0 = 10'd461; b_exp1 = 10'd882; b_exp2 = 10'd258; b_exp3 = 10'd92;
a_sign0 = 4'd16; a_sign1 = 4'd16; a_sign2 = 4'd16; a_sign3 = 4'd0;
b_sign0 = 4'd16; b_sign1 = 4'd6; b_sign2 = 4'd14; b_sign3 = 4'd11;
@(posedge clk_i);
a_mant0 = 8'd110; a_mant1 = 8'd34; a_mant2 = 8'd144; a_mant3 = 8'd183;
b_mant0 = 8'd249; b_mant1 = 8'd163; b_mant2 = 8'd250; b_mant3 = 8'd0;
a_exp0 = 10'd1; a_exp1 = 10'd351; a_exp2 = 10'd498; a_exp3 = 10'd411;
b_exp0 = 10'd837; b_exp1 = 10'd164; b_exp2 = 10'd324; b_exp3 = 10'd516;
a_sign0 = 4'd3; a_sign1 = 4'd5; a_sign2 = 4'd1; a_sign3 = 4'd5;
b_sign0 = 4'd12; b_sign1 = 4'd9; b_sign2 = 4'd8; b_sign3 = 4'd12;
@(posedge clk_i);
shared_exps0 = 8'd136;
shared_exps1 = 8'd119;
a_mant0 = 8'd167; a_mant1 = 8'd93; a_mant2 = 8'd214; a_mant3 = 8'd105;
b_mant0 = 8'd110; b_mant1 = 8'd190; b_mant2 = 8'd150; b_mant3 = 8'd1;
a_exp0 = 10'd150; a_exp1 = 10'd889; a_exp2 = 10'd922; a_exp3 = 10'd1008;
b_exp0 = 10'd642; b_exp1 = 10'd377; b_exp2 = 10'd215; b_exp3 = 10'd942;
a_sign0 = 4'd5; a_sign1 = 4'd0; a_sign2 = 4'd10; a_sign3 = 4'd5;
b_sign0 = 4'd14; b_sign1 = 4'd5; b_sign2 = 4'd7; b_sign3 = 4'd6;
@(posedge clk_i);
a_mant0 = 8'd77; a_mant1 = 8'd212; a_mant2 = 8'd183; a_mant3 = 8'd201;
b_mant0 = 8'd60; b_mant1 = 8'd175; b_mant2 = 8'd178; b_mant3 = 8'd4;
a_exp0 = 10'd142; a_exp1 = 10'd821; a_exp2 = 10'd619; a_exp3 = 10'd402;
b_exp0 = 10'd628; b_exp1 = 10'd68; b_exp2 = 10'd998; b_exp3 = 10'd878;
a_sign0 = 4'd3; a_sign1 = 4'd7; a_sign2 = 4'd3; a_sign3 = 4'd11;
b_sign0 = 4'd3; b_sign1 = 4'd12; b_sign2 = 4'd1; b_sign3 = 4'd14;
@(posedge clk_i);
a_mant0 = 8'd101; a_mant1 = 8'd35; a_mant2 = 8'd230; a_mant3 = 8'd51;
b_mant0 = 8'd189; b_mant1 = 8'd161; b_mant2 = 8'd47; b_mant3 = 8'd154;
a_exp0 = 10'd979; a_exp1 = 10'd223; a_exp2 = 10'd258; a_exp3 = 10'd108;
b_exp0 = 10'd391; b_exp1 = 10'd259; b_exp2 = 10'd178; b_exp3 = 10'd405;
a_sign0 = 4'd3; a_sign1 = 4'd1; a_sign2 = 4'd0; a_sign3 = 4'd11;
b_sign0 = 4'd7; b_sign1 = 4'd13; b_sign2 = 4'd13; b_sign3 = 4'd3;
@(posedge clk_i);
a_mant0 = 8'd199; a_mant1 = 8'd197; a_mant2 = 8'd128; a_mant3 = 8'd93;
b_mant0 = 8'd50; b_mant1 = 8'd229; b_mant2 = 8'd245; b_mant3 = 8'd69;
a_exp0 = 10'd868; a_exp1 = 10'd817; a_exp2 = 10'd416; a_exp3 = 10'd322;
b_exp0 = 10'd866; b_exp1 = 10'd208; b_exp2 = 10'd85; b_exp3 = 10'd480;
a_sign0 = 4'd15; a_sign1 = 4'd6; a_sign2 = 4'd0; a_sign3 = 4'd10;
b_sign0 = 4'd3; b_sign1 = 4'd15; b_sign2 = 4'd4; b_sign3 = 4'd4;
@(posedge clk_i);
a_mant0 = 8'd239; a_mant1 = 8'd143; a_mant2 = 8'd245; a_mant3 = 8'd94;
b_mant0 = 8'd70; b_mant1 = 8'd234; b_mant2 = 8'd228; b_mant3 = 8'd230;
a_exp0 = 10'd286; a_exp1 = 10'd822; a_exp2 = 10'd632; a_exp3 = 10'd2;
b_exp0 = 10'd458; b_exp1 = 10'd886; b_exp2 = 10'd262; b_exp3 = 10'd303;
a_sign0 = 4'd9; a_sign1 = 4'd12; a_sign2 = 4'd13; a_sign3 = 4'd5;
b_sign0 = 4'd8; b_sign1 = 4'd6; b_sign2 = 4'd2; b_sign3 = 4'd11;
@(posedge clk_i);
a_mant0 = 8'd93; a_mant1 = 8'd96; a_mant2 = 8'd227; a_mant3 = 8'd115;
b_mant0 = 8'd50; b_mant1 = 8'd98; b_mant2 = 8'd35; b_mant3 = 8'd234;
a_exp0 = 10'd21; a_exp1 = 10'd738; a_exp2 = 10'd759; a_exp3 = 10'd778;
b_exp0 = 10'd787; b_exp1 = 10'd324; b_exp2 = 10'd782; b_exp3 = 10'd13;
a_sign0 = 4'd16; a_sign1 = 4'd0; a_sign2 = 4'd15; a_sign3 = 4'd5;
b_sign0 = 4'd2; b_sign1 = 4'd13; b_sign2 = 4'd13; b_sign3 = 4'd7;
@(posedge clk_i);
a_mant0 = 8'd255; a_mant1 = 8'd160; a_mant2 = 8'd237; a_mant3 = 8'd113;
b_mant0 = 8'd82; b_mant1 = 8'd237; b_mant2 = 8'd111; b_mant3 = 8'd80;
a_exp0 = 10'd908; a_exp1 = 10'd238; a_exp2 = 10'd280; a_exp3 = 10'd364;
b_exp0 = 10'd435; b_exp1 = 10'd840; b_exp2 = 10'd130; b_exp3 = 10'd425;
a_sign0 = 4'd15; a_sign1 = 4'd14; a_sign2 = 4'd13; a_sign3 = 4'd10;
b_sign0 = 4'd9; b_sign1 = 4'd11; b_sign2 = 4'd0; b_sign3 = 4'd8;
@(posedge clk_i);
a_mant0 = 8'd167; a_mant1 = 8'd160; a_mant2 = 8'd50; a_mant3 = 8'd81;
b_mant0 = 8'd188; b_mant1 = 8'd233; b_mant2 = 8'd218; b_mant3 = 8'd156;
a_exp0 = 10'd941; a_exp1 = 10'd929; a_exp2 = 10'd65; a_exp3 = 10'd943;
b_exp0 = 10'd102; b_exp1 = 10'd93; b_exp2 = 10'd147; b_exp3 = 10'd886;
a_sign0 = 4'd9; a_sign1 = 4'd9; a_sign2 = 4'd6; a_sign3 = 4'd15;
b_sign0 = 4'd4; b_sign1 = 4'd7; b_sign2 = 4'd0; b_sign3 = 4'd4;
@(posedge clk_i);
shared_exps0 = 8'd128;
shared_exps1 = 8'd132;
a_mant0 = 8'd21; a_mant1 = 8'd86; a_mant2 = 8'd157; a_mant3 = 8'd5;
b_mant0 = 8'd187; b_mant1 = 8'd3; b_mant2 = 8'd236; b_mant3 = 8'd59;
a_exp0 = 10'd723; a_exp1 = 10'd572; a_exp2 = 10'd209; a_exp3 = 10'd905;
b_exp0 = 10'd470; b_exp1 = 10'd362; b_exp2 = 10'd197; b_exp3 = 10'd195;
a_sign0 = 4'd4; a_sign1 = 4'd2; a_sign2 = 4'd6; a_sign3 = 4'd8;
b_sign0 = 4'd0; b_sign1 = 4'd14; b_sign2 = 4'd7; b_sign3 = 4'd16;
@(posedge clk_i);
a_mant0 = 8'd140; a_mant1 = 8'd140; a_mant2 = 8'd38; a_mant3 = 8'd149;
b_mant0 = 8'd252; b_mant1 = 8'd102; b_mant2 = 8'd119; b_mant3 = 8'd24;
a_exp0 = 10'd203; a_exp1 = 10'd283; a_exp2 = 10'd169; a_exp3 = 10'd222;
b_exp0 = 10'd827; b_exp1 = 10'd28; b_exp2 = 10'd97; b_exp3 = 10'd344;
a_sign0 = 4'd12; a_sign1 = 4'd8; a_sign2 = 4'd8; a_sign3 = 4'd2;
b_sign0 = 4'd14; b_sign1 = 4'd10; b_sign2 = 4'd2; b_sign3 = 4'd12;
@(posedge clk_i);
a_mant0 = 8'd231; a_mant1 = 8'd195; a_mant2 = 8'd161; a_mant3 = 8'd138;
b_mant0 = 8'd128; b_mant1 = 8'd254; b_mant2 = 8'd116; b_mant3 = 8'd129;
a_exp0 = 10'd422; a_exp1 = 10'd797; a_exp2 = 10'd309; a_exp3 = 10'd268;
b_exp0 = 10'd593; b_exp1 = 10'd631; b_exp2 = 10'd467; b_exp3 = 10'd341;
a_sign0 = 4'd12; a_sign1 = 4'd7; a_sign2 = 4'd13; a_sign3 = 4'd9;
b_sign0 = 4'd6; b_sign1 = 4'd6; b_sign2 = 4'd15; b_sign3 = 4'd14;
@(posedge clk_i);
a_mant0 = 8'd73; a_mant1 = 8'd51; a_mant2 = 8'd78; a_mant3 = 8'd58;
b_mant0 = 8'd186; b_mant1 = 8'd80; b_mant2 = 8'd209; b_mant3 = 8'd17;
a_exp0 = 10'd130; a_exp1 = 10'd14; a_exp2 = 10'd299; a_exp3 = 10'd421;
b_exp0 = 10'd617; b_exp1 = 10'd123; b_exp2 = 10'd540; b_exp3 = 10'd978;
a_sign0 = 4'd0; a_sign1 = 4'd8; a_sign2 = 4'd8; a_sign3 = 4'd14;
b_sign0 = 4'd10; b_sign1 = 4'd16; b_sign2 = 4'd16; b_sign3 = 4'd9;
@(posedge clk_i);
a_mant0 = 8'd107; a_mant1 = 8'd17; a_mant2 = 8'd11; a_mant3 = 8'd47;
b_mant0 = 8'd7; b_mant1 = 8'd172; b_mant2 = 8'd72; b_mant3 = 8'd136;
a_exp0 = 10'd368; a_exp1 = 10'd673; a_exp2 = 10'd797; a_exp3 = 10'd811;
b_exp0 = 10'd629; b_exp1 = 10'd950; b_exp2 = 10'd768; b_exp3 = 10'd316;
a_sign0 = 4'd12; a_sign1 = 4'd7; a_sign2 = 4'd9; a_sign3 = 4'd14;
b_sign0 = 4'd7; b_sign1 = 4'd13; b_sign2 = 4'd15; b_sign3 = 4'd9;
@(posedge clk_i);
a_mant0 = 8'd23; a_mant1 = 8'd153; a_mant2 = 8'd31; a_mant3 = 8'd3;
b_mant0 = 8'd158; b_mant1 = 8'd109; b_mant2 = 8'd80; b_mant3 = 8'd28;
a_exp0 = 10'd216; a_exp1 = 10'd758; a_exp2 = 10'd717; a_exp3 = 10'd129;
b_exp0 = 10'd167; b_exp1 = 10'd324; b_exp2 = 10'd62; b_exp3 = 10'd685;
a_sign0 = 4'd13; a_sign1 = 4'd4; a_sign2 = 4'd14; a_sign3 = 4'd14;
b_sign0 = 4'd1; b_sign1 = 4'd14; b_sign2 = 4'd7; b_sign3 = 4'd7;
@(posedge clk_i);
a_mant0 = 8'd237; a_mant1 = 8'd42; a_mant2 = 8'd225; a_mant3 = 8'd15;
b_mant0 = 8'd38; b_mant1 = 8'd219; b_mant2 = 8'd204; b_mant3 = 8'd115;
a_exp0 = 10'd715; a_exp1 = 10'd925; a_exp2 = 10'd973; a_exp3 = 10'd810;
b_exp0 = 10'd907; b_exp1 = 10'd904; b_exp2 = 10'd59; b_exp3 = 10'd261;
a_sign0 = 4'd4; a_sign1 = 4'd2; a_sign2 = 4'd10; a_sign3 = 4'd4;
b_sign0 = 4'd7; b_sign1 = 4'd0; b_sign2 = 4'd3; b_sign3 = 4'd15;
@(posedge clk_i);
a_mant0 = 8'd48; a_mant1 = 8'd229; a_mant2 = 8'd215; a_mant3 = 8'd28;
b_mant0 = 8'd45; b_mant1 = 8'd176; b_mant2 = 8'd45; b_mant3 = 8'd43;
a_exp0 = 10'd422; a_exp1 = 10'd219; a_exp2 = 10'd66; a_exp3 = 10'd634;
b_exp0 = 10'd953; b_exp1 = 10'd886; b_exp2 = 10'd142; b_exp3 = 10'd358;
a_sign0 = 4'd14; a_sign1 = 4'd5; a_sign2 = 4'd11; a_sign3 = 4'd7;
b_sign0 = 4'd5; b_sign1 = 4'd5; b_sign2 = 4'd16; b_sign3 = 4'd11;
@(posedge clk_i);
shared_exps0 = 8'd147;
shared_exps1 = 8'd124;
a_mant0 = 8'd113; a_mant1 = 8'd69; a_mant2 = 8'd82; a_mant3 = 8'd246;
b_mant0 = 8'd100; b_mant1 = 8'd221; b_mant2 = 8'd73; b_mant3 = 8'd232;
a_exp0 = 10'd971; a_exp1 = 10'd818; a_exp2 = 10'd395; a_exp3 = 10'd863;
b_exp0 = 10'd790; b_exp1 = 10'd126; b_exp2 = 10'd722; b_exp3 = 10'd388;
a_sign0 = 4'd9; a_sign1 = 4'd9; a_sign2 = 4'd7; a_sign3 = 4'd0;
b_sign0 = 4'd7; b_sign1 = 4'd6; b_sign2 = 4'd16; b_sign3 = 4'd8;
@(posedge clk_i);
a_mant0 = 8'd174; a_mant1 = 8'd130; a_mant2 = 8'd233; a_mant3 = 8'd40;
b_mant0 = 8'd46; b_mant1 = 8'd124; b_mant2 = 8'd190; b_mant3 = 8'd247;
a_exp0 = 10'd373; a_exp1 = 10'd603; a_exp2 = 10'd893; a_exp3 = 10'd764;
b_exp0 = 10'd378; b_exp1 = 10'd625; b_exp2 = 10'd846; b_exp3 = 10'd699;
a_sign0 = 4'd5; a_sign1 = 4'd8; a_sign2 = 4'd1; a_sign3 = 4'd8;
b_sign0 = 4'd11; b_sign1 = 4'd1; b_sign2 = 4'd16; b_sign3 = 4'd2;
@(posedge clk_i);
a_mant0 = 8'd218; a_mant1 = 8'd111; a_mant2 = 8'd83; a_mant3 = 8'd205;
b_mant0 = 8'd253; b_mant1 = 8'd191; b_mant2 = 8'd124; b_mant3 = 8'd219;
a_exp0 = 10'd639; a_exp1 = 10'd763; a_exp2 = 10'd205; a_exp3 = 10'd1009;
b_exp0 = 10'd649; b_exp1 = 10'd184; b_exp2 = 10'd662; b_exp3 = 10'd434;
a_sign0 = 4'd9; a_sign1 = 4'd0; a_sign2 = 4'd1; a_sign3 = 4'd6;
b_sign0 = 4'd6; b_sign1 = 4'd14; b_sign2 = 4'd15; b_sign3 = 4'd0;
@(posedge clk_i);
a_mant0 = 8'd12; a_mant1 = 8'd176; a_mant2 = 8'd244; a_mant3 = 8'd132;
b_mant0 = 8'd254; b_mant1 = 8'd188; b_mant2 = 8'd127; b_mant3 = 8'd56;
a_exp0 = 10'd225; a_exp1 = 10'd318; a_exp2 = 10'd695; a_exp3 = 10'd107;
b_exp0 = 10'd3; b_exp1 = 10'd191; b_exp2 = 10'd454; b_exp3 = 10'd508;
a_sign0 = 4'd0; a_sign1 = 4'd12; a_sign2 = 4'd9; a_sign3 = 4'd4;
b_sign0 = 4'd14; b_sign1 = 4'd14; b_sign2 = 4'd16; b_sign3 = 4'd6;
@(posedge clk_i);
a_mant0 = 8'd177; a_mant1 = 8'd37; a_mant2 = 8'd140; a_mant3 = 8'd212;
b_mant0 = 8'd124; b_mant1 = 8'd81; b_mant2 = 8'd191; b_mant3 = 8'd113;
a_exp0 = 10'd881; a_exp1 = 10'd608; a_exp2 = 10'd733; a_exp3 = 10'd773;
b_exp0 = 10'd605; b_exp1 = 10'd857; b_exp2 = 10'd671; b_exp3 = 10'd399;
a_sign0 = 4'd11; a_sign1 = 4'd8; a_sign2 = 4'd10; a_sign3 = 4'd10;
b_sign0 = 4'd12; b_sign1 = 4'd11; b_sign2 = 4'd7; b_sign3 = 4'd10;
@(posedge clk_i);
a_mant0 = 8'd200; a_mant1 = 8'd47; a_mant2 = 8'd39; a_mant3 = 8'd82;
b_mant0 = 8'd228; b_mant1 = 8'd246; b_mant2 = 8'd126; b_mant3 = 8'd131;
a_exp0 = 10'd965; a_exp1 = 10'd872; a_exp2 = 10'd54; a_exp3 = 10'd957;
b_exp0 = 10'd22; b_exp1 = 10'd967; b_exp2 = 10'd255; b_exp3 = 10'd423;
a_sign0 = 4'd10; a_sign1 = 4'd6; a_sign2 = 4'd10; a_sign3 = 4'd12;
b_sign0 = 4'd8; b_sign1 = 4'd15; b_sign2 = 4'd12; b_sign3 = 4'd13;
@(posedge clk_i);
a_mant0 = 8'd18; a_mant1 = 8'd116; a_mant2 = 8'd173; a_mant3 = 8'd0;
b_mant0 = 8'd43; b_mant1 = 8'd44; b_mant2 = 8'd167; b_mant3 = 8'd128;
a_exp0 = 10'd974; a_exp1 = 10'd99; a_exp2 = 10'd1010; a_exp3 = 10'd239;
b_exp0 = 10'd71; b_exp1 = 10'd156; b_exp2 = 10'd203; b_exp3 = 10'd901;
a_sign0 = 4'd14; a_sign1 = 4'd9; a_sign2 = 4'd5; a_sign3 = 4'd8;
b_sign0 = 4'd16; b_sign1 = 4'd1; b_sign2 = 4'd7; b_sign3 = 4'd4;
@(posedge clk_i);
a_mant0 = 8'd168; a_mant1 = 8'd133; a_mant2 = 8'd111; a_mant3 = 8'd57;
b_mant0 = 8'd146; b_mant1 = 8'd174; b_mant2 = 8'd48; b_mant3 = 8'd245;
a_exp0 = 10'd38; a_exp1 = 10'd172; a_exp2 = 10'd119; a_exp3 = 10'd460;
b_exp0 = 10'd668; b_exp1 = 10'd415; b_exp2 = 10'd250; b_exp3 = 10'd834;
a_sign0 = 4'd11; a_sign1 = 4'd7; a_sign2 = 4'd9; a_sign3 = 4'd13;
b_sign0 = 4'd8; b_sign1 = 4'd12; b_sign2 = 4'd14; b_sign3 = 4'd16;
@(posedge clk_i);
shared_exps0 = 8'd143;
shared_exps1 = 8'd137;
rstn = 0;
@(posedge clk_i);
rstn = 1;
a_mant0 = 8'd54; a_mant1 = 8'd54; a_mant2 = 8'd159; a_mant3 = 8'd227;
b_mant0 = 8'd2; b_mant1 = 8'd161; b_mant2 = 8'd223; b_mant3 = 8'd79;
a_exp0 = 10'd808; a_exp1 = 10'd436; a_exp2 = 10'd842; a_exp3 = 10'd527;
b_exp0 = 10'd363; b_exp1 = 10'd680; b_exp2 = 10'd363; b_exp3 = 10'd825;
a_sign0 = 4'd10; a_sign1 = 4'd2; a_sign2 = 4'd10; a_sign3 = 4'd7;
b_sign0 = 4'd6; b_sign1 = 4'd6; b_sign2 = 4'd4; b_sign3 = 4'd1;
@(posedge clk_i);
a_mant0 = 8'd62; a_mant1 = 8'd210; a_mant2 = 8'd220; a_mant3 = 8'd172;
b_mant0 = 8'd240; b_mant1 = 8'd135; b_mant2 = 8'd19; b_mant3 = 8'd79;
a_exp0 = 10'd530; a_exp1 = 10'd861; a_exp2 = 10'd973; a_exp3 = 10'd155;
b_exp0 = 10'd796; b_exp1 = 10'd588; b_exp2 = 10'd847; b_exp3 = 10'd704;
a_sign0 = 4'd6; a_sign1 = 4'd8; a_sign2 = 4'd13; a_sign3 = 4'd10;
b_sign0 = 4'd16; b_sign1 = 4'd12; b_sign2 = 4'd1; b_sign3 = 4'd5;
@(posedge clk_i);
a_mant0 = 8'd36; a_mant1 = 8'd176; a_mant2 = 8'd53; a_mant3 = 8'd21;
b_mant0 = 8'd231; b_mant1 = 8'd87; b_mant2 = 8'd52; b_mant3 = 8'd176;
a_exp0 = 10'd384; a_exp1 = 10'd469; a_exp2 = 10'd558; a_exp3 = 10'd652;
b_exp0 = 10'd264; b_exp1 = 10'd506; b_exp2 = 10'd270; b_exp3 = 10'd899;
a_sign0 = 4'd12; a_sign1 = 4'd3; a_sign2 = 4'd6; a_sign3 = 4'd2;
b_sign0 = 4'd12; b_sign1 = 4'd0; b_sign2 = 4'd1; b_sign3 = 4'd4;
@(posedge clk_i);
a_mant0 = 8'd154; a_mant1 = 8'd38; a_mant2 = 8'd164; a_mant3 = 8'd14;
b_mant0 = 8'd215; b_mant1 = 8'd45; b_mant2 = 8'd249; b_mant3 = 8'd37;
a_exp0 = 10'd346; a_exp1 = 10'd951; a_exp2 = 10'd595; a_exp3 = 10'd979;
b_exp0 = 10'd794; b_exp1 = 10'd834; b_exp2 = 10'd984; b_exp3 = 10'd25;
a_sign0 = 4'd15; a_sign1 = 4'd11; a_sign2 = 4'd14; a_sign3 = 4'd13;
b_sign0 = 4'd13; b_sign1 = 4'd6; b_sign2 = 4'd5; b_sign3 = 4'd4;
@(posedge clk_i);
a_mant0 = 8'd18; a_mant1 = 8'd118; a_mant2 = 8'd249; a_mant3 = 8'd193;
b_mant0 = 8'd144; b_mant1 = 8'd134; b_mant2 = 8'd138; b_mant3 = 8'd83;
a_exp0 = 10'd550; a_exp1 = 10'd326; a_exp2 = 10'd429; a_exp3 = 10'd24;
b_exp0 = 10'd331; b_exp1 = 10'd316; b_exp2 = 10'd477; b_exp3 = 10'd856;
a_sign0 = 4'd0; a_sign1 = 4'd5; a_sign2 = 4'd12; a_sign3 = 4'd6;
b_sign0 = 4'd12; b_sign1 = 4'd6; b_sign2 = 4'd13; b_sign3 = 4'd10;
@(posedge clk_i);
a_mant0 = 8'd36; a_mant1 = 8'd151; a_mant2 = 8'd248; a_mant3 = 8'd223;
b_mant0 = 8'd144; b_mant1 = 8'd170; b_mant2 = 8'd184; b_mant3 = 8'd175;
a_exp0 = 10'd985; a_exp1 = 10'd143; a_exp2 = 10'd543; a_exp3 = 10'd183;
b_exp0 = 10'd985; b_exp1 = 10'd472; b_exp2 = 10'd17; b_exp3 = 10'd690;
a_sign0 = 4'd16; a_sign1 = 4'd4; a_sign2 = 4'd3; a_sign3 = 4'd11;
b_sign0 = 4'd7; b_sign1 = 4'd10; b_sign2 = 4'd10; b_sign3 = 4'd3;
@(posedge clk_i);
a_mant0 = 8'd245; a_mant1 = 8'd81; a_mant2 = 8'd28; a_mant3 = 8'd121;
b_mant0 = 8'd34; b_mant1 = 8'd92; b_mant2 = 8'd190; b_mant3 = 8'd29;
a_exp0 = 10'd510; a_exp1 = 10'd296; a_exp2 = 10'd106; a_exp3 = 10'd872;
b_exp0 = 10'd300; b_exp1 = 10'd69; b_exp2 = 10'd933; b_exp3 = 10'd681;
a_sign0 = 4'd14; a_sign1 = 4'd9; a_sign2 = 4'd7; a_sign3 = 4'd12;
b_sign0 = 4'd4; b_sign1 = 4'd11; b_sign2 = 4'd2; b_sign3 = 4'd7;
@(posedge clk_i);
shared_exps0 = 8'd151;
shared_exps1 = 8'd141;
a_mant0 = 8'd133; a_mant1 = 8'd124; a_mant2 = 8'd135; a_mant3 = 8'd101;
b_mant0 = 8'd221; b_mant1 = 8'd30; b_mant2 = 8'd218; b_mant3 = 8'd79;
a_exp0 = 10'd479; a_exp1 = 10'd983; a_exp2 = 10'd301; a_exp3 = 10'd456;
b_exp0 = 10'd832; b_exp1 = 10'd215; b_exp2 = 10'd597; b_exp3 = 10'd370;
a_sign0 = 4'd3; a_sign1 = 4'd16; a_sign2 = 4'd7; a_sign3 = 4'd14;
b_sign0 = 4'd2; b_sign1 = 4'd3; b_sign2 = 4'd8; b_sign3 = 4'd16;
@(posedge clk_i);
a_mant0 = 8'd252; a_mant1 = 8'd189; a_mant2 = 8'd67; a_mant3 = 8'd185;
b_mant0 = 8'd123; b_mant1 = 8'd140; b_mant2 = 8'd195; b_mant3 = 8'd18;
a_exp0 = 10'd549; a_exp1 = 10'd823; a_exp2 = 10'd344; a_exp3 = 10'd641;
b_exp0 = 10'd951; b_exp1 = 10'd673; b_exp2 = 10'd49; b_exp3 = 10'd460;
a_sign0 = 4'd7; a_sign1 = 4'd2; a_sign2 = 4'd11; a_sign3 = 4'd9;
b_sign0 = 4'd12; b_sign1 = 4'd7; b_sign2 = 4'd7; b_sign3 = 4'd13;
@(posedge clk_i);
a_mant0 = 8'd191; a_mant1 = 8'd135; a_mant2 = 8'd28; a_mant3 = 8'd209;
b_mant0 = 8'd217; b_mant1 = 8'd235; b_mant2 = 8'd1; b_mant3 = 8'd214;
a_exp0 = 10'd397; a_exp1 = 10'd363; a_exp2 = 10'd285; a_exp3 = 10'd794;
b_exp0 = 10'd593; b_exp1 = 10'd65; b_exp2 = 10'd675; b_exp3 = 10'd284;
a_sign0 = 4'd12; a_sign1 = 4'd1; a_sign2 = 4'd14; a_sign3 = 4'd7;
b_sign0 = 4'd13; b_sign1 = 4'd4; b_sign2 = 4'd15; b_sign3 = 4'd4;
@(posedge clk_i);
a_mant0 = 8'd68; a_mant1 = 8'd60; a_mant2 = 8'd16; a_mant3 = 8'd199;
b_mant0 = 8'd201; b_mant1 = 8'd194; b_mant2 = 8'd35; b_mant3 = 8'd22;
a_exp0 = 10'd511; a_exp1 = 10'd1016; a_exp2 = 10'd178; a_exp3 = 10'd873;
b_exp0 = 10'd885; b_exp1 = 10'd760; b_exp2 = 10'd801; b_exp3 = 10'd417;
a_sign0 = 4'd9; a_sign1 = 4'd1; a_sign2 = 4'd5; a_sign3 = 4'd1;
b_sign0 = 4'd15; b_sign1 = 4'd14; b_sign2 = 4'd15; b_sign3 = 4'd8;
@(posedge clk_i);
a_mant0 = 8'd3; a_mant1 = 8'd203; a_mant2 = 8'd135; a_mant3 = 8'd216;
b_mant0 = 8'd66; b_mant1 = 8'd91; b_mant2 = 8'd95; b_mant3 = 8'd108;
a_exp0 = 10'd14; a_exp1 = 10'd383; a_exp2 = 10'd897; a_exp3 = 10'd36;
b_exp0 = 10'd749; b_exp1 = 10'd963; b_exp2 = 10'd87; b_exp3 = 10'd25;
a_sign0 = 4'd0; a_sign1 = 4'd0; a_sign2 = 4'd10; a_sign3 = 4'd5;
b_sign0 = 4'd5; b_sign1 = 4'd9; b_sign2 = 4'd8; b_sign3 = 4'd16;
@(posedge clk_i);
a_mant0 = 8'd111; a_mant1 = 8'd51; a_mant2 = 8'd91; a_mant3 = 8'd16;
b_mant0 = 8'd207; b_mant1 = 8'd171; b_mant2 = 8'd60; b_mant3 = 8'd85;
a_exp0 = 10'd235; a_exp1 = 10'd744; a_exp2 = 10'd648; a_exp3 = 10'd247;
b_exp0 = 10'd984; b_exp1 = 10'd25; b_exp2 = 10'd469; b_exp3 = 10'd336;
a_sign0 = 4'd3; a_sign1 = 4'd11; a_sign2 = 4'd1; a_sign3 = 4'd0;
b_sign0 = 4'd1; b_sign1 = 4'd15; b_sign2 = 4'd15; b_sign3 = 4'd7;
@(posedge clk_i);
a_mant0 = 8'd236; a_mant1 = 8'd89; a_mant2 = 8'd213; a_mant3 = 8'd211;
b_mant0 = 8'd64; b_mant1 = 8'd117; b_mant2 = 8'd118; b_mant3 = 8'd43;
a_exp0 = 10'd579; a_exp1 = 10'd559; a_exp2 = 10'd181; a_exp3 = 10'd694;
b_exp0 = 10'd505; b_exp1 = 10'd546; b_exp2 = 10'd846; b_exp3 = 10'd478;
a_sign0 = 4'd8; a_sign1 = 4'd0; a_sign2 = 4'd14; a_sign3 = 4'd3;
b_sign0 = 4'd13; b_sign1 = 4'd13; b_sign2 = 4'd10; b_sign3 = 4'd3;
@(posedge clk_i);
a_mant0 = 8'd7; a_mant1 = 8'd40; a_mant2 = 8'd152; a_mant3 = 8'd140;
b_mant0 = 8'd99; b_mant1 = 8'd50; b_mant2 = 8'd150; b_mant3 = 8'd211;
a_exp0 = 10'd857; a_exp1 = 10'd883; a_exp2 = 10'd885; a_exp3 = 10'd370;
b_exp0 = 10'd84; b_exp1 = 10'd812; b_exp2 = 10'd209; b_exp3 = 10'd546;
a_sign0 = 4'd9; a_sign1 = 4'd10; a_sign2 = 4'd3; a_sign3 = 4'd9;
b_sign0 = 4'd0; b_sign1 = 4'd15; b_sign2 = 4'd11; b_sign3 = 4'd8;
@(posedge clk_i);
shared_exps0 = 8'd128;
shared_exps1 = 8'd118;
a_mant0 = 8'd216; a_mant1 = 8'd188; a_mant2 = 8'd212; a_mant3 = 8'd77;
b_mant0 = 8'd52; b_mant1 = 8'd161; b_mant2 = 8'd244; b_mant3 = 8'd18;
a_exp0 = 10'd742; a_exp1 = 10'd125; a_exp2 = 10'd928; a_exp3 = 10'd631;
b_exp0 = 10'd441; b_exp1 = 10'd110; b_exp2 = 10'd284; b_exp3 = 10'd836;
a_sign0 = 4'd14; a_sign1 = 4'd0; a_sign2 = 4'd9; a_sign3 = 4'd15;
b_sign0 = 4'd14; b_sign1 = 4'd4; b_sign2 = 4'd13; b_sign3 = 4'd13;
@(posedge clk_i);
a_mant0 = 8'd100; a_mant1 = 8'd107; a_mant2 = 8'd81; a_mant3 = 8'd226;
b_mant0 = 8'd237; b_mant1 = 8'd108; b_mant2 = 8'd200; b_mant3 = 8'd16;
a_exp0 = 10'd988; a_exp1 = 10'd818; a_exp2 = 10'd881; a_exp3 = 10'd689;
b_exp0 = 10'd464; b_exp1 = 10'd534; b_exp2 = 10'd214; b_exp3 = 10'd1013;
a_sign0 = 4'd4; a_sign1 = 4'd12; a_sign2 = 4'd1; a_sign3 = 4'd15;
b_sign0 = 4'd8; b_sign1 = 4'd1; b_sign2 = 4'd16; b_sign3 = 4'd6;
@(posedge clk_i);
a_mant0 = 8'd158; a_mant1 = 8'd183; a_mant2 = 8'd170; a_mant3 = 8'd127;
b_mant0 = 8'd116; b_mant1 = 8'd84; b_mant2 = 8'd42; b_mant3 = 8'd231;
a_exp0 = 10'd661; a_exp1 = 10'd952; a_exp2 = 10'd23; a_exp3 = 10'd79;
b_exp0 = 10'd101; b_exp1 = 10'd682; b_exp2 = 10'd637; b_exp3 = 10'd969;
a_sign0 = 4'd4; a_sign1 = 4'd7; a_sign2 = 4'd4; a_sign3 = 4'd4;
b_sign0 = 4'd16; b_sign1 = 4'd2; b_sign2 = 4'd5; b_sign3 = 4'd14;
@(posedge clk_i);
a_mant0 = 8'd99; a_mant1 = 8'd236; a_mant2 = 8'd238; a_mant3 = 8'd221;
b_mant0 = 8'd67; b_mant1 = 8'd18; b_mant2 = 8'd68; b_mant3 = 8'd44;
a_exp0 = 10'd432; a_exp1 = 10'd138; a_exp2 = 10'd888; a_exp3 = 10'd983;
b_exp0 = 10'd651; b_exp1 = 10'd31; b_exp2 = 10'd899; b_exp3 = 10'd834;
a_sign0 = 4'd1; a_sign1 = 4'd13; a_sign2 = 4'd14; a_sign3 = 4'd4;
b_sign0 = 4'd13; b_sign1 = 4'd9; b_sign2 = 4'd13; b_sign3 = 4'd0;
@(posedge clk_i);
a_mant0 = 8'd24; a_mant1 = 8'd240; a_mant2 = 8'd134; a_mant3 = 8'd54;
b_mant0 = 8'd38; b_mant1 = 8'd31; b_mant2 = 8'd136; b_mant3 = 8'd13;
a_exp0 = 10'd461; a_exp1 = 10'd169; a_exp2 = 10'd963; a_exp3 = 10'd1006;
b_exp0 = 10'd929; b_exp1 = 10'd608; b_exp2 = 10'd987; b_exp3 = 10'd797;
a_sign0 = 4'd7; a_sign1 = 4'd13; a_sign2 = 4'd14; a_sign3 = 4'd7;
b_sign0 = 4'd11; b_sign1 = 4'd12; b_sign2 = 4'd3; b_sign3 = 4'd4;
@(posedge clk_i);
a_mant0 = 8'd95; a_mant1 = 8'd34; a_mant2 = 8'd137; a_mant3 = 8'd174;
b_mant0 = 8'd161; b_mant1 = 8'd113; b_mant2 = 8'd59; b_mant3 = 8'd233;
a_exp0 = 10'd10; a_exp1 = 10'd340; a_exp2 = 10'd206; a_exp3 = 10'd345;
b_exp0 = 10'd721; b_exp1 = 10'd248; b_exp2 = 10'd233; b_exp3 = 10'd300;
a_sign0 = 4'd6; a_sign1 = 4'd0; a_sign2 = 4'd6; a_sign3 = 4'd14;
b_sign0 = 4'd9; b_sign1 = 4'd10; b_sign2 = 4'd7; b_sign3 = 4'd2;
@(posedge clk_i);
a_mant0 = 8'd209; a_mant1 = 8'd146; a_mant2 = 8'd112; a_mant3 = 8'd120;
b_mant0 = 8'd179; b_mant1 = 8'd61; b_mant2 = 8'd206; b_mant3 = 8'd177;
a_exp0 = 10'd665; a_exp1 = 10'd23; a_exp2 = 10'd956; a_exp3 = 10'd11;
b_exp0 = 10'd988; b_exp1 = 10'd294; b_exp2 = 10'd260; b_exp3 = 10'd617;
a_sign0 = 4'd10; a_sign1 = 4'd2; a_sign2 = 4'd10; a_sign3 = 4'd9;
b_sign0 = 4'd9; b_sign1 = 4'd1; b_sign2 = 4'd0; b_sign3 = 4'd8;
@(posedge clk_i);
a_mant0 = 8'd103; a_mant1 = 8'd233; a_mant2 = 8'd255; a_mant3 = 8'd231;
b_mant0 = 8'd251; b_mant1 = 8'd133; b_mant2 = 8'd81; b_mant3 = 8'd115;
a_exp0 = 10'd927; a_exp1 = 10'd421; a_exp2 = 10'd379; a_exp3 = 10'd305;
b_exp0 = 10'd123; b_exp1 = 10'd437; b_exp2 = 10'd462; b_exp3 = 10'd888;
a_sign0 = 4'd1; a_sign1 = 4'd5; a_sign2 = 4'd14; a_sign3 = 4'd16;
b_sign0 = 4'd16; b_sign1 = 4'd3; b_sign2 = 4'd12; b_sign3 = 4'd1;
@(posedge clk_i);
shared_exps0 = 8'd126;
shared_exps1 = 8'd95;
a_mant0 = 8'd10; a_mant1 = 8'd60; a_mant2 = 8'd215; a_mant3 = 8'd242;
b_mant0 = 8'd201; b_mant1 = 8'd202; b_mant2 = 8'd54; b_mant3 = 8'd181;
a_exp0 = 10'd765; a_exp1 = 10'd69; a_exp2 = 10'd314; a_exp3 = 10'd439;
b_exp0 = 10'd867; b_exp1 = 10'd664; b_exp2 = 10'd285; b_exp3 = 10'd238;
a_sign0 = 4'd14; a_sign1 = 4'd10; a_sign2 = 4'd4; a_sign3 = 4'd14;
b_sign0 = 4'd5; b_sign1 = 4'd11; b_sign2 = 4'd6; b_sign3 = 4'd6;
@(posedge clk_i);
a_mant0 = 8'd118; a_mant1 = 8'd248; a_mant2 = 8'd124; a_mant3 = 8'd160;
b_mant0 = 8'd147; b_mant1 = 8'd168; b_mant2 = 8'd216; b_mant3 = 8'd179;
a_exp0 = 10'd737; a_exp1 = 10'd905; a_exp2 = 10'd651; a_exp3 = 10'd216;
b_exp0 = 10'd646; b_exp1 = 10'd193; b_exp2 = 10'd491; b_exp3 = 10'd870;
a_sign0 = 4'd3; a_sign1 = 4'd5; a_sign2 = 4'd15; a_sign3 = 4'd13;
b_sign0 = 4'd0; b_sign1 = 4'd9; b_sign2 = 4'd0; b_sign3 = 4'd5;
@(posedge clk_i);
a_mant0 = 8'd181; a_mant1 = 8'd108; a_mant2 = 8'd42; a_mant3 = 8'd110;
b_mant0 = 8'd111; b_mant1 = 8'd66; b_mant2 = 8'd176; b_mant3 = 8'd231;
a_exp0 = 10'd84; a_exp1 = 10'd326; a_exp2 = 10'd210; a_exp3 = 10'd25;
b_exp0 = 10'd76; b_exp1 = 10'd817; b_exp2 = 10'd429; b_exp3 = 10'd323;
a_sign0 = 4'd13; a_sign1 = 4'd8; a_sign2 = 4'd0; a_sign3 = 4'd16;
b_sign0 = 4'd11; b_sign1 = 4'd11; b_sign2 = 4'd6; b_sign3 = 4'd4;
@(posedge clk_i);
a_mant0 = 8'd149; a_mant1 = 8'd23; a_mant2 = 8'd82; a_mant3 = 8'd240;
b_mant0 = 8'd39; b_mant1 = 8'd237; b_mant2 = 8'd239; b_mant3 = 8'd49;
a_exp0 = 10'd751; a_exp1 = 10'd600; a_exp2 = 10'd787; a_exp3 = 10'd637;
b_exp0 = 10'd847; b_exp1 = 10'd819; b_exp2 = 10'd142; b_exp3 = 10'd264;
a_sign0 = 4'd15; a_sign1 = 4'd12; a_sign2 = 4'd9; a_sign3 = 4'd12;
b_sign0 = 4'd8; b_sign1 = 4'd1; b_sign2 = 4'd16; b_sign3 = 4'd14;
@(posedge clk_i);
a_mant0 = 8'd145; a_mant1 = 8'd99; a_mant2 = 8'd220; a_mant3 = 8'd3;
b_mant0 = 8'd89; b_mant1 = 8'd68; b_mant2 = 8'd88; b_mant3 = 8'd69;
a_exp0 = 10'd725; a_exp1 = 10'd319; a_exp2 = 10'd12; a_exp3 = 10'd266;
b_exp0 = 10'd410; b_exp1 = 10'd444; b_exp2 = 10'd234; b_exp3 = 10'd968;
a_sign0 = 4'd4; a_sign1 = 4'd6; a_sign2 = 4'd4; a_sign3 = 4'd6;
b_sign0 = 4'd15; b_sign1 = 4'd10; b_sign2 = 4'd3; b_sign3 = 4'd14;
@(posedge clk_i);
a_mant0 = 8'd35; a_mant1 = 8'd243; a_mant2 = 8'd181; a_mant3 = 8'd84;
b_mant0 = 8'd0; b_mant1 = 8'd166; b_mant2 = 8'd212; b_mant3 = 8'd30;
a_exp0 = 10'd523; a_exp1 = 10'd647; a_exp2 = 10'd736; a_exp3 = 10'd558;
b_exp0 = 10'd769; b_exp1 = 10'd1006; b_exp2 = 10'd980; b_exp3 = 10'd224;
a_sign0 = 4'd15; a_sign1 = 4'd11; a_sign2 = 4'd10; a_sign3 = 4'd16;
b_sign0 = 4'd16; b_sign1 = 4'd15; b_sign2 = 4'd1; b_sign3 = 4'd12;
@(posedge clk_i);
a_mant0 = 8'd9; a_mant1 = 8'd167; a_mant2 = 8'd30; a_mant3 = 8'd127;
b_mant0 = 8'd233; b_mant1 = 8'd15; b_mant2 = 8'd84; b_mant3 = 8'd250;
a_exp0 = 10'd413; a_exp1 = 10'd312; a_exp2 = 10'd975; a_exp3 = 10'd275;
b_exp0 = 10'd161; b_exp1 = 10'd475; b_exp2 = 10'd998; b_exp3 = 10'd989;
a_sign0 = 4'd12; a_sign1 = 4'd13; a_sign2 = 4'd0; a_sign3 = 4'd9;
b_sign0 = 4'd7; b_sign1 = 4'd0; b_sign2 = 4'd9; b_sign3 = 4'd14;
@(posedge clk_i);
a_mant0 = 8'd41; a_mant1 = 8'd211; a_mant2 = 8'd189; a_mant3 = 8'd172;
b_mant0 = 8'd12; b_mant1 = 8'd172; b_mant2 = 8'd18; b_mant3 = 8'd233;
a_exp0 = 10'd866; a_exp1 = 10'd566; a_exp2 = 10'd199; a_exp3 = 10'd241;
b_exp0 = 10'd769; b_exp1 = 10'd842; b_exp2 = 10'd844; b_exp3 = 10'd755;
a_sign0 = 4'd5; a_sign1 = 4'd14; a_sign2 = 4'd6; a_sign3 = 4'd10;
b_sign0 = 4'd2; b_sign1 = 4'd5; b_sign2 = 4'd7; b_sign3 = 4'd6;
@(posedge clk_i);
shared_exps0 = 8'd139;
shared_exps1 = 8'd146;
rstn = 0;
@(posedge clk_i);
rstn = 1;
a_mant0 = 8'd74; a_mant1 = 8'd188; a_mant2 = 8'd108; a_mant3 = 8'd109;
b_mant0 = 8'd203; b_mant1 = 8'd226; b_mant2 = 8'd159; b_mant3 = 8'd118;
a_exp0 = 10'd122; a_exp1 = 10'd465; a_exp2 = 10'd508; a_exp3 = 10'd52;
b_exp0 = 10'd294; b_exp1 = 10'd781; b_exp2 = 10'd287; b_exp3 = 10'd879;
a_sign0 = 4'd14; a_sign1 = 4'd4; a_sign2 = 4'd1; a_sign3 = 4'd10;
b_sign0 = 4'd5; b_sign1 = 4'd5; b_sign2 = 4'd14; b_sign3 = 4'd6;
@(posedge clk_i);
a_mant0 = 8'd107; a_mant1 = 8'd96; a_mant2 = 8'd211; a_mant3 = 8'd246;
b_mant0 = 8'd232; b_mant1 = 8'd182; b_mant2 = 8'd101; b_mant3 = 8'd4;
a_exp0 = 10'd402; a_exp1 = 10'd692; a_exp2 = 10'd493; a_exp3 = 10'd33;
b_exp0 = 10'd784; b_exp1 = 10'd61; b_exp2 = 10'd8; b_exp3 = 10'd549;
a_sign0 = 4'd6; a_sign1 = 4'd14; a_sign2 = 4'd2; a_sign3 = 4'd12;
b_sign0 = 4'd10; b_sign1 = 4'd13; b_sign2 = 4'd15; b_sign3 = 4'd16;
@(posedge clk_i);
a_mant0 = 8'd186; a_mant1 = 8'd169; a_mant2 = 8'd95; a_mant3 = 8'd137;
b_mant0 = 8'd123; b_mant1 = 8'd87; b_mant2 = 8'd55; b_mant3 = 8'd246;
a_exp0 = 10'd841; a_exp1 = 10'd622; a_exp2 = 10'd646; a_exp3 = 10'd450;
b_exp0 = 10'd542; b_exp1 = 10'd841; b_exp2 = 10'd465; b_exp3 = 10'd66;
a_sign0 = 4'd9; a_sign1 = 4'd9; a_sign2 = 4'd13; a_sign3 = 4'd16;
b_sign0 = 4'd4; b_sign1 = 4'd13; b_sign2 = 4'd3; b_sign3 = 4'd12;
@(posedge clk_i);
a_mant0 = 8'd187; a_mant1 = 8'd110; a_mant2 = 8'd253; a_mant3 = 8'd183;
b_mant0 = 8'd36; b_mant1 = 8'd58; b_mant2 = 8'd140; b_mant3 = 8'd120;
a_exp0 = 10'd409; a_exp1 = 10'd628; a_exp2 = 10'd700; a_exp3 = 10'd444;
b_exp0 = 10'd260; b_exp1 = 10'd639; b_exp2 = 10'd964; b_exp3 = 10'd216;
a_sign0 = 4'd0; a_sign1 = 4'd8; a_sign2 = 4'd11; a_sign3 = 4'd16;
b_sign0 = 4'd12; b_sign1 = 4'd4; b_sign2 = 4'd15; b_sign3 = 4'd10;
@(posedge clk_i);
a_mant0 = 8'd3; a_mant1 = 8'd240; a_mant2 = 8'd175; a_mant3 = 8'd153;
b_mant0 = 8'd118; b_mant1 = 8'd12; b_mant2 = 8'd232; b_mant3 = 8'd76;
a_exp0 = 10'd93; a_exp1 = 10'd918; a_exp2 = 10'd838; a_exp3 = 10'd134;
b_exp0 = 10'd972; b_exp1 = 10'd465; b_exp2 = 10'd688; b_exp3 = 10'd864;
a_sign0 = 4'd16; a_sign1 = 4'd4; a_sign2 = 4'd4; a_sign3 = 4'd0;
b_sign0 = 4'd7; b_sign1 = 4'd13; b_sign2 = 4'd2; b_sign3 = 4'd7;
@(posedge clk_i);
a_mant0 = 8'd218; a_mant1 = 8'd95; a_mant2 = 8'd144; a_mant3 = 8'd94;
b_mant0 = 8'd146; b_mant1 = 8'd126; b_mant2 = 8'd5; b_mant3 = 8'd79;
a_exp0 = 10'd887; a_exp1 = 10'd602; a_exp2 = 10'd444; a_exp3 = 10'd201;
b_exp0 = 10'd759; b_exp1 = 10'd277; b_exp2 = 10'd96; b_exp3 = 10'd446;
a_sign0 = 4'd12; a_sign1 = 4'd10; a_sign2 = 4'd10; a_sign3 = 4'd7;
b_sign0 = 4'd14; b_sign1 = 4'd12; b_sign2 = 4'd11; b_sign3 = 4'd8;
@(posedge clk_i);
a_mant0 = 8'd145; a_mant1 = 8'd6; a_mant2 = 8'd235; a_mant3 = 8'd244;
b_mant0 = 8'd54; b_mant1 = 8'd239; b_mant2 = 8'd159; b_mant3 = 8'd25;
a_exp0 = 10'd625; a_exp1 = 10'd526; a_exp2 = 10'd694; a_exp3 = 10'd710;
b_exp0 = 10'd117; b_exp1 = 10'd541; b_exp2 = 10'd285; b_exp3 = 10'd231;
a_sign0 = 4'd1; a_sign1 = 4'd16; a_sign2 = 4'd10; a_sign3 = 4'd10;
b_sign0 = 4'd2; b_sign1 = 4'd16; b_sign2 = 4'd10; b_sign3 = 4'd3;
@(posedge clk_i);
shared_exps0 = 8'd122;
shared_exps1 = 8'd127;
a_mant0 = 8'd192; a_mant1 = 8'd109; a_mant2 = 8'd99; a_mant3 = 8'd141;
b_mant0 = 8'd183; b_mant1 = 8'd54; b_mant2 = 8'd216; b_mant3 = 8'd0;
a_exp0 = 10'd744; a_exp1 = 10'd394; a_exp2 = 10'd994; a_exp3 = 10'd29;
b_exp0 = 10'd744; b_exp1 = 10'd413; b_exp2 = 10'd60; b_exp3 = 10'd762;
a_sign0 = 4'd13; a_sign1 = 4'd1; a_sign2 = 4'd12; a_sign3 = 4'd14;
b_sign0 = 4'd12; b_sign1 = 4'd10; b_sign2 = 4'd2; b_sign3 = 4'd11;
@(posedge clk_i);
a_mant0 = 8'd122; a_mant1 = 8'd71; a_mant2 = 8'd223; a_mant3 = 8'd14;
b_mant0 = 8'd251; b_mant1 = 8'd194; b_mant2 = 8'd179; b_mant3 = 8'd108;
a_exp0 = 10'd28; a_exp1 = 10'd248; a_exp2 = 10'd952; a_exp3 = 10'd204;
b_exp0 = 10'd622; b_exp1 = 10'd880; b_exp2 = 10'd680; b_exp3 = 10'd299;
a_sign0 = 4'd13; a_sign1 = 4'd0; a_sign2 = 4'd2; a_sign3 = 4'd10;
b_sign0 = 4'd5; b_sign1 = 4'd6; b_sign2 = 4'd6; b_sign3 = 4'd1;
@(posedge clk_i);
a_mant0 = 8'd115; a_mant1 = 8'd244; a_mant2 = 8'd91; a_mant3 = 8'd5;
b_mant0 = 8'd23; b_mant1 = 8'd40; b_mant2 = 8'd92; b_mant3 = 8'd228;
a_exp0 = 10'd6; a_exp1 = 10'd243; a_exp2 = 10'd514; a_exp3 = 10'd908;
b_exp0 = 10'd520; b_exp1 = 10'd485; b_exp2 = 10'd949; b_exp3 = 10'd388;
a_sign0 = 4'd5; a_sign1 = 4'd4; a_sign2 = 4'd3; a_sign3 = 4'd0;
b_sign0 = 4'd5; b_sign1 = 4'd13; b_sign2 = 4'd7; b_sign3 = 4'd15;
@(posedge clk_i);
a_mant0 = 8'd84; a_mant1 = 8'd10; a_mant2 = 8'd18; a_mant3 = 8'd226;
b_mant0 = 8'd251; b_mant1 = 8'd211; b_mant2 = 8'd67; b_mant3 = 8'd62;
a_exp0 = 10'd221; a_exp1 = 10'd946; a_exp2 = 10'd145; a_exp3 = 10'd177;
b_exp0 = 10'd316; b_exp1 = 10'd427; b_exp2 = 10'd60; b_exp3 = 10'd429;
a_sign0 = 4'd5; a_sign1 = 4'd16; a_sign2 = 4'd9; a_sign3 = 4'd15;
b_sign0 = 4'd11; b_sign1 = 4'd5; b_sign2 = 4'd6; b_sign3 = 4'd0;
@(posedge clk_i);
a_mant0 = 8'd114; a_mant1 = 8'd209; a_mant2 = 8'd179; a_mant3 = 8'd79;
b_mant0 = 8'd25; b_mant1 = 8'd127; b_mant2 = 8'd222; b_mant3 = 8'd248;
a_exp0 = 10'd1004; a_exp1 = 10'd347; a_exp2 = 10'd516; a_exp3 = 10'd680;
b_exp0 = 10'd684; b_exp1 = 10'd286; b_exp2 = 10'd250; b_exp3 = 10'd560;
a_sign0 = 4'd9; a_sign1 = 4'd7; a_sign2 = 4'd6; a_sign3 = 4'd13;
b_sign0 = 4'd6; b_sign1 = 4'd6; b_sign2 = 4'd9; b_sign3 = 4'd11;
@(posedge clk_i);
a_mant0 = 8'd95; a_mant1 = 8'd181; a_mant2 = 8'd241; a_mant3 = 8'd116;
b_mant0 = 8'd32; b_mant1 = 8'd177; b_mant2 = 8'd78; b_mant3 = 8'd187;
a_exp0 = 10'd966; a_exp1 = 10'd115; a_exp2 = 10'd541; a_exp3 = 10'd499;
b_exp0 = 10'd320; b_exp1 = 10'd696; b_exp2 = 10'd516; b_exp3 = 10'd992;
a_sign0 = 4'd2; a_sign1 = 4'd5; a_sign2 = 4'd14; a_sign3 = 4'd12;
b_sign0 = 4'd0; b_sign1 = 4'd10; b_sign2 = 4'd2; b_sign3 = 4'd12;
@(posedge clk_i);
a_mant0 = 8'd82; a_mant1 = 8'd181; a_mant2 = 8'd58; a_mant3 = 8'd13;
b_mant0 = 8'd159; b_mant1 = 8'd234; b_mant2 = 8'd21; b_mant3 = 8'd193;
a_exp0 = 10'd790; a_exp1 = 10'd498; a_exp2 = 10'd613; a_exp3 = 10'd0;
b_exp0 = 10'd440; b_exp1 = 10'd504; b_exp2 = 10'd310; b_exp3 = 10'd750;
a_sign0 = 4'd4; a_sign1 = 4'd10; a_sign2 = 4'd11; a_sign3 = 4'd6;
b_sign0 = 4'd16; b_sign1 = 4'd4; b_sign2 = 4'd14; b_sign3 = 4'd7;
@(posedge clk_i);
a_mant0 = 8'd134; a_mant1 = 8'd12; a_mant2 = 8'd208; a_mant3 = 8'd7;
b_mant0 = 8'd13; b_mant1 = 8'd165; b_mant2 = 8'd39; b_mant3 = 8'd23;
a_exp0 = 10'd86; a_exp1 = 10'd58; a_exp2 = 10'd996; a_exp3 = 10'd223;
b_exp0 = 10'd836; b_exp1 = 10'd107; b_exp2 = 10'd819; b_exp3 = 10'd402;
a_sign0 = 4'd15; a_sign1 = 4'd10; a_sign2 = 4'd7; a_sign3 = 4'd14;
b_sign0 = 4'd9; b_sign1 = 4'd6; b_sign2 = 4'd14; b_sign3 = 4'd6;
@(posedge clk_i);
shared_exps0 = 8'd154;
shared_exps1 = 8'd109;
a_mant0 = 8'd164; a_mant1 = 8'd111; a_mant2 = 8'd211; a_mant3 = 8'd181;
b_mant0 = 8'd57; b_mant1 = 8'd208; b_mant2 = 8'd48; b_mant3 = 8'd6;
a_exp0 = 10'd613; a_exp1 = 10'd500; a_exp2 = 10'd304; a_exp3 = 10'd410;
b_exp0 = 10'd195; b_exp1 = 10'd1000; b_exp2 = 10'd349; b_exp3 = 10'd248;
a_sign0 = 4'd4; a_sign1 = 4'd15; a_sign2 = 4'd12; a_sign3 = 4'd16;
b_sign0 = 4'd16; b_sign1 = 4'd5; b_sign2 = 4'd0; b_sign3 = 4'd3;
@(posedge clk_i);
a_mant0 = 8'd76; a_mant1 = 8'd187; a_mant2 = 8'd123; a_mant3 = 8'd165;
b_mant0 = 8'd219; b_mant1 = 8'd166; b_mant2 = 8'd248; b_mant3 = 8'd130;
a_exp0 = 10'd373; a_exp1 = 10'd991; a_exp2 = 10'd203; a_exp3 = 10'd751;
b_exp0 = 10'd316; b_exp1 = 10'd775; b_exp2 = 10'd284; b_exp3 = 10'd106;
a_sign0 = 4'd3; a_sign1 = 4'd12; a_sign2 = 4'd12; a_sign3 = 4'd6;
b_sign0 = 4'd6; b_sign1 = 4'd9; b_sign2 = 4'd3; b_sign3 = 4'd9;
@(posedge clk_i);
a_mant0 = 8'd150; a_mant1 = 8'd134; a_mant2 = 8'd168; a_mant3 = 8'd141;
b_mant0 = 8'd222; b_mant1 = 8'd110; b_mant2 = 8'd72; b_mant3 = 8'd190;
a_exp0 = 10'd922; a_exp1 = 10'd791; a_exp2 = 10'd480; a_exp3 = 10'd337;
b_exp0 = 10'd984; b_exp1 = 10'd718; b_exp2 = 10'd403; b_exp3 = 10'd19;
a_sign0 = 4'd15; a_sign1 = 4'd15; a_sign2 = 4'd15; a_sign3 = 4'd11;
b_sign0 = 4'd3; b_sign1 = 4'd6; b_sign2 = 4'd0; b_sign3 = 4'd5;
@(posedge clk_i);
a_mant0 = 8'd149; a_mant1 = 8'd207; a_mant2 = 8'd28; a_mant3 = 8'd128;
b_mant0 = 8'd24; b_mant1 = 8'd107; b_mant2 = 8'd62; b_mant3 = 8'd191;
a_exp0 = 10'd7; a_exp1 = 10'd48; a_exp2 = 10'd335; a_exp3 = 10'd943;
b_exp0 = 10'd123; b_exp1 = 10'd74; b_exp2 = 10'd916; b_exp3 = 10'd509;
a_sign0 = 4'd15; a_sign1 = 4'd1; a_sign2 = 4'd4; a_sign3 = 4'd7;
b_sign0 = 4'd9; b_sign1 = 4'd10; b_sign2 = 4'd0; b_sign3 = 4'd16;
@(posedge clk_i);
a_mant0 = 8'd119; a_mant1 = 8'd166; a_mant2 = 8'd185; a_mant3 = 8'd64;
b_mant0 = 8'd104; b_mant1 = 8'd94; b_mant2 = 8'd82; b_mant3 = 8'd219;
a_exp0 = 10'd317; a_exp1 = 10'd363; a_exp2 = 10'd329; a_exp3 = 10'd944;
b_exp0 = 10'd863; b_exp1 = 10'd619; b_exp2 = 10'd46; b_exp3 = 10'd58;
a_sign0 = 4'd16; a_sign1 = 4'd3; a_sign2 = 4'd7; a_sign3 = 4'd1;
b_sign0 = 4'd7; b_sign1 = 4'd0; b_sign2 = 4'd7; b_sign3 = 4'd2;
@(posedge clk_i);
a_mant0 = 8'd8; a_mant1 = 8'd36; a_mant2 = 8'd215; a_mant3 = 8'd71;
b_mant0 = 8'd16; b_mant1 = 8'd121; b_mant2 = 8'd80; b_mant3 = 8'd241;
a_exp0 = 10'd740; a_exp1 = 10'd959; a_exp2 = 10'd389; a_exp3 = 10'd433;
b_exp0 = 10'd581; b_exp1 = 10'd29; b_exp2 = 10'd446; b_exp3 = 10'd308;
a_sign0 = 4'd15; a_sign1 = 4'd0; a_sign2 = 4'd6; a_sign3 = 4'd15;
b_sign0 = 4'd5; b_sign1 = 4'd14; b_sign2 = 4'd13; b_sign3 = 4'd0;
@(posedge clk_i);
a_mant0 = 8'd39; a_mant1 = 8'd31; a_mant2 = 8'd171; a_mant3 = 8'd232;
b_mant0 = 8'd45; b_mant1 = 8'd90; b_mant2 = 8'd133; b_mant3 = 8'd142;
a_exp0 = 10'd791; a_exp1 = 10'd527; a_exp2 = 10'd443; a_exp3 = 10'd702;
b_exp0 = 10'd998; b_exp1 = 10'd899; b_exp2 = 10'd1015; b_exp3 = 10'd560;
a_sign0 = 4'd11; a_sign1 = 4'd8; a_sign2 = 4'd12; a_sign3 = 4'd1;
b_sign0 = 4'd10; b_sign1 = 4'd11; b_sign2 = 4'd3; b_sign3 = 4'd1;
@(posedge clk_i);
a_mant0 = 8'd117; a_mant1 = 8'd168; a_mant2 = 8'd122; a_mant3 = 8'd74;
b_mant0 = 8'd134; b_mant1 = 8'd197; b_mant2 = 8'd145; b_mant3 = 8'd114;
a_exp0 = 10'd498; a_exp1 = 10'd772; a_exp2 = 10'd865; a_exp3 = 10'd238;
b_exp0 = 10'd579; b_exp1 = 10'd147; b_exp2 = 10'd471; b_exp3 = 10'd827;
a_sign0 = 4'd10; a_sign1 = 4'd12; a_sign2 = 4'd12; a_sign3 = 4'd1;
b_sign0 = 4'd14; b_sign1 = 4'd12; b_sign2 = 4'd0; b_sign3 = 4'd14;
@(posedge clk_i);
shared_exps0 = 8'd159;
shared_exps1 = 8'd106;
a_mant0 = 8'd42; a_mant1 = 8'd243; a_mant2 = 8'd178; a_mant3 = 8'd27;
b_mant0 = 8'd252; b_mant1 = 8'd212; b_mant2 = 8'd185; b_mant3 = 8'd123;
a_exp0 = 10'd896; a_exp1 = 10'd330; a_exp2 = 10'd886; a_exp3 = 10'd817;
b_exp0 = 10'd3; b_exp1 = 10'd879; b_exp2 = 10'd67; b_exp3 = 10'd159;
a_sign0 = 4'd5; a_sign1 = 4'd12; a_sign2 = 4'd5; a_sign3 = 4'd14;
b_sign0 = 4'd10; b_sign1 = 4'd12; b_sign2 = 4'd8; b_sign3 = 4'd6;
@(posedge clk_i);
a_mant0 = 8'd5; a_mant1 = 8'd213; a_mant2 = 8'd38; a_mant3 = 8'd117;
b_mant0 = 8'd62; b_mant1 = 8'd192; b_mant2 = 8'd253; b_mant3 = 8'd190;
a_exp0 = 10'd758; a_exp1 = 10'd1018; a_exp2 = 10'd834; a_exp3 = 10'd661;
b_exp0 = 10'd235; b_exp1 = 10'd700; b_exp2 = 10'd44; b_exp3 = 10'd863;
a_sign0 = 4'd10; a_sign1 = 4'd1; a_sign2 = 4'd11; a_sign3 = 4'd12;
b_sign0 = 4'd2; b_sign1 = 4'd0; b_sign2 = 4'd4; b_sign3 = 4'd13;
@(posedge clk_i);
a_mant0 = 8'd107; a_mant1 = 8'd2; a_mant2 = 8'd141; a_mant3 = 8'd48;
b_mant0 = 8'd180; b_mant1 = 8'd192; b_mant2 = 8'd63; b_mant3 = 8'd197;
a_exp0 = 10'd603; a_exp1 = 10'd543; a_exp2 = 10'd946; a_exp3 = 10'd1009;
b_exp0 = 10'd920; b_exp1 = 10'd124; b_exp2 = 10'd195; b_exp3 = 10'd113;
a_sign0 = 4'd0; a_sign1 = 4'd15; a_sign2 = 4'd9; a_sign3 = 4'd11;
b_sign0 = 4'd12; b_sign1 = 4'd16; b_sign2 = 4'd0; b_sign3 = 4'd8;
@(posedge clk_i);
a_mant0 = 8'd245; a_mant1 = 8'd160; a_mant2 = 8'd115; a_mant3 = 8'd149;
b_mant0 = 8'd134; b_mant1 = 8'd169; b_mant2 = 8'd87; b_mant3 = 8'd125;
a_exp0 = 10'd418; a_exp1 = 10'd964; a_exp2 = 10'd1008; a_exp3 = 10'd512;
b_exp0 = 10'd15; b_exp1 = 10'd105; b_exp2 = 10'd447; b_exp3 = 10'd549;
a_sign0 = 4'd15; a_sign1 = 4'd0; a_sign2 = 4'd1; a_sign3 = 4'd9;
b_sign0 = 4'd3; b_sign1 = 4'd10; b_sign2 = 4'd1; b_sign3 = 4'd10;
@(posedge clk_i);
a_mant0 = 8'd199; a_mant1 = 8'd45; a_mant2 = 8'd62; a_mant3 = 8'd62;
b_mant0 = 8'd90; b_mant1 = 8'd206; b_mant2 = 8'd107; b_mant3 = 8'd237;
a_exp0 = 10'd372; a_exp1 = 10'd694; a_exp2 = 10'd309; a_exp3 = 10'd943;
b_exp0 = 10'd703; b_exp1 = 10'd542; b_exp2 = 10'd699; b_exp3 = 10'd804;
a_sign0 = 4'd15; a_sign1 = 4'd15; a_sign2 = 4'd0; a_sign3 = 4'd2;
b_sign0 = 4'd4; b_sign1 = 4'd0; b_sign2 = 4'd10; b_sign3 = 4'd4;
@(posedge clk_i);
a_mant0 = 8'd151; a_mant1 = 8'd93; a_mant2 = 8'd159; a_mant3 = 8'd213;
b_mant0 = 8'd58; b_mant1 = 8'd228; b_mant2 = 8'd90; b_mant3 = 8'd150;
a_exp0 = 10'd861; a_exp1 = 10'd884; a_exp2 = 10'd91; a_exp3 = 10'd721;
b_exp0 = 10'd148; b_exp1 = 10'd50; b_exp2 = 10'd505; b_exp3 = 10'd257;
a_sign0 = 4'd3; a_sign1 = 4'd3; a_sign2 = 4'd11; a_sign3 = 4'd13;
b_sign0 = 4'd9; b_sign1 = 4'd10; b_sign2 = 4'd8; b_sign3 = 4'd0;
@(posedge clk_i);
a_mant0 = 8'd62; a_mant1 = 8'd209; a_mant2 = 8'd176; a_mant3 = 8'd209;
b_mant0 = 8'd106; b_mant1 = 8'd74; b_mant2 = 8'd214; b_mant3 = 8'd67;
a_exp0 = 10'd200; a_exp1 = 10'd862; a_exp2 = 10'd786; a_exp3 = 10'd881;
b_exp0 = 10'd822; b_exp1 = 10'd859; b_exp2 = 10'd56; b_exp3 = 10'd349;
a_sign0 = 4'd7; a_sign1 = 4'd15; a_sign2 = 4'd5; a_sign3 = 4'd13;
b_sign0 = 4'd11; b_sign1 = 4'd8; b_sign2 = 4'd4; b_sign3 = 4'd8;
@(posedge clk_i);
a_mant0 = 8'd146; a_mant1 = 8'd241; a_mant2 = 8'd13; a_mant3 = 8'd208;
b_mant0 = 8'd88; b_mant1 = 8'd210; b_mant2 = 8'd253; b_mant3 = 8'd126;
a_exp0 = 10'd869; a_exp1 = 10'd462; a_exp2 = 10'd56; a_exp3 = 10'd708;
b_exp0 = 10'd146; b_exp1 = 10'd949; b_exp2 = 10'd140; b_exp3 = 10'd335;
a_sign0 = 4'd16; a_sign1 = 4'd14; a_sign2 = 4'd10; a_sign3 = 4'd15;
b_sign0 = 4'd13; b_sign1 = 4'd11; b_sign2 = 4'd5; b_sign3 = 4'd14;
@(posedge clk_i);
shared_exps0 = 8'd131;
shared_exps1 = 8'd122;
rstn = 0;
@(posedge clk_i);
rstn = 1;
a_mant0 = 8'd251; a_mant1 = 8'd117; a_mant2 = 8'd130; a_mant3 = 8'd194;
b_mant0 = 8'd22; b_mant1 = 8'd95; b_mant2 = 8'd132; b_mant3 = 8'd203;
a_exp0 = 10'd776; a_exp1 = 10'd874; a_exp2 = 10'd432; a_exp3 = 10'd496;
b_exp0 = 10'd180; b_exp1 = 10'd363; b_exp2 = 10'd773; b_exp3 = 10'd772;
a_sign0 = 4'd2; a_sign1 = 4'd10; a_sign2 = 4'd8; a_sign3 = 4'd1;
b_sign0 = 4'd15; b_sign1 = 4'd11; b_sign2 = 4'd15; b_sign3 = 4'd1;
@(posedge clk_i);
a_mant0 = 8'd36; a_mant1 = 8'd106; a_mant2 = 8'd235; a_mant3 = 8'd146;
b_mant0 = 8'd103; b_mant1 = 8'd181; b_mant2 = 8'd37; b_mant3 = 8'd31;
a_exp0 = 10'd754; a_exp1 = 10'd486; a_exp2 = 10'd657; a_exp3 = 10'd206;
b_exp0 = 10'd618; b_exp1 = 10'd0; b_exp2 = 10'd895; b_exp3 = 10'd649;
a_sign0 = 4'd2; a_sign1 = 4'd6; a_sign2 = 4'd14; a_sign3 = 4'd4;
b_sign0 = 4'd11; b_sign1 = 4'd11; b_sign2 = 4'd10; b_sign3 = 4'd9;
@(posedge clk_i);
a_mant0 = 8'd157; a_mant1 = 8'd193; a_mant2 = 8'd44; a_mant3 = 8'd128;
b_mant0 = 8'd143; b_mant1 = 8'd219; b_mant2 = 8'd248; b_mant3 = 8'd138;
a_exp0 = 10'd680; a_exp1 = 10'd521; a_exp2 = 10'd28; a_exp3 = 10'd150;
b_exp0 = 10'd194; b_exp1 = 10'd247; b_exp2 = 10'd381; b_exp3 = 10'd29;
a_sign0 = 4'd16; a_sign1 = 4'd10; a_sign2 = 4'd7; a_sign3 = 4'd6;
b_sign0 = 4'd6; b_sign1 = 4'd11; b_sign2 = 4'd13; b_sign3 = 4'd0;
@(posedge clk_i);
a_mant0 = 8'd31; a_mant1 = 8'd193; a_mant2 = 8'd127; a_mant3 = 8'd132;
b_mant0 = 8'd38; b_mant1 = 8'd92; b_mant2 = 8'd9; b_mant3 = 8'd160;
a_exp0 = 10'd125; a_exp1 = 10'd159; a_exp2 = 10'd1001; a_exp3 = 10'd895;
b_exp0 = 10'd481; b_exp1 = 10'd47; b_exp2 = 10'd902; b_exp3 = 10'd401;
a_sign0 = 4'd6; a_sign1 = 4'd0; a_sign2 = 4'd16; a_sign3 = 4'd0;
b_sign0 = 4'd0; b_sign1 = 4'd12; b_sign2 = 4'd6; b_sign3 = 4'd1;
@(posedge clk_i);
a_mant0 = 8'd125; a_mant1 = 8'd240; a_mant2 = 8'd200; a_mant3 = 8'd112;
b_mant0 = 8'd213; b_mant1 = 8'd40; b_mant2 = 8'd128; b_mant3 = 8'd89;
a_exp0 = 10'd907; a_exp1 = 10'd1010; a_exp2 = 10'd541; a_exp3 = 10'd655;
b_exp0 = 10'd49; b_exp1 = 10'd393; b_exp2 = 10'd1001; b_exp3 = 10'd208;
a_sign0 = 4'd10; a_sign1 = 4'd16; a_sign2 = 4'd12; a_sign3 = 4'd14;
b_sign0 = 4'd1; b_sign1 = 4'd7; b_sign2 = 4'd5; b_sign3 = 4'd10;
@(posedge clk_i);
a_mant0 = 8'd122; a_mant1 = 8'd132; a_mant2 = 8'd60; a_mant3 = 8'd190;
b_mant0 = 8'd223; b_mant1 = 8'd148; b_mant2 = 8'd92; b_mant3 = 8'd131;
a_exp0 = 10'd1; a_exp1 = 10'd986; a_exp2 = 10'd478; a_exp3 = 10'd809;
b_exp0 = 10'd667; b_exp1 = 10'd351; b_exp2 = 10'd317; b_exp3 = 10'd618;
a_sign0 = 4'd6; a_sign1 = 4'd4; a_sign2 = 4'd14; a_sign3 = 4'd14;
b_sign0 = 4'd12; b_sign1 = 4'd6; b_sign2 = 4'd4; b_sign3 = 4'd15;
@(posedge clk_i);
a_mant0 = 8'd130; a_mant1 = 8'd197; a_mant2 = 8'd75; a_mant3 = 8'd46;
b_mant0 = 8'd141; b_mant1 = 8'd79; b_mant2 = 8'd189; b_mant3 = 8'd85;
a_exp0 = 10'd256; a_exp1 = 10'd32; a_exp2 = 10'd575; a_exp3 = 10'd929;
b_exp0 = 10'd766; b_exp1 = 10'd891; b_exp2 = 10'd785; b_exp3 = 10'd71;
a_sign0 = 4'd0; a_sign1 = 4'd2; a_sign2 = 4'd6; a_sign3 = 4'd10;
b_sign0 = 4'd14; b_sign1 = 4'd12; b_sign2 = 4'd9; b_sign3 = 4'd15;
@(posedge clk_i);
shared_exps0 = 8'd124;
shared_exps1 = 8'd147;
a_mant0 = 8'd200; a_mant1 = 8'd20; a_mant2 = 8'd83; a_mant3 = 8'd99;
b_mant0 = 8'd154; b_mant1 = 8'd189; b_mant2 = 8'd47; b_mant3 = 8'd4;
a_exp0 = 10'd848; a_exp1 = 10'd881; a_exp2 = 10'd645; a_exp3 = 10'd466;
b_exp0 = 10'd537; b_exp1 = 10'd145; b_exp2 = 10'd997; b_exp3 = 10'd843;
a_sign0 = 4'd7; a_sign1 = 4'd3; a_sign2 = 4'd16; a_sign3 = 4'd2;
b_sign0 = 4'd8; b_sign1 = 4'd7; b_sign2 = 4'd2; b_sign3 = 4'd5;
@(posedge clk_i);
a_mant0 = 8'd189; a_mant1 = 8'd34; a_mant2 = 8'd235; a_mant3 = 8'd153;
b_mant0 = 8'd80; b_mant1 = 8'd101; b_mant2 = 8'd185; b_mant3 = 8'd13;
a_exp0 = 10'd984; a_exp1 = 10'd943; a_exp2 = 10'd106; a_exp3 = 10'd196;
b_exp0 = 10'd464; b_exp1 = 10'd954; b_exp2 = 10'd984; b_exp3 = 10'd598;
a_sign0 = 4'd2; a_sign1 = 4'd10; a_sign2 = 4'd8; a_sign3 = 4'd3;
b_sign0 = 4'd1; b_sign1 = 4'd13; b_sign2 = 4'd1; b_sign3 = 4'd7;
@(posedge clk_i);
a_mant0 = 8'd126; a_mant1 = 8'd163; a_mant2 = 8'd80; a_mant3 = 8'd228;
b_mant0 = 8'd52; b_mant1 = 8'd38; b_mant2 = 8'd10; b_mant3 = 8'd169;
a_exp0 = 10'd691; a_exp1 = 10'd360; a_exp2 = 10'd987; a_exp3 = 10'd138;
b_exp0 = 10'd155; b_exp1 = 10'd235; b_exp2 = 10'd790; b_exp3 = 10'd48;
a_sign0 = 4'd16; a_sign1 = 4'd5; a_sign2 = 4'd11; a_sign3 = 4'd8;
b_sign0 = 4'd1; b_sign1 = 4'd13; b_sign2 = 4'd8; b_sign3 = 4'd13;
@(posedge clk_i);
a_mant0 = 8'd211; a_mant1 = 8'd44; a_mant2 = 8'd210; a_mant3 = 8'd202;
b_mant0 = 8'd107; b_mant1 = 8'd146; b_mant2 = 8'd138; b_mant3 = 8'd178;
a_exp0 = 10'd785; a_exp1 = 10'd278; a_exp2 = 10'd958; a_exp3 = 10'd239;
b_exp0 = 10'd336; b_exp1 = 10'd260; b_exp2 = 10'd924; b_exp3 = 10'd944;
a_sign0 = 4'd14; a_sign1 = 4'd4; a_sign2 = 4'd16; a_sign3 = 4'd0;
b_sign0 = 4'd10; b_sign1 = 4'd12; b_sign2 = 4'd6; b_sign3 = 4'd11;
@(posedge clk_i);
a_mant0 = 8'd87; a_mant1 = 8'd103; a_mant2 = 8'd90; a_mant3 = 8'd66;
b_mant0 = 8'd105; b_mant1 = 8'd40; b_mant2 = 8'd155; b_mant3 = 8'd68;
a_exp0 = 10'd828; a_exp1 = 10'd854; a_exp2 = 10'd722; a_exp3 = 10'd634;
b_exp0 = 10'd27; b_exp1 = 10'd621; b_exp2 = 10'd575; b_exp3 = 10'd144;
a_sign0 = 4'd2; a_sign1 = 4'd5; a_sign2 = 4'd15; a_sign3 = 4'd6;
b_sign0 = 4'd10; b_sign1 = 4'd15; b_sign2 = 4'd12; b_sign3 = 4'd2;
@(posedge clk_i);
a_mant0 = 8'd223; a_mant1 = 8'd205; a_mant2 = 8'd246; a_mant3 = 8'd64;
b_mant0 = 8'd146; b_mant1 = 8'd220; b_mant2 = 8'd169; b_mant3 = 8'd26;
a_exp0 = 10'd868; a_exp1 = 10'd912; a_exp2 = 10'd989; a_exp3 = 10'd547;
b_exp0 = 10'd867; b_exp1 = 10'd1017; b_exp2 = 10'd880; b_exp3 = 10'd523;
a_sign0 = 4'd0; a_sign1 = 4'd10; a_sign2 = 4'd9; a_sign3 = 4'd9;
b_sign0 = 4'd14; b_sign1 = 4'd6; b_sign2 = 4'd10; b_sign3 = 4'd12;
@(posedge clk_i);
a_mant0 = 8'd213; a_mant1 = 8'd167; a_mant2 = 8'd109; a_mant3 = 8'd52;
b_mant0 = 8'd193; b_mant1 = 8'd253; b_mant2 = 8'd136; b_mant3 = 8'd207;
a_exp0 = 10'd289; a_exp1 = 10'd977; a_exp2 = 10'd179; a_exp3 = 10'd613;
b_exp0 = 10'd928; b_exp1 = 10'd968; b_exp2 = 10'd851; b_exp3 = 10'd738;
a_sign0 = 4'd9; a_sign1 = 4'd11; a_sign2 = 4'd6; a_sign3 = 4'd16;
b_sign0 = 4'd3; b_sign1 = 4'd15; b_sign2 = 4'd7; b_sign3 = 4'd3;
@(posedge clk_i);
a_mant0 = 8'd30; a_mant1 = 8'd37; a_mant2 = 8'd167; a_mant3 = 8'd165;
b_mant0 = 8'd163; b_mant1 = 8'd137; b_mant2 = 8'd14; b_mant3 = 8'd246;
a_exp0 = 10'd431; a_exp1 = 10'd384; a_exp2 = 10'd545; a_exp3 = 10'd15;
b_exp0 = 10'd84; b_exp1 = 10'd244; b_exp2 = 10'd507; b_exp3 = 10'd785;
a_sign0 = 4'd5; a_sign1 = 4'd14; a_sign2 = 4'd8; a_sign3 = 4'd6;
b_sign0 = 4'd12; b_sign1 = 4'd10; b_sign2 = 4'd7; b_sign3 = 4'd0;
@(posedge clk_i);
shared_exps0 = 8'd148;
shared_exps1 = 8'd123;
a_mant0 = 8'd215; a_mant1 = 8'd201; a_mant2 = 8'd39; a_mant3 = 8'd26;
b_mant0 = 8'd15; b_mant1 = 8'd97; b_mant2 = 8'd170; b_mant3 = 8'd187;
a_exp0 = 10'd783; a_exp1 = 10'd994; a_exp2 = 10'd280; a_exp3 = 10'd31;
b_exp0 = 10'd380; b_exp1 = 10'd330; b_exp2 = 10'd326; b_exp3 = 10'd380;
a_sign0 = 4'd6; a_sign1 = 4'd11; a_sign2 = 4'd7; a_sign3 = 4'd13;
b_sign0 = 4'd7; b_sign1 = 4'd8; b_sign2 = 4'd13; b_sign3 = 4'd3;
@(posedge clk_i);
a_mant0 = 8'd101; a_mant1 = 8'd184; a_mant2 = 8'd121; a_mant3 = 8'd206;
b_mant0 = 8'd11; b_mant1 = 8'd31; b_mant2 = 8'd117; b_mant3 = 8'd100;
a_exp0 = 10'd405; a_exp1 = 10'd229; a_exp2 = 10'd1013; a_exp3 = 10'd944;
b_exp0 = 10'd44; b_exp1 = 10'd211; b_exp2 = 10'd163; b_exp3 = 10'd695;
a_sign0 = 4'd5; a_sign1 = 4'd9; a_sign2 = 4'd0; a_sign3 = 4'd9;
b_sign0 = 4'd7; b_sign1 = 4'd5; b_sign2 = 4'd2; b_sign3 = 4'd16;
@(posedge clk_i);
a_mant0 = 8'd81; a_mant1 = 8'd143; a_mant2 = 8'd132; a_mant3 = 8'd53;
b_mant0 = 8'd243; b_mant1 = 8'd237; b_mant2 = 8'd86; b_mant3 = 8'd104;
a_exp0 = 10'd615; a_exp1 = 10'd761; a_exp2 = 10'd787; a_exp3 = 10'd857;
b_exp0 = 10'd557; b_exp1 = 10'd978; b_exp2 = 10'd909; b_exp3 = 10'd551;
a_sign0 = 4'd0; a_sign1 = 4'd1; a_sign2 = 4'd12; a_sign3 = 4'd13;
b_sign0 = 4'd6; b_sign1 = 4'd9; b_sign2 = 4'd16; b_sign3 = 4'd11;
@(posedge clk_i);
a_mant0 = 8'd243; a_mant1 = 8'd116; a_mant2 = 8'd151; a_mant3 = 8'd166;
b_mant0 = 8'd43; b_mant1 = 8'd235; b_mant2 = 8'd27; b_mant3 = 8'd218;
a_exp0 = 10'd204; a_exp1 = 10'd750; a_exp2 = 10'd435; a_exp3 = 10'd234;
b_exp0 = 10'd780; b_exp1 = 10'd144; b_exp2 = 10'd1017; b_exp3 = 10'd318;
a_sign0 = 4'd11; a_sign1 = 4'd1; a_sign2 = 4'd2; a_sign3 = 4'd2;
b_sign0 = 4'd8; b_sign1 = 4'd5; b_sign2 = 4'd2; b_sign3 = 4'd6;
@(posedge clk_i);
a_mant0 = 8'd116; a_mant1 = 8'd67; a_mant2 = 8'd220; a_mant3 = 8'd184;
b_mant0 = 8'd227; b_mant1 = 8'd170; b_mant2 = 8'd31; b_mant3 = 8'd244;
a_exp0 = 10'd438; a_exp1 = 10'd937; a_exp2 = 10'd491; a_exp3 = 10'd56;
b_exp0 = 10'd398; b_exp1 = 10'd497; b_exp2 = 10'd28; b_exp3 = 10'd40;
a_sign0 = 4'd14; a_sign1 = 4'd15; a_sign2 = 4'd6; a_sign3 = 4'd1;
b_sign0 = 4'd9; b_sign1 = 4'd4; b_sign2 = 4'd5; b_sign3 = 4'd16;
@(posedge clk_i);
a_mant0 = 8'd13; a_mant1 = 8'd130; a_mant2 = 8'd242; a_mant3 = 8'd140;
b_mant0 = 8'd73; b_mant1 = 8'd90; b_mant2 = 8'd180; b_mant3 = 8'd111;
a_exp0 = 10'd383; a_exp1 = 10'd226; a_exp2 = 10'd12; a_exp3 = 10'd229;
b_exp0 = 10'd585; b_exp1 = 10'd315; b_exp2 = 10'd64; b_exp3 = 10'd127;
a_sign0 = 4'd1; a_sign1 = 4'd10; a_sign2 = 4'd11; a_sign3 = 4'd16;
b_sign0 = 4'd15; b_sign1 = 4'd11; b_sign2 = 4'd14; b_sign3 = 4'd8;
@(posedge clk_i);
a_mant0 = 8'd198; a_mant1 = 8'd149; a_mant2 = 8'd198; a_mant3 = 8'd40;
b_mant0 = 8'd83; b_mant1 = 8'd154; b_mant2 = 8'd189; b_mant3 = 8'd18;
a_exp0 = 10'd804; a_exp1 = 10'd825; a_exp2 = 10'd998; a_exp3 = 10'd444;
b_exp0 = 10'd474; b_exp1 = 10'd950; b_exp2 = 10'd75; b_exp3 = 10'd27;
a_sign0 = 4'd6; a_sign1 = 4'd15; a_sign2 = 4'd5; a_sign3 = 4'd10;
b_sign0 = 4'd6; b_sign1 = 4'd11; b_sign2 = 4'd7; b_sign3 = 4'd1;
@(posedge clk_i);
a_mant0 = 8'd112; a_mant1 = 8'd161; a_mant2 = 8'd75; a_mant3 = 8'd66;
b_mant0 = 8'd190; b_mant1 = 8'd77; b_mant2 = 8'd237; b_mant3 = 8'd247;
a_exp0 = 10'd772; a_exp1 = 10'd804; a_exp2 = 10'd634; a_exp3 = 10'd310;
b_exp0 = 10'd759; b_exp1 = 10'd752; b_exp2 = 10'd140; b_exp3 = 10'd134;
a_sign0 = 4'd0; a_sign1 = 4'd10; a_sign2 = 4'd12; a_sign3 = 4'd6;
b_sign0 = 4'd13; b_sign1 = 4'd5; b_sign2 = 4'd6; b_sign3 = 4'd2;
@(posedge clk_i);
shared_exps0 = 8'd133;
shared_exps1 = 8'd148;
a_mant0 = 8'd115; a_mant1 = 8'd173; a_mant2 = 8'd246; a_mant3 = 8'd45;
b_mant0 = 8'd167; b_mant1 = 8'd37; b_mant2 = 8'd207; b_mant3 = 8'd0;
a_exp0 = 10'd263; a_exp1 = 10'd1016; a_exp2 = 10'd220; a_exp3 = 10'd378;
b_exp0 = 10'd276; b_exp1 = 10'd826; b_exp2 = 10'd836; b_exp3 = 10'd166;
a_sign0 = 4'd8; a_sign1 = 4'd15; a_sign2 = 4'd13; a_sign3 = 4'd1;
b_sign0 = 4'd3; b_sign1 = 4'd1; b_sign2 = 4'd11; b_sign3 = 4'd0;
@(posedge clk_i);
a_mant0 = 8'd16; a_mant1 = 8'd162; a_mant2 = 8'd30; a_mant3 = 8'd188;
b_mant0 = 8'd66; b_mant1 = 8'd204; b_mant2 = 8'd54; b_mant3 = 8'd110;
a_exp0 = 10'd52; a_exp1 = 10'd248; a_exp2 = 10'd625; a_exp3 = 10'd354;
b_exp0 = 10'd540; b_exp1 = 10'd131; b_exp2 = 10'd359; b_exp3 = 10'd686;
a_sign0 = 4'd4; a_sign1 = 4'd2; a_sign2 = 4'd6; a_sign3 = 4'd10;
b_sign0 = 4'd6; b_sign1 = 4'd2; b_sign2 = 4'd1; b_sign3 = 4'd8;
@(posedge clk_i);
a_mant0 = 8'd229; a_mant1 = 8'd54; a_mant2 = 8'd80; a_mant3 = 8'd25;
b_mant0 = 8'd210; b_mant1 = 8'd252; b_mant2 = 8'd80; b_mant3 = 8'd196;
a_exp0 = 10'd344; a_exp1 = 10'd279; a_exp2 = 10'd849; a_exp3 = 10'd625;
b_exp0 = 10'd622; b_exp1 = 10'd908; b_exp2 = 10'd326; b_exp3 = 10'd427;
a_sign0 = 4'd11; a_sign1 = 4'd16; a_sign2 = 4'd9; a_sign3 = 4'd15;
b_sign0 = 4'd7; b_sign1 = 4'd7; b_sign2 = 4'd4; b_sign3 = 4'd16;
@(posedge clk_i);
a_mant0 = 8'd174; a_mant1 = 8'd8; a_mant2 = 8'd10; a_mant3 = 8'd90;
b_mant0 = 8'd228; b_mant1 = 8'd96; b_mant2 = 8'd158; b_mant3 = 8'd133;
a_exp0 = 10'd95; a_exp1 = 10'd476; a_exp2 = 10'd631; a_exp3 = 10'd477;
b_exp0 = 10'd1019; b_exp1 = 10'd864; b_exp2 = 10'd279; b_exp3 = 10'd247;
a_sign0 = 4'd12; a_sign1 = 4'd14; a_sign2 = 4'd9; a_sign3 = 4'd6;
b_sign0 = 4'd5; b_sign1 = 4'd2; b_sign2 = 4'd5; b_sign3 = 4'd4;
@(posedge clk_i);
a_mant0 = 8'd104; a_mant1 = 8'd173; a_mant2 = 8'd113; a_mant3 = 8'd38;
b_mant0 = 8'd69; b_mant1 = 8'd174; b_mant2 = 8'd39; b_mant3 = 8'd12;
a_exp0 = 10'd467; a_exp1 = 10'd807; a_exp2 = 10'd579; a_exp3 = 10'd300;
b_exp0 = 10'd345; b_exp1 = 10'd455; b_exp2 = 10'd76; b_exp3 = 10'd473;
a_sign0 = 4'd5; a_sign1 = 4'd14; a_sign2 = 4'd11; a_sign3 = 4'd6;
b_sign0 = 4'd8; b_sign1 = 4'd8; b_sign2 = 4'd6; b_sign3 = 4'd13;
@(posedge clk_i);
a_mant0 = 8'd188; a_mant1 = 8'd85; a_mant2 = 8'd100; a_mant3 = 8'd162;
b_mant0 = 8'd84; b_mant1 = 8'd238; b_mant2 = 8'd135; b_mant3 = 8'd122;
a_exp0 = 10'd631; a_exp1 = 10'd492; a_exp2 = 10'd571; a_exp3 = 10'd105;
b_exp0 = 10'd62; b_exp1 = 10'd966; b_exp2 = 10'd160; b_exp3 = 10'd244;
a_sign0 = 4'd4; a_sign1 = 4'd15; a_sign2 = 4'd1; a_sign3 = 4'd7;
b_sign0 = 4'd5; b_sign1 = 4'd14; b_sign2 = 4'd13; b_sign3 = 4'd10;
@(posedge clk_i);
a_mant0 = 8'd84; a_mant1 = 8'd100; a_mant2 = 8'd108; a_mant3 = 8'd152;
b_mant0 = 8'd117; b_mant1 = 8'd86; b_mant2 = 8'd81; b_mant3 = 8'd93;
a_exp0 = 10'd873; a_exp1 = 10'd735; a_exp2 = 10'd162; a_exp3 = 10'd401;
b_exp0 = 10'd656; b_exp1 = 10'd653; b_exp2 = 10'd563; b_exp3 = 10'd572;
a_sign0 = 4'd11; a_sign1 = 4'd2; a_sign2 = 4'd11; a_sign3 = 4'd5;
b_sign0 = 4'd3; b_sign1 = 4'd10; b_sign2 = 4'd2; b_sign3 = 4'd13;
@(posedge clk_i);
a_mant0 = 8'd55; a_mant1 = 8'd85; a_mant2 = 8'd117; a_mant3 = 8'd23;
b_mant0 = 8'd47; b_mant1 = 8'd44; b_mant2 = 8'd8; b_mant3 = 8'd92;
a_exp0 = 10'd840; a_exp1 = 10'd775; a_exp2 = 10'd791; a_exp3 = 10'd270;
b_exp0 = 10'd163; b_exp1 = 10'd364; b_exp2 = 10'd718; b_exp3 = 10'd427;
a_sign0 = 4'd14; a_sign1 = 4'd4; a_sign2 = 4'd0; a_sign3 = 4'd4;
b_sign0 = 4'd16; b_sign1 = 4'd12; b_sign2 = 4'd10; b_sign3 = 4'd12;
@(posedge clk_i);
shared_exps0 = 8'd159;
shared_exps1 = 8'd110;
rstn = 0;
@(posedge clk_i);
rstn = 1;
a_mant0 = 8'd156; a_mant1 = 8'd132; a_mant2 = 8'd196; a_mant3 = 8'd245;
b_mant0 = 8'd120; b_mant1 = 8'd137; b_mant2 = 8'd108; b_mant3 = 8'd250;
a_exp0 = 10'd833; a_exp1 = 10'd783; a_exp2 = 10'd476; a_exp3 = 10'd411;
b_exp0 = 10'd1002; b_exp1 = 10'd550; b_exp2 = 10'd487; b_exp3 = 10'd396;
a_sign0 = 4'd11; a_sign1 = 4'd10; a_sign2 = 4'd13; a_sign3 = 4'd3;
b_sign0 = 4'd1; b_sign1 = 4'd12; b_sign2 = 4'd1; b_sign3 = 4'd4;
@(posedge clk_i);
a_mant0 = 8'd89; a_mant1 = 8'd37; a_mant2 = 8'd89; a_mant3 = 8'd45;
b_mant0 = 8'd146; b_mant1 = 8'd49; b_mant2 = 8'd137; b_mant3 = 8'd141;
a_exp0 = 10'd769; a_exp1 = 10'd861; a_exp2 = 10'd192; a_exp3 = 10'd989;
b_exp0 = 10'd441; b_exp1 = 10'd574; b_exp2 = 10'd407; b_exp3 = 10'd244;
a_sign0 = 4'd7; a_sign1 = 4'd8; a_sign2 = 4'd2; a_sign3 = 4'd2;
b_sign0 = 4'd8; b_sign1 = 4'd16; b_sign2 = 4'd10; b_sign3 = 4'd11;
@(posedge clk_i);
a_mant0 = 8'd153; a_mant1 = 8'd35; a_mant2 = 8'd179; a_mant3 = 8'd231;
b_mant0 = 8'd26; b_mant1 = 8'd245; b_mant2 = 8'd157; b_mant3 = 8'd62;
a_exp0 = 10'd571; a_exp1 = 10'd574; a_exp2 = 10'd272; a_exp3 = 10'd688;
b_exp0 = 10'd1002; b_exp1 = 10'd787; b_exp2 = 10'd818; b_exp3 = 10'd418;
a_sign0 = 4'd2; a_sign1 = 4'd5; a_sign2 = 4'd9; a_sign3 = 4'd4;
b_sign0 = 4'd4; b_sign1 = 4'd0; b_sign2 = 4'd6; b_sign3 = 4'd15;
@(posedge clk_i);
a_mant0 = 8'd246; a_mant1 = 8'd67; a_mant2 = 8'd12; a_mant3 = 8'd93;
b_mant0 = 8'd74; b_mant1 = 8'd63; b_mant2 = 8'd174; b_mant3 = 8'd28;
a_exp0 = 10'd962; a_exp1 = 10'd963; a_exp2 = 10'd32; a_exp3 = 10'd750;
b_exp0 = 10'd129; b_exp1 = 10'd276; b_exp2 = 10'd510; b_exp3 = 10'd636;
a_sign0 = 4'd4; a_sign1 = 4'd6; a_sign2 = 4'd15; a_sign3 = 4'd8;
b_sign0 = 4'd11; b_sign1 = 4'd0; b_sign2 = 4'd15; b_sign3 = 4'd5;
@(posedge clk_i);
a_mant0 = 8'd28; a_mant1 = 8'd184; a_mant2 = 8'd82; a_mant3 = 8'd194;
b_mant0 = 8'd198; b_mant1 = 8'd96; b_mant2 = 8'd56; b_mant3 = 8'd55;
a_exp0 = 10'd575; a_exp1 = 10'd286; a_exp2 = 10'd7; a_exp3 = 10'd679;
b_exp0 = 10'd215; b_exp1 = 10'd115; b_exp2 = 10'd643; b_exp3 = 10'd507;
a_sign0 = 4'd16; a_sign1 = 4'd2; a_sign2 = 4'd12; a_sign3 = 4'd5;
b_sign0 = 4'd3; b_sign1 = 4'd2; b_sign2 = 4'd3; b_sign3 = 4'd4;
@(posedge clk_i);
a_mant0 = 8'd157; a_mant1 = 8'd115; a_mant2 = 8'd145; a_mant3 = 8'd5;
b_mant0 = 8'd78; b_mant1 = 8'd11; b_mant2 = 8'd222; b_mant3 = 8'd97;
a_exp0 = 10'd368; a_exp1 = 10'd812; a_exp2 = 10'd832; a_exp3 = 10'd77;
b_exp0 = 10'd628; b_exp1 = 10'd910; b_exp2 = 10'd568; b_exp3 = 10'd549;
a_sign0 = 4'd12; a_sign1 = 4'd16; a_sign2 = 4'd15; a_sign3 = 4'd5;
b_sign0 = 4'd2; b_sign1 = 4'd8; b_sign2 = 4'd13; b_sign3 = 4'd4;
@(posedge clk_i);
a_mant0 = 8'd251; a_mant1 = 8'd202; a_mant2 = 8'd196; a_mant3 = 8'd165;
b_mant0 = 8'd104; b_mant1 = 8'd93; b_mant2 = 8'd51; b_mant3 = 8'd71;
a_exp0 = 10'd421; a_exp1 = 10'd202; a_exp2 = 10'd549; a_exp3 = 10'd829;
b_exp0 = 10'd768; b_exp1 = 10'd534; b_exp2 = 10'd686; b_exp3 = 10'd894;
a_sign0 = 4'd2; a_sign1 = 4'd14; a_sign2 = 4'd2; a_sign3 = 4'd8;
b_sign0 = 4'd7; b_sign1 = 4'd8; b_sign2 = 4'd5; b_sign3 = 4'd12;
@(posedge clk_i);
shared_exps0 = 8'd127;
shared_exps1 = 8'd161;
a_mant0 = 8'd181; a_mant1 = 8'd175; a_mant2 = 8'd160; a_mant3 = 8'd158;
b_mant0 = 8'd47; b_mant1 = 8'd222; b_mant2 = 8'd1; b_mant3 = 8'd78;
a_exp0 = 10'd599; a_exp1 = 10'd126; a_exp2 = 10'd2; a_exp3 = 10'd556;
b_exp0 = 10'd758; b_exp1 = 10'd537; b_exp2 = 10'd828; b_exp3 = 10'd550;
a_sign0 = 4'd12; a_sign1 = 4'd7; a_sign2 = 4'd3; a_sign3 = 4'd12;
b_sign0 = 4'd3; b_sign1 = 4'd11; b_sign2 = 4'd6; b_sign3 = 4'd14;
@(posedge clk_i);
a_mant0 = 8'd64; a_mant1 = 8'd255; a_mant2 = 8'd55; a_mant3 = 8'd255;
b_mant0 = 8'd40; b_mant1 = 8'd110; b_mant2 = 8'd219; b_mant3 = 8'd211;
a_exp0 = 10'd717; a_exp1 = 10'd748; a_exp2 = 10'd908; a_exp3 = 10'd244;
b_exp0 = 10'd77; b_exp1 = 10'd26; b_exp2 = 10'd863; b_exp3 = 10'd883;
a_sign0 = 4'd8; a_sign1 = 4'd11; a_sign2 = 4'd10; a_sign3 = 4'd16;
b_sign0 = 4'd2; b_sign1 = 4'd5; b_sign2 = 4'd9; b_sign3 = 4'd9;
@(posedge clk_i);
a_mant0 = 8'd98; a_mant1 = 8'd193; a_mant2 = 8'd15; a_mant3 = 8'd38;
b_mant0 = 8'd43; b_mant1 = 8'd26; b_mant2 = 8'd183; b_mant3 = 8'd61;
a_exp0 = 10'd161; a_exp1 = 10'd708; a_exp2 = 10'd978; a_exp3 = 10'd693;
b_exp0 = 10'd817; b_exp1 = 10'd461; b_exp2 = 10'd712; b_exp3 = 10'd464;
a_sign0 = 4'd0; a_sign1 = 4'd13; a_sign2 = 4'd12; a_sign3 = 4'd5;
b_sign0 = 4'd5; b_sign1 = 4'd11; b_sign2 = 4'd8; b_sign3 = 4'd2;
@(posedge clk_i);
a_mant0 = 8'd57; a_mant1 = 8'd244; a_mant2 = 8'd64; a_mant3 = 8'd52;
b_mant0 = 8'd246; b_mant1 = 8'd88; b_mant2 = 8'd19; b_mant3 = 8'd128;
a_exp0 = 10'd662; a_exp1 = 10'd389; a_exp2 = 10'd958; a_exp3 = 10'd34;
b_exp0 = 10'd590; b_exp1 = 10'd963; b_exp2 = 10'd796; b_exp3 = 10'd798;
a_sign0 = 4'd3; a_sign1 = 4'd0; a_sign2 = 4'd14; a_sign3 = 4'd15;
b_sign0 = 4'd6; b_sign1 = 4'd2; b_sign2 = 4'd10; b_sign3 = 4'd12;
@(posedge clk_i);
a_mant0 = 8'd43; a_mant1 = 8'd77; a_mant2 = 8'd199; a_mant3 = 8'd39;
b_mant0 = 8'd199; b_mant1 = 8'd79; b_mant2 = 8'd126; b_mant3 = 8'd75;
a_exp0 = 10'd60; a_exp1 = 10'd176; a_exp2 = 10'd939; a_exp3 = 10'd324;
b_exp0 = 10'd713; b_exp1 = 10'd516; b_exp2 = 10'd924; b_exp3 = 10'd662;
a_sign0 = 4'd8; a_sign1 = 4'd5; a_sign2 = 4'd14; a_sign3 = 4'd9;
b_sign0 = 4'd1; b_sign1 = 4'd13; b_sign2 = 4'd12; b_sign3 = 4'd0;
@(posedge clk_i);
a_mant0 = 8'd61; a_mant1 = 8'd161; a_mant2 = 8'd222; a_mant3 = 8'd202;
b_mant0 = 8'd57; b_mant1 = 8'd46; b_mant2 = 8'd11; b_mant3 = 8'd23;
a_exp0 = 10'd284; a_exp1 = 10'd935; a_exp2 = 10'd669; a_exp3 = 10'd558;
b_exp0 = 10'd394; b_exp1 = 10'd901; b_exp2 = 10'd885; b_exp3 = 10'd294;
a_sign0 = 4'd11; a_sign1 = 4'd14; a_sign2 = 4'd4; a_sign3 = 4'd1;
b_sign0 = 4'd14; b_sign1 = 4'd10; b_sign2 = 4'd6; b_sign3 = 4'd4;
@(posedge clk_i);
a_mant0 = 8'd238; a_mant1 = 8'd15; a_mant2 = 8'd67; a_mant3 = 8'd231;
b_mant0 = 8'd134; b_mant1 = 8'd252; b_mant2 = 8'd138; b_mant3 = 8'd194;
a_exp0 = 10'd961; a_exp1 = 10'd285; a_exp2 = 10'd169; a_exp3 = 10'd585;
b_exp0 = 10'd823; b_exp1 = 10'd95; b_exp2 = 10'd997; b_exp3 = 10'd496;
a_sign0 = 4'd3; a_sign1 = 4'd13; a_sign2 = 4'd16; a_sign3 = 4'd15;
b_sign0 = 4'd7; b_sign1 = 4'd10; b_sign2 = 4'd10; b_sign3 = 4'd1;
@(posedge clk_i);
a_mant0 = 8'd51; a_mant1 = 8'd184; a_mant2 = 8'd61; a_mant3 = 8'd50;
b_mant0 = 8'd49; b_mant1 = 8'd242; b_mant2 = 8'd18; b_mant3 = 8'd130;
a_exp0 = 10'd455; a_exp1 = 10'd253; a_exp2 = 10'd818; a_exp3 = 10'd1019;
b_exp0 = 10'd356; b_exp1 = 10'd137; b_exp2 = 10'd543; b_exp3 = 10'd185;
a_sign0 = 4'd13; a_sign1 = 4'd2; a_sign2 = 4'd14; a_sign3 = 4'd4;
b_sign0 = 4'd10; b_sign1 = 4'd0; b_sign2 = 4'd3; b_sign3 = 4'd3;
@(posedge clk_i);
shared_exps0 = 8'd120;
shared_exps1 = 8'd121;
a_mant0 = 8'd54; a_mant1 = 8'd201; a_mant2 = 8'd70; a_mant3 = 8'd216;
b_mant0 = 8'd134; b_mant1 = 8'd89; b_mant2 = 8'd155; b_mant3 = 8'd15;
a_exp0 = 10'd943; a_exp1 = 10'd743; a_exp2 = 10'd760; a_exp3 = 10'd830;
b_exp0 = 10'd877; b_exp1 = 10'd115; b_exp2 = 10'd130; b_exp3 = 10'd369;
a_sign0 = 4'd7; a_sign1 = 4'd10; a_sign2 = 4'd4; a_sign3 = 4'd6;
b_sign0 = 4'd4; b_sign1 = 4'd8; b_sign2 = 4'd15; b_sign3 = 4'd10;
@(posedge clk_i);
a_mant0 = 8'd130; a_mant1 = 8'd243; a_mant2 = 8'd115; a_mant3 = 8'd120;
b_mant0 = 8'd199; b_mant1 = 8'd149; b_mant2 = 8'd242; b_mant3 = 8'd169;
a_exp0 = 10'd906; a_exp1 = 10'd691; a_exp2 = 10'd14; a_exp3 = 10'd560;
b_exp0 = 10'd82; b_exp1 = 10'd815; b_exp2 = 10'd499; b_exp3 = 10'd666;
a_sign0 = 4'd5; a_sign1 = 4'd11; a_sign2 = 4'd14; a_sign3 = 4'd6;
b_sign0 = 4'd3; b_sign1 = 4'd8; b_sign2 = 4'd8; b_sign3 = 4'd15;
@(posedge clk_i);
a_mant0 = 8'd205; a_mant1 = 8'd42; a_mant2 = 8'd28; a_mant3 = 8'd57;
b_mant0 = 8'd121; b_mant1 = 8'd202; b_mant2 = 8'd189; b_mant3 = 8'd150;
a_exp0 = 10'd834; a_exp1 = 10'd4; a_exp2 = 10'd688; a_exp3 = 10'd256;
b_exp0 = 10'd32; b_exp1 = 10'd683; b_exp2 = 10'd411; b_exp3 = 10'd1000;
a_sign0 = 4'd14; a_sign1 = 4'd4; a_sign2 = 4'd1; a_sign3 = 4'd5;
b_sign0 = 4'd3; b_sign1 = 4'd8; b_sign2 = 4'd8; b_sign3 = 4'd12;
@(posedge clk_i);
a_mant0 = 8'd20; a_mant1 = 8'd254; a_mant2 = 8'd181; a_mant3 = 8'd15;
b_mant0 = 8'd88; b_mant1 = 8'd10; b_mant2 = 8'd222; b_mant3 = 8'd11;
a_exp0 = 10'd51; a_exp1 = 10'd386; a_exp2 = 10'd838; a_exp3 = 10'd5;
b_exp0 = 10'd13; b_exp1 = 10'd424; b_exp2 = 10'd603; b_exp3 = 10'd902;
a_sign0 = 4'd12; a_sign1 = 4'd6; a_sign2 = 4'd3; a_sign3 = 4'd3;
b_sign0 = 4'd2; b_sign1 = 4'd5; b_sign2 = 4'd0; b_sign3 = 4'd7;
@(posedge clk_i);
a_mant0 = 8'd108; a_mant1 = 8'd161; a_mant2 = 8'd104; a_mant3 = 8'd190;
b_mant0 = 8'd229; b_mant1 = 8'd34; b_mant2 = 8'd75; b_mant3 = 8'd234;
a_exp0 = 10'd807; a_exp1 = 10'd399; a_exp2 = 10'd742; a_exp3 = 10'd888;
b_exp0 = 10'd430; b_exp1 = 10'd585; b_exp2 = 10'd426; b_exp3 = 10'd83;
a_sign0 = 4'd1; a_sign1 = 4'd8; a_sign2 = 4'd7; a_sign3 = 4'd5;
b_sign0 = 4'd13; b_sign1 = 4'd12; b_sign2 = 4'd13; b_sign3 = 4'd16;
@(posedge clk_i);
a_mant0 = 8'd128; a_mant1 = 8'd255; a_mant2 = 8'd81; a_mant3 = 8'd43;
b_mant0 = 8'd232; b_mant1 = 8'd96; b_mant2 = 8'd42; b_mant3 = 8'd80;
a_exp0 = 10'd386; a_exp1 = 10'd612; a_exp2 = 10'd948; a_exp3 = 10'd255;
b_exp0 = 10'd79; b_exp1 = 10'd995; b_exp2 = 10'd728; b_exp3 = 10'd912;
a_sign0 = 4'd6; a_sign1 = 4'd4; a_sign2 = 4'd6; a_sign3 = 4'd9;
b_sign0 = 4'd6; b_sign1 = 4'd3; b_sign2 = 4'd15; b_sign3 = 4'd7;
@(posedge clk_i);
a_mant0 = 8'd199; a_mant1 = 8'd253; a_mant2 = 8'd108; a_mant3 = 8'd157;
b_mant0 = 8'd98; b_mant1 = 8'd216; b_mant2 = 8'd72; b_mant3 = 8'd82;
a_exp0 = 10'd382; a_exp1 = 10'd802; a_exp2 = 10'd601; a_exp3 = 10'd252;
b_exp0 = 10'd200; b_exp1 = 10'd106; b_exp2 = 10'd685; b_exp3 = 10'd16;
a_sign0 = 4'd15; a_sign1 = 4'd7; a_sign2 = 4'd15; a_sign3 = 4'd10;
b_sign0 = 4'd4; b_sign1 = 4'd13; b_sign2 = 4'd0; b_sign3 = 4'd6;
@(posedge clk_i);
a_mant0 = 8'd13; a_mant1 = 8'd8; a_mant2 = 8'd76; a_mant3 = 8'd17;
b_mant0 = 8'd141; b_mant1 = 8'd225; b_mant2 = 8'd248; b_mant3 = 8'd130;
a_exp0 = 10'd53; a_exp1 = 10'd215; a_exp2 = 10'd984; a_exp3 = 10'd977;
b_exp0 = 10'd664; b_exp1 = 10'd93; b_exp2 = 10'd83; b_exp3 = 10'd713;
a_sign0 = 4'd15; a_sign1 = 4'd10; a_sign2 = 4'd1; a_sign3 = 4'd13;
b_sign0 = 4'd3; b_sign1 = 4'd3; b_sign2 = 4'd3; b_sign3 = 4'd2;
@(posedge clk_i);
shared_exps0 = 8'd118;
shared_exps1 = 8'd99;
a_mant0 = 8'd117; a_mant1 = 8'd86; a_mant2 = 8'd116; a_mant3 = 8'd19;
b_mant0 = 8'd191; b_mant1 = 8'd166; b_mant2 = 8'd218; b_mant3 = 8'd208;
a_exp0 = 10'd530; a_exp1 = 10'd332; a_exp2 = 10'd824; a_exp3 = 10'd395;
b_exp0 = 10'd518; b_exp1 = 10'd56; b_exp2 = 10'd724; b_exp3 = 10'd96;
a_sign0 = 4'd14; a_sign1 = 4'd16; a_sign2 = 4'd2; a_sign3 = 4'd0;
b_sign0 = 4'd12; b_sign1 = 4'd15; b_sign2 = 4'd12; b_sign3 = 4'd10;
@(posedge clk_i);
a_mant0 = 8'd5; a_mant1 = 8'd36; a_mant2 = 8'd13; a_mant3 = 8'd92;
b_mant0 = 8'd73; b_mant1 = 8'd254; b_mant2 = 8'd192; b_mant3 = 8'd105;
a_exp0 = 10'd217; a_exp1 = 10'd176; a_exp2 = 10'd325; a_exp3 = 10'd988;
b_exp0 = 10'd63; b_exp1 = 10'd911; b_exp2 = 10'd272; b_exp3 = 10'd584;
a_sign0 = 4'd10; a_sign1 = 4'd5; a_sign2 = 4'd15; a_sign3 = 4'd8;
b_sign0 = 4'd4; b_sign1 = 4'd7; b_sign2 = 4'd13; b_sign3 = 4'd6;
@(posedge clk_i);
a_mant0 = 8'd129; a_mant1 = 8'd44; a_mant2 = 8'd72; a_mant3 = 8'd47;
b_mant0 = 8'd98; b_mant1 = 8'd133; b_mant2 = 8'd213; b_mant3 = 8'd26;
a_exp0 = 10'd868; a_exp1 = 10'd722; a_exp2 = 10'd426; a_exp3 = 10'd567;
b_exp0 = 10'd37; b_exp1 = 10'd127; b_exp2 = 10'd534; b_exp3 = 10'd711;
a_sign0 = 4'd4; a_sign1 = 4'd16; a_sign2 = 4'd16; a_sign3 = 4'd3;
b_sign0 = 4'd10; b_sign1 = 4'd10; b_sign2 = 4'd15; b_sign3 = 4'd3;
@(posedge clk_i);
a_mant0 = 8'd91; a_mant1 = 8'd112; a_mant2 = 8'd116; a_mant3 = 8'd44;
b_mant0 = 8'd105; b_mant1 = 8'd163; b_mant2 = 8'd102; b_mant3 = 8'd253;
a_exp0 = 10'd553; a_exp1 = 10'd169; a_exp2 = 10'd409; a_exp3 = 10'd671;
b_exp0 = 10'd284; b_exp1 = 10'd794; b_exp2 = 10'd689; b_exp3 = 10'd483;
a_sign0 = 4'd8; a_sign1 = 4'd5; a_sign2 = 4'd8; a_sign3 = 4'd10;
b_sign0 = 4'd2; b_sign1 = 4'd4; b_sign2 = 4'd7; b_sign3 = 4'd14;
@(posedge clk_i);
a_mant0 = 8'd68; a_mant1 = 8'd255; a_mant2 = 8'd40; a_mant3 = 8'd235;
b_mant0 = 8'd11; b_mant1 = 8'd215; b_mant2 = 8'd38; b_mant3 = 8'd127;
a_exp0 = 10'd301; a_exp1 = 10'd372; a_exp2 = 10'd749; a_exp3 = 10'd526;
b_exp0 = 10'd876; b_exp1 = 10'd212; b_exp2 = 10'd366; b_exp3 = 10'd476;
a_sign0 = 4'd10; a_sign1 = 4'd6; a_sign2 = 4'd3; a_sign3 = 4'd16;
b_sign0 = 4'd0; b_sign1 = 4'd2; b_sign2 = 4'd16; b_sign3 = 4'd6;
@(posedge clk_i);
a_mant0 = 8'd111; a_mant1 = 8'd142; a_mant2 = 8'd151; a_mant3 = 8'd75;
b_mant0 = 8'd217; b_mant1 = 8'd239; b_mant2 = 8'd129; b_mant3 = 8'd184;
a_exp0 = 10'd907; a_exp1 = 10'd243; a_exp2 = 10'd977; a_exp3 = 10'd268;
b_exp0 = 10'd199; b_exp1 = 10'd377; b_exp2 = 10'd270; b_exp3 = 10'd745;
a_sign0 = 4'd0; a_sign1 = 4'd0; a_sign2 = 4'd2; a_sign3 = 4'd9;
b_sign0 = 4'd14; b_sign1 = 4'd9; b_sign2 = 4'd2; b_sign3 = 4'd4;
@(posedge clk_i);
a_mant0 = 8'd145; a_mant1 = 8'd56; a_mant2 = 8'd61; a_mant3 = 8'd103;
b_mant0 = 8'd192; b_mant1 = 8'd75; b_mant2 = 8'd20; b_mant3 = 8'd96;
a_exp0 = 10'd862; a_exp1 = 10'd578; a_exp2 = 10'd116; a_exp3 = 10'd500;
b_exp0 = 10'd470; b_exp1 = 10'd386; b_exp2 = 10'd591; b_exp3 = 10'd492;
a_sign0 = 4'd10; a_sign1 = 4'd15; a_sign2 = 4'd4; a_sign3 = 4'd1;
b_sign0 = 4'd13; b_sign1 = 4'd7; b_sign2 = 4'd1; b_sign3 = 4'd13;
@(posedge clk_i);
a_mant0 = 8'd231; a_mant1 = 8'd12; a_mant2 = 8'd226; a_mant3 = 8'd175;
b_mant0 = 8'd237; b_mant1 = 8'd108; b_mant2 = 8'd181; b_mant3 = 8'd164;
a_exp0 = 10'd22; a_exp1 = 10'd582; a_exp2 = 10'd469; a_exp3 = 10'd175;
b_exp0 = 10'd117; b_exp1 = 10'd74; b_exp2 = 10'd670; b_exp3 = 10'd824;
a_sign0 = 4'd7; a_sign1 = 4'd0; a_sign2 = 4'd14; a_sign3 = 4'd7;
b_sign0 = 4'd15; b_sign1 = 4'd4; b_sign2 = 4'd10; b_sign3 = 4'd13;
@(posedge clk_i);
shared_exps0 = 8'd130;
shared_exps1 = 8'd141;
rstn = 0;
@(posedge clk_i);
rstn = 1;
a_mant0 = 8'd76; a_mant1 = 8'd233; a_mant2 = 8'd189; a_mant3 = 8'd158;
b_mant0 = 8'd75; b_mant1 = 8'd133; b_mant2 = 8'd122; b_mant3 = 8'd9;
a_exp0 = 10'd1016; a_exp1 = 10'd461; a_exp2 = 10'd214; a_exp3 = 10'd743;
b_exp0 = 10'd423; b_exp1 = 10'd435; b_exp2 = 10'd988; b_exp3 = 10'd183;
a_sign0 = 4'd5; a_sign1 = 4'd16; a_sign2 = 4'd13; a_sign3 = 4'd0;
b_sign0 = 4'd6; b_sign1 = 4'd15; b_sign2 = 4'd1; b_sign3 = 4'd3;
@(posedge clk_i);
a_mant0 = 8'd84; a_mant1 = 8'd104; a_mant2 = 8'd204; a_mant3 = 8'd119;
b_mant0 = 8'd246; b_mant1 = 8'd63; b_mant2 = 8'd150; b_mant3 = 8'd90;
a_exp0 = 10'd981; a_exp1 = 10'd887; a_exp2 = 10'd247; a_exp3 = 10'd102;
b_exp0 = 10'd839; b_exp1 = 10'd279; b_exp2 = 10'd446; b_exp3 = 10'd886;
a_sign0 = 4'd13; a_sign1 = 4'd5; a_sign2 = 4'd9; a_sign3 = 4'd11;
b_sign0 = 4'd0; b_sign1 = 4'd12; b_sign2 = 4'd13; b_sign3 = 4'd7;
@(posedge clk_i);
a_mant0 = 8'd191; a_mant1 = 8'd0; a_mant2 = 8'd145; a_mant3 = 8'd253;
b_mant0 = 8'd163; b_mant1 = 8'd202; b_mant2 = 8'd25; b_mant3 = 8'd81;
a_exp0 = 10'd671; a_exp1 = 10'd982; a_exp2 = 10'd460; a_exp3 = 10'd224;
b_exp0 = 10'd582; b_exp1 = 10'd990; b_exp2 = 10'd418; b_exp3 = 10'd471;
a_sign0 = 4'd8; a_sign1 = 4'd9; a_sign2 = 4'd3; a_sign3 = 4'd0;
b_sign0 = 4'd16; b_sign1 = 4'd0; b_sign2 = 4'd16; b_sign3 = 4'd9;
@(posedge clk_i);
a_mant0 = 8'd133; a_mant1 = 8'd29; a_mant2 = 8'd153; a_mant3 = 8'd12;
b_mant0 = 8'd41; b_mant1 = 8'd151; b_mant2 = 8'd90; b_mant3 = 8'd66;
a_exp0 = 10'd39; a_exp1 = 10'd374; a_exp2 = 10'd714; a_exp3 = 10'd711;
b_exp0 = 10'd617; b_exp1 = 10'd648; b_exp2 = 10'd244; b_exp3 = 10'd449;
a_sign0 = 4'd13; a_sign1 = 4'd4; a_sign2 = 4'd3; a_sign3 = 4'd5;
b_sign0 = 4'd11; b_sign1 = 4'd1; b_sign2 = 4'd16; b_sign3 = 4'd12;
@(posedge clk_i);
a_mant0 = 8'd222; a_mant1 = 8'd23; a_mant2 = 8'd155; a_mant3 = 8'd234;
b_mant0 = 8'd37; b_mant1 = 8'd199; b_mant2 = 8'd63; b_mant3 = 8'd36;
a_exp0 = 10'd505; a_exp1 = 10'd470; a_exp2 = 10'd919; a_exp3 = 10'd597;
b_exp0 = 10'd476; b_exp1 = 10'd299; b_exp2 = 10'd997; b_exp3 = 10'd390;
a_sign0 = 4'd0; a_sign1 = 4'd8; a_sign2 = 4'd11; a_sign3 = 4'd8;
b_sign0 = 4'd2; b_sign1 = 4'd11; b_sign2 = 4'd10; b_sign3 = 4'd4;
@(posedge clk_i);
a_mant0 = 8'd84; a_mant1 = 8'd45; a_mant2 = 8'd16; a_mant3 = 8'd113;
b_mant0 = 8'd195; b_mant1 = 8'd153; b_mant2 = 8'd175; b_mant3 = 8'd73;
a_exp0 = 10'd1011; a_exp1 = 10'd388; a_exp2 = 10'd822; a_exp3 = 10'd2;
b_exp0 = 10'd156; b_exp1 = 10'd229; b_exp2 = 10'd923; b_exp3 = 10'd186;
a_sign0 = 4'd13; a_sign1 = 4'd15; a_sign2 = 4'd4; a_sign3 = 4'd4;
b_sign0 = 4'd5; b_sign1 = 4'd9; b_sign2 = 4'd2; b_sign3 = 4'd0;
@(posedge clk_i);
a_mant0 = 8'd243; a_mant1 = 8'd204; a_mant2 = 8'd61; a_mant3 = 8'd22;
b_mant0 = 8'd19; b_mant1 = 8'd12; b_mant2 = 8'd56; b_mant3 = 8'd199;
a_exp0 = 10'd964; a_exp1 = 10'd450; a_exp2 = 10'd267; a_exp3 = 10'd340;
b_exp0 = 10'd989; b_exp1 = 10'd2; b_exp2 = 10'd907; b_exp3 = 10'd576;
a_sign0 = 4'd14; a_sign1 = 4'd13; a_sign2 = 4'd2; a_sign3 = 4'd2;
b_sign0 = 4'd15; b_sign1 = 4'd6; b_sign2 = 4'd6; b_sign3 = 4'd0;
@(posedge clk_i);
shared_exps0 = 8'd134;
shared_exps1 = 8'd114;
a_mant0 = 8'd72; a_mant1 = 8'd236; a_mant2 = 8'd87; a_mant3 = 8'd42;
b_mant0 = 8'd228; b_mant1 = 8'd12; b_mant2 = 8'd255; b_mant3 = 8'd205;
a_exp0 = 10'd74; a_exp1 = 10'd936; a_exp2 = 10'd738; a_exp3 = 10'd665;
b_exp0 = 10'd545; b_exp1 = 10'd532; b_exp2 = 10'd469; b_exp3 = 10'd860;
a_sign0 = 4'd0; a_sign1 = 4'd5; a_sign2 = 4'd5; a_sign3 = 4'd9;
b_sign0 = 4'd6; b_sign1 = 4'd13; b_sign2 = 4'd1; b_sign3 = 4'd13;
@(posedge clk_i);
a_mant0 = 8'd85; a_mant1 = 8'd96; a_mant2 = 8'd129; a_mant3 = 8'd255;
b_mant0 = 8'd172; b_mant1 = 8'd13; b_mant2 = 8'd130; b_mant3 = 8'd42;
a_exp0 = 10'd272; a_exp1 = 10'd36; a_exp2 = 10'd320; a_exp3 = 10'd664;
b_exp0 = 10'd232; b_exp1 = 10'd815; b_exp2 = 10'd182; b_exp3 = 10'd267;
a_sign0 = 4'd3; a_sign1 = 4'd15; a_sign2 = 4'd7; a_sign3 = 4'd4;
b_sign0 = 4'd5; b_sign1 = 4'd6; b_sign2 = 4'd4; b_sign3 = 4'd5;
@(posedge clk_i);
a_mant0 = 8'd117; a_mant1 = 8'd144; a_mant2 = 8'd204; a_mant3 = 8'd252;
b_mant0 = 8'd204; b_mant1 = 8'd30; b_mant2 = 8'd92; b_mant3 = 8'd196;
a_exp0 = 10'd401; a_exp1 = 10'd889; a_exp2 = 10'd508; a_exp3 = 10'd1000;
b_exp0 = 10'd409; b_exp1 = 10'd687; b_exp2 = 10'd139; b_exp3 = 10'd710;
a_sign0 = 4'd5; a_sign1 = 4'd15; a_sign2 = 4'd3; a_sign3 = 4'd12;
b_sign0 = 4'd16; b_sign1 = 4'd1; b_sign2 = 4'd2; b_sign3 = 4'd13;
@(posedge clk_i);
a_mant0 = 8'd166; a_mant1 = 8'd179; a_mant2 = 8'd141; a_mant3 = 8'd105;
b_mant0 = 8'd19; b_mant1 = 8'd45; b_mant2 = 8'd186; b_mant3 = 8'd110;
a_exp0 = 10'd528; a_exp1 = 10'd920; a_exp2 = 10'd250; a_exp3 = 10'd856;
b_exp0 = 10'd16; b_exp1 = 10'd662; b_exp2 = 10'd56; b_exp3 = 10'd193;
a_sign0 = 4'd11; a_sign1 = 4'd3; a_sign2 = 4'd1; a_sign3 = 4'd5;
b_sign0 = 4'd11; b_sign1 = 4'd1; b_sign2 = 4'd0; b_sign3 = 4'd9;
@(posedge clk_i);
a_mant0 = 8'd148; a_mant1 = 8'd40; a_mant2 = 8'd130; a_mant3 = 8'd226;
b_mant0 = 8'd186; b_mant1 = 8'd156; b_mant2 = 8'd135; b_mant3 = 8'd81;
a_exp0 = 10'd743; a_exp1 = 10'd367; a_exp2 = 10'd925; a_exp3 = 10'd92;
b_exp0 = 10'd986; b_exp1 = 10'd577; b_exp2 = 10'd839; b_exp3 = 10'd879;
a_sign0 = 4'd5; a_sign1 = 4'd1; a_sign2 = 4'd7; a_sign3 = 4'd6;
b_sign0 = 4'd4; b_sign1 = 4'd10; b_sign2 = 4'd7; b_sign3 = 4'd5;
@(posedge clk_i);
a_mant0 = 8'd156; a_mant1 = 8'd197; a_mant2 = 8'd44; a_mant3 = 8'd95;
b_mant0 = 8'd187; b_mant1 = 8'd14; b_mant2 = 8'd218; b_mant3 = 8'd47;
a_exp0 = 10'd695; a_exp1 = 10'd733; a_exp2 = 10'd675; a_exp3 = 10'd227;
b_exp0 = 10'd134; b_exp1 = 10'd17; b_exp2 = 10'd114; b_exp3 = 10'd696;
a_sign0 = 4'd11; a_sign1 = 4'd14; a_sign2 = 4'd6; a_sign3 = 4'd15;
b_sign0 = 4'd1; b_sign1 = 4'd16; b_sign2 = 4'd13; b_sign3 = 4'd0;
@(posedge clk_i);
a_mant0 = 8'd93; a_mant1 = 8'd68; a_mant2 = 8'd225; a_mant3 = 8'd209;
b_mant0 = 8'd51; b_mant1 = 8'd15; b_mant2 = 8'd133; b_mant3 = 8'd227;
a_exp0 = 10'd387; a_exp1 = 10'd481; a_exp2 = 10'd91; a_exp3 = 10'd26;
b_exp0 = 10'd200; b_exp1 = 10'd34; b_exp2 = 10'd426; b_exp3 = 10'd576;
a_sign0 = 4'd15; a_sign1 = 4'd11; a_sign2 = 4'd7; a_sign3 = 4'd0;
b_sign0 = 4'd6; b_sign1 = 4'd9; b_sign2 = 4'd8; b_sign3 = 4'd1;
@(posedge clk_i);
a_mant0 = 8'd223; a_mant1 = 8'd180; a_mant2 = 8'd230; a_mant3 = 8'd157;
b_mant0 = 8'd91; b_mant1 = 8'd178; b_mant2 = 8'd42; b_mant3 = 8'd78;
a_exp0 = 10'd363; a_exp1 = 10'd428; a_exp2 = 10'd724; a_exp3 = 10'd496;
b_exp0 = 10'd987; b_exp1 = 10'd340; b_exp2 = 10'd115; b_exp3 = 10'd1011;
a_sign0 = 4'd5; a_sign1 = 4'd5; a_sign2 = 4'd7; a_sign3 = 4'd5;
b_sign0 = 4'd5; b_sign1 = 4'd11; b_sign2 = 4'd1; b_sign3 = 4'd14;
@(posedge clk_i);
shared_exps0 = 8'd116;
shared_exps1 = 8'd138;
a_mant0 = 8'd180; a_mant1 = 8'd209; a_mant2 = 8'd28; a_mant3 = 8'd8;
b_mant0 = 8'd44; b_mant1 = 8'd32; b_mant2 = 8'd203; b_mant3 = 8'd241;
a_exp0 = 10'd4; a_exp1 = 10'd828; a_exp2 = 10'd75; a_exp3 = 10'd263;
b_exp0 = 10'd764; b_exp1 = 10'd587; b_exp2 = 10'd55; b_exp3 = 10'd1011;
a_sign0 = 4'd12; a_sign1 = 4'd7; a_sign2 = 4'd5; a_sign3 = 4'd15;
b_sign0 = 4'd5; b_sign1 = 4'd4; b_sign2 = 4'd11; b_sign3 = 4'd16;
@(posedge clk_i);
a_mant0 = 8'd165; a_mant1 = 8'd138; a_mant2 = 8'd172; a_mant3 = 8'd127;
b_mant0 = 8'd192; b_mant1 = 8'd217; b_mant2 = 8'd126; b_mant3 = 8'd39;
a_exp0 = 10'd952; a_exp1 = 10'd76; a_exp2 = 10'd866; a_exp3 = 10'd109;
b_exp0 = 10'd29; b_exp1 = 10'd493; b_exp2 = 10'd326; b_exp3 = 10'd188;
a_sign0 = 4'd7; a_sign1 = 4'd12; a_sign2 = 4'd13; a_sign3 = 4'd8;
b_sign0 = 4'd0; b_sign1 = 4'd11; b_sign2 = 4'd10; b_sign3 = 4'd11;
@(posedge clk_i);
a_mant0 = 8'd152; a_mant1 = 8'd36; a_mant2 = 8'd183; a_mant3 = 8'd33;
b_mant0 = 8'd112; b_mant1 = 8'd152; b_mant2 = 8'd203; b_mant3 = 8'd214;
a_exp0 = 10'd317; a_exp1 = 10'd150; a_exp2 = 10'd479; a_exp3 = 10'd671;
b_exp0 = 10'd319; b_exp1 = 10'd438; b_exp2 = 10'd791; b_exp3 = 10'd190;
a_sign0 = 4'd9; a_sign1 = 4'd3; a_sign2 = 4'd16; a_sign3 = 4'd12;
b_sign0 = 4'd0; b_sign1 = 4'd10; b_sign2 = 4'd3; b_sign3 = 4'd14;
@(posedge clk_i);
a_mant0 = 8'd105; a_mant1 = 8'd142; a_mant2 = 8'd106; a_mant3 = 8'd115;
b_mant0 = 8'd80; b_mant1 = 8'd104; b_mant2 = 8'd34; b_mant3 = 8'd89;
a_exp0 = 10'd131; a_exp1 = 10'd310; a_exp2 = 10'd335; a_exp3 = 10'd60;
b_exp0 = 10'd608; b_exp1 = 10'd677; b_exp2 = 10'd1002; b_exp3 = 10'd645;
a_sign0 = 4'd5; a_sign1 = 4'd5; a_sign2 = 4'd13; a_sign3 = 4'd7;
b_sign0 = 4'd2; b_sign1 = 4'd9; b_sign2 = 4'd4; b_sign3 = 4'd9;
@(posedge clk_i);
a_mant0 = 8'd100; a_mant1 = 8'd70; a_mant2 = 8'd45; a_mant3 = 8'd250;
b_mant0 = 8'd233; b_mant1 = 8'd113; b_mant2 = 8'd200; b_mant3 = 8'd95;
a_exp0 = 10'd99; a_exp1 = 10'd514; a_exp2 = 10'd253; a_exp3 = 10'd225;
b_exp0 = 10'd316; b_exp1 = 10'd20; b_exp2 = 10'd777; b_exp3 = 10'd443;
a_sign0 = 4'd0; a_sign1 = 4'd6; a_sign2 = 4'd11; a_sign3 = 4'd7;
b_sign0 = 4'd16; b_sign1 = 4'd7; b_sign2 = 4'd16; b_sign3 = 4'd3;
@(posedge clk_i);
a_mant0 = 8'd100; a_mant1 = 8'd7; a_mant2 = 8'd72; a_mant3 = 8'd189;
b_mant0 = 8'd110; b_mant1 = 8'd139; b_mant2 = 8'd34; b_mant3 = 8'd169;
a_exp0 = 10'd316; a_exp1 = 10'd353; a_exp2 = 10'd742; a_exp3 = 10'd238;
b_exp0 = 10'd679; b_exp1 = 10'd50; b_exp2 = 10'd736; b_exp3 = 10'd177;
a_sign0 = 4'd10; a_sign1 = 4'd10; a_sign2 = 4'd0; a_sign3 = 4'd4;
b_sign0 = 4'd15; b_sign1 = 4'd13; b_sign2 = 4'd9; b_sign3 = 4'd15;
@(posedge clk_i);
a_mant0 = 8'd149; a_mant1 = 8'd129; a_mant2 = 8'd66; a_mant3 = 8'd218;
b_mant0 = 8'd154; b_mant1 = 8'd252; b_mant2 = 8'd189; b_mant3 = 8'd109;
a_exp0 = 10'd970; a_exp1 = 10'd301; a_exp2 = 10'd505; a_exp3 = 10'd212;
b_exp0 = 10'd862; b_exp1 = 10'd699; b_exp2 = 10'd379; b_exp3 = 10'd673;
a_sign0 = 4'd2; a_sign1 = 4'd6; a_sign2 = 4'd4; a_sign3 = 4'd2;
b_sign0 = 4'd7; b_sign1 = 4'd3; b_sign2 = 4'd16; b_sign3 = 4'd12;
@(posedge clk_i);
a_mant0 = 8'd114; a_mant1 = 8'd68; a_mant2 = 8'd45; a_mant3 = 8'd10;
b_mant0 = 8'd136; b_mant1 = 8'd153; b_mant2 = 8'd95; b_mant3 = 8'd104;
a_exp0 = 10'd173; a_exp1 = 10'd422; a_exp2 = 10'd425; a_exp3 = 10'd763;
b_exp0 = 10'd712; b_exp1 = 10'd595; b_exp2 = 10'd590; b_exp3 = 10'd248;
a_sign0 = 4'd8; a_sign1 = 4'd10; a_sign2 = 4'd7; a_sign3 = 4'd0;
b_sign0 = 4'd9; b_sign1 = 4'd3; b_sign2 = 4'd13; b_sign3 = 4'd3;
@(posedge clk_i);
shared_exps0 = 8'd118;
shared_exps1 = 8'd151;
a_mant0 = 8'd120; a_mant1 = 8'd167; a_mant2 = 8'd108; a_mant3 = 8'd103;
b_mant0 = 8'd99; b_mant1 = 8'd251; b_mant2 = 8'd18; b_mant3 = 8'd241;
a_exp0 = 10'd981; a_exp1 = 10'd769; a_exp2 = 10'd987; a_exp3 = 10'd658;
b_exp0 = 10'd999; b_exp1 = 10'd824; b_exp2 = 10'd114; b_exp3 = 10'd357;
a_sign0 = 4'd9; a_sign1 = 4'd4; a_sign2 = 4'd2; a_sign3 = 4'd13;
b_sign0 = 4'd9; b_sign1 = 4'd12; b_sign2 = 4'd9; b_sign3 = 4'd10;
@(posedge clk_i);
a_mant0 = 8'd148; a_mant1 = 8'd59; a_mant2 = 8'd170; a_mant3 = 8'd136;
b_mant0 = 8'd63; b_mant1 = 8'd42; b_mant2 = 8'd61; b_mant3 = 8'd89;
a_exp0 = 10'd215; a_exp1 = 10'd830; a_exp2 = 10'd267; a_exp3 = 10'd567;
b_exp0 = 10'd354; b_exp1 = 10'd1005; b_exp2 = 10'd454; b_exp3 = 10'd349;
a_sign0 = 4'd8; a_sign1 = 4'd14; a_sign2 = 4'd13; a_sign3 = 4'd8;
b_sign0 = 4'd4; b_sign1 = 4'd4; b_sign2 = 4'd7; b_sign3 = 4'd11;
@(posedge clk_i);
a_mant0 = 8'd90; a_mant1 = 8'd17; a_mant2 = 8'd81; a_mant3 = 8'd172;
b_mant0 = 8'd148; b_mant1 = 8'd254; b_mant2 = 8'd98; b_mant3 = 8'd111;
a_exp0 = 10'd880; a_exp1 = 10'd770; a_exp2 = 10'd518; a_exp3 = 10'd741;
b_exp0 = 10'd733; b_exp1 = 10'd442; b_exp2 = 10'd804; b_exp3 = 10'd481;
a_sign0 = 4'd2; a_sign1 = 4'd13; a_sign2 = 4'd16; a_sign3 = 4'd7;
b_sign0 = 4'd7; b_sign1 = 4'd8; b_sign2 = 4'd4; b_sign3 = 4'd12;
@(posedge clk_i);
a_mant0 = 8'd49; a_mant1 = 8'd188; a_mant2 = 8'd240; a_mant3 = 8'd188;
b_mant0 = 8'd95; b_mant1 = 8'd19; b_mant2 = 8'd88; b_mant3 = 8'd23;
a_exp0 = 10'd171; a_exp1 = 10'd59; a_exp2 = 10'd665; a_exp3 = 10'd992;
b_exp0 = 10'd621; b_exp1 = 10'd245; b_exp2 = 10'd699; b_exp3 = 10'd107;
a_sign0 = 4'd15; a_sign1 = 4'd12; a_sign2 = 4'd2; a_sign3 = 4'd4;
b_sign0 = 4'd0; b_sign1 = 4'd8; b_sign2 = 4'd6; b_sign3 = 4'd1;
@(posedge clk_i);
a_mant0 = 8'd123; a_mant1 = 8'd38; a_mant2 = 8'd28; a_mant3 = 8'd78;
b_mant0 = 8'd145; b_mant1 = 8'd156; b_mant2 = 8'd99; b_mant3 = 8'd239;
a_exp0 = 10'd765; a_exp1 = 10'd87; a_exp2 = 10'd911; a_exp3 = 10'd772;
b_exp0 = 10'd726; b_exp1 = 10'd461; b_exp2 = 10'd821; b_exp3 = 10'd927;
a_sign0 = 4'd16; a_sign1 = 4'd8; a_sign2 = 4'd4; a_sign3 = 4'd8;
b_sign0 = 4'd5; b_sign1 = 4'd4; b_sign2 = 4'd6; b_sign3 = 4'd14;
@(posedge clk_i);
a_mant0 = 8'd113; a_mant1 = 8'd102; a_mant2 = 8'd169; a_mant3 = 8'd79;
b_mant0 = 8'd50; b_mant1 = 8'd170; b_mant2 = 8'd243; b_mant3 = 8'd128;
a_exp0 = 10'd637; a_exp1 = 10'd858; a_exp2 = 10'd469; a_exp3 = 10'd99;
b_exp0 = 10'd603; b_exp1 = 10'd118; b_exp2 = 10'd462; b_exp3 = 10'd624;
a_sign0 = 4'd5; a_sign1 = 4'd6; a_sign2 = 4'd4; a_sign3 = 4'd7;
b_sign0 = 4'd2; b_sign1 = 4'd15; b_sign2 = 4'd5; b_sign3 = 4'd12;
@(posedge clk_i);
a_mant0 = 8'd86; a_mant1 = 8'd245; a_mant2 = 8'd138; a_mant3 = 8'd109;
b_mant0 = 8'd137; b_mant1 = 8'd182; b_mant2 = 8'd167; b_mant3 = 8'd185;
a_exp0 = 10'd640; a_exp1 = 10'd775; a_exp2 = 10'd134; a_exp3 = 10'd572;
b_exp0 = 10'd585; b_exp1 = 10'd737; b_exp2 = 10'd303; b_exp3 = 10'd405;
a_sign0 = 4'd10; a_sign1 = 4'd13; a_sign2 = 4'd12; a_sign3 = 4'd0;
b_sign0 = 4'd8; b_sign1 = 4'd3; b_sign2 = 4'd10; b_sign3 = 4'd1;
@(posedge clk_i);
a_mant0 = 8'd61; a_mant1 = 8'd48; a_mant2 = 8'd152; a_mant3 = 8'd180;
b_mant0 = 8'd210; b_mant1 = 8'd191; b_mant2 = 8'd48; b_mant3 = 8'd174;
a_exp0 = 10'd620; a_exp1 = 10'd526; a_exp2 = 10'd985; a_exp3 = 10'd925;
b_exp0 = 10'd425; b_exp1 = 10'd1009; b_exp2 = 10'd112; b_exp3 = 10'd362;
a_sign0 = 4'd0; a_sign1 = 4'd16; a_sign2 = 4'd13; a_sign3 = 4'd16;
b_sign0 = 4'd14; b_sign1 = 4'd5; b_sign2 = 4'd1; b_sign3 = 4'd13;
@(posedge clk_i);
shared_exps0 = 8'd123;
shared_exps1 = 8'd125;
rstn = 0;
@(posedge clk_i);
rstn = 1;
a_mant0 = 8'd68; a_mant1 = 8'd205; a_mant2 = 8'd154; a_mant3 = 8'd58;
b_mant0 = 8'd158; b_mant1 = 8'd163; b_mant2 = 8'd9; b_mant3 = 8'd192;
a_exp0 = 10'd542; a_exp1 = 10'd126; a_exp2 = 10'd64; a_exp3 = 10'd862;
b_exp0 = 10'd875; b_exp1 = 10'd371; b_exp2 = 10'd588; b_exp3 = 10'd333;
a_sign0 = 4'd8; a_sign1 = 4'd6; a_sign2 = 4'd12; a_sign3 = 4'd16;
b_sign0 = 4'd13; b_sign1 = 4'd14; b_sign2 = 4'd0; b_sign3 = 4'd7;
@(posedge clk_i);
a_mant0 = 8'd210; a_mant1 = 8'd37; a_mant2 = 8'd40; a_mant3 = 8'd242;
b_mant0 = 8'd238; b_mant1 = 8'd173; b_mant2 = 8'd244; b_mant3 = 8'd230;
a_exp0 = 10'd803; a_exp1 = 10'd260; a_exp2 = 10'd982; a_exp3 = 10'd57;
b_exp0 = 10'd36; b_exp1 = 10'd769; b_exp2 = 10'd908; b_exp3 = 10'd359;
a_sign0 = 4'd11; a_sign1 = 4'd3; a_sign2 = 4'd11; a_sign3 = 4'd2;
b_sign0 = 4'd1; b_sign1 = 4'd5; b_sign2 = 4'd1; b_sign3 = 4'd7;
@(posedge clk_i);
a_mant0 = 8'd150; a_mant1 = 8'd255; a_mant2 = 8'd195; a_mant3 = 8'd12;
b_mant0 = 8'd178; b_mant1 = 8'd137; b_mant2 = 8'd114; b_mant3 = 8'd144;
a_exp0 = 10'd463; a_exp1 = 10'd349; a_exp2 = 10'd250; a_exp3 = 10'd470;
b_exp0 = 10'd98; b_exp1 = 10'd48; b_exp2 = 10'd504; b_exp3 = 10'd129;
a_sign0 = 4'd12; a_sign1 = 4'd13; a_sign2 = 4'd4; a_sign3 = 4'd12;
b_sign0 = 4'd5; b_sign1 = 4'd9; b_sign2 = 4'd13; b_sign3 = 4'd9;
@(posedge clk_i);
a_mant0 = 8'd107; a_mant1 = 8'd144; a_mant2 = 8'd1; a_mant3 = 8'd201;
b_mant0 = 8'd210; b_mant1 = 8'd34; b_mant2 = 8'd94; b_mant3 = 8'd134;
a_exp0 = 10'd15; a_exp1 = 10'd226; a_exp2 = 10'd526; a_exp3 = 10'd336;
b_exp0 = 10'd996; b_exp1 = 10'd670; b_exp2 = 10'd314; b_exp3 = 10'd591;
a_sign0 = 4'd16; a_sign1 = 4'd8; a_sign2 = 4'd9; a_sign3 = 4'd3;
b_sign0 = 4'd11; b_sign1 = 4'd13; b_sign2 = 4'd15; b_sign3 = 4'd10;
@(posedge clk_i);
a_mant0 = 8'd4; a_mant1 = 8'd63; a_mant2 = 8'd205; a_mant3 = 8'd241;
b_mant0 = 8'd39; b_mant1 = 8'd228; b_mant2 = 8'd14; b_mant3 = 8'd85;
a_exp0 = 10'd895; a_exp1 = 10'd580; a_exp2 = 10'd696; a_exp3 = 10'd365;
b_exp0 = 10'd899; b_exp1 = 10'd769; b_exp2 = 10'd729; b_exp3 = 10'd821;
a_sign0 = 4'd10; a_sign1 = 4'd0; a_sign2 = 4'd1; a_sign3 = 4'd0;
b_sign0 = 4'd10; b_sign1 = 4'd6; b_sign2 = 4'd6; b_sign3 = 4'd3;
@(posedge clk_i);
a_mant0 = 8'd185; a_mant1 = 8'd73; a_mant2 = 8'd28; a_mant3 = 8'd253;
b_mant0 = 8'd211; b_mant1 = 8'd91; b_mant2 = 8'd26; b_mant3 = 8'd218;
a_exp0 = 10'd420; a_exp1 = 10'd473; a_exp2 = 10'd495; a_exp3 = 10'd972;
b_exp0 = 10'd458; b_exp1 = 10'd131; b_exp2 = 10'd950; b_exp3 = 10'd264;
a_sign0 = 4'd11; a_sign1 = 4'd14; a_sign2 = 4'd13; a_sign3 = 4'd11;
b_sign0 = 4'd1; b_sign1 = 4'd2; b_sign2 = 4'd16; b_sign3 = 4'd12;
@(posedge clk_i);
a_mant0 = 8'd77; a_mant1 = 8'd62; a_mant2 = 8'd64; a_mant3 = 8'd200;
b_mant0 = 8'd92; b_mant1 = 8'd83; b_mant2 = 8'd255; b_mant3 = 8'd127;
a_exp0 = 10'd974; a_exp1 = 10'd451; a_exp2 = 10'd1012; a_exp3 = 10'd528;
b_exp0 = 10'd16; b_exp1 = 10'd632; b_exp2 = 10'd148; b_exp3 = 10'd862;
a_sign0 = 4'd10; a_sign1 = 4'd12; a_sign2 = 4'd12; a_sign3 = 4'd0;
b_sign0 = 4'd0; b_sign1 = 4'd15; b_sign2 = 4'd12; b_sign3 = 4'd16;
@(posedge clk_i);
shared_exps0 = 8'd158;
shared_exps1 = 8'd126;
a_mant0 = 8'd220; a_mant1 = 8'd185; a_mant2 = 8'd184; a_mant3 = 8'd115;
b_mant0 = 8'd66; b_mant1 = 8'd140; b_mant2 = 8'd2; b_mant3 = 8'd86;
a_exp0 = 10'd730; a_exp1 = 10'd672; a_exp2 = 10'd426; a_exp3 = 10'd381;
b_exp0 = 10'd175; b_exp1 = 10'd50; b_exp2 = 10'd611; b_exp3 = 10'd110;
a_sign0 = 4'd2; a_sign1 = 4'd14; a_sign2 = 4'd0; a_sign3 = 4'd6;
b_sign0 = 4'd6; b_sign1 = 4'd15; b_sign2 = 4'd10; b_sign3 = 4'd9;
@(posedge clk_i);
a_mant0 = 8'd72; a_mant1 = 8'd176; a_mant2 = 8'd14; a_mant3 = 8'd75;
b_mant0 = 8'd69; b_mant1 = 8'd28; b_mant2 = 8'd182; b_mant3 = 8'd88;
a_exp0 = 10'd139; a_exp1 = 10'd483; a_exp2 = 10'd955; a_exp3 = 10'd831;
b_exp0 = 10'd193; b_exp1 = 10'd456; b_exp2 = 10'd818; b_exp3 = 10'd424;
a_sign0 = 4'd4; a_sign1 = 4'd7; a_sign2 = 4'd4; a_sign3 = 4'd15;
b_sign0 = 4'd6; b_sign1 = 4'd15; b_sign2 = 4'd15; b_sign3 = 4'd16;
@(posedge clk_i);
a_mant0 = 8'd250; a_mant1 = 8'd47; a_mant2 = 8'd40; a_mant3 = 8'd209;
b_mant0 = 8'd38; b_mant1 = 8'd145; b_mant2 = 8'd207; b_mant3 = 8'd211;
a_exp0 = 10'd662; a_exp1 = 10'd383; a_exp2 = 10'd681; a_exp3 = 10'd669;
b_exp0 = 10'd570; b_exp1 = 10'd129; b_exp2 = 10'd797; b_exp3 = 10'd927;
a_sign0 = 4'd5; a_sign1 = 4'd7; a_sign2 = 4'd11; a_sign3 = 4'd7;
b_sign0 = 4'd16; b_sign1 = 4'd13; b_sign2 = 4'd3; b_sign3 = 4'd11;
@(posedge clk_i);
a_mant0 = 8'd223; a_mant1 = 8'd23; a_mant2 = 8'd78; a_mant3 = 8'd10;
b_mant0 = 8'd217; b_mant1 = 8'd167; b_mant2 = 8'd175; b_mant3 = 8'd137;
a_exp0 = 10'd645; a_exp1 = 10'd874; a_exp2 = 10'd262; a_exp3 = 10'd24;
b_exp0 = 10'd781; b_exp1 = 10'd68; b_exp2 = 10'd616; b_exp3 = 10'd972;
a_sign0 = 4'd12; a_sign1 = 4'd13; a_sign2 = 4'd13; a_sign3 = 4'd5;
b_sign0 = 4'd9; b_sign1 = 4'd14; b_sign2 = 4'd13; b_sign3 = 4'd2;
@(posedge clk_i);
a_mant0 = 8'd138; a_mant1 = 8'd17; a_mant2 = 8'd94; a_mant3 = 8'd180;
b_mant0 = 8'd120; b_mant1 = 8'd113; b_mant2 = 8'd223; b_mant3 = 8'd107;
a_exp0 = 10'd336; a_exp1 = 10'd132; a_exp2 = 10'd477; a_exp3 = 10'd976;
b_exp0 = 10'd68; b_exp1 = 10'd384; b_exp2 = 10'd741; b_exp3 = 10'd470;
a_sign0 = 4'd0; a_sign1 = 4'd2; a_sign2 = 4'd7; a_sign3 = 4'd15;
b_sign0 = 4'd2; b_sign1 = 4'd8; b_sign2 = 4'd8; b_sign3 = 4'd6;
@(posedge clk_i);
a_mant0 = 8'd214; a_mant1 = 8'd143; a_mant2 = 8'd135; a_mant3 = 8'd207;
b_mant0 = 8'd99; b_mant1 = 8'd239; b_mant2 = 8'd34; b_mant3 = 8'd100;
a_exp0 = 10'd872; a_exp1 = 10'd297; a_exp2 = 10'd146; a_exp3 = 10'd1007;
b_exp0 = 10'd332; b_exp1 = 10'd614; b_exp2 = 10'd504; b_exp3 = 10'd640;
a_sign0 = 4'd1; a_sign1 = 4'd12; a_sign2 = 4'd13; a_sign3 = 4'd5;
b_sign0 = 4'd7; b_sign1 = 4'd13; b_sign2 = 4'd13; b_sign3 = 4'd6;
@(posedge clk_i);
a_mant0 = 8'd163; a_mant1 = 8'd195; a_mant2 = 8'd61; a_mant3 = 8'd222;
b_mant0 = 8'd30; b_mant1 = 8'd243; b_mant2 = 8'd12; b_mant3 = 8'd22;
a_exp0 = 10'd988; a_exp1 = 10'd174; a_exp2 = 10'd297; a_exp3 = 10'd654;
b_exp0 = 10'd277; b_exp1 = 10'd897; b_exp2 = 10'd200; b_exp3 = 10'd353;
a_sign0 = 4'd5; a_sign1 = 4'd5; a_sign2 = 4'd5; a_sign3 = 4'd15;
b_sign0 = 4'd10; b_sign1 = 4'd2; b_sign2 = 4'd0; b_sign3 = 4'd7;
@(posedge clk_i);
a_mant0 = 8'd102; a_mant1 = 8'd229; a_mant2 = 8'd239; a_mant3 = 8'd69;
b_mant0 = 8'd90; b_mant1 = 8'd59; b_mant2 = 8'd46; b_mant3 = 8'd2;
a_exp0 = 10'd321; a_exp1 = 10'd666; a_exp2 = 10'd133; a_exp3 = 10'd14;
b_exp0 = 10'd145; b_exp1 = 10'd888; b_exp2 = 10'd698; b_exp3 = 10'd524;
a_sign0 = 4'd6; a_sign1 = 4'd13; a_sign2 = 4'd11; a_sign3 = 4'd4;
b_sign0 = 4'd2; b_sign1 = 4'd0; b_sign2 = 4'd6; b_sign3 = 4'd0;
@(posedge clk_i);
shared_exps0 = 8'd125;
shared_exps1 = 8'd130;
a_mant0 = 8'd40; a_mant1 = 8'd68; a_mant2 = 8'd128; a_mant3 = 8'd48;
b_mant0 = 8'd186; b_mant1 = 8'd218; b_mant2 = 8'd48; b_mant3 = 8'd196;
a_exp0 = 10'd610; a_exp1 = 10'd227; a_exp2 = 10'd381; a_exp3 = 10'd67;
b_exp0 = 10'd261; b_exp1 = 10'd681; b_exp2 = 10'd740; b_exp3 = 10'd811;
a_sign0 = 4'd7; a_sign1 = 4'd8; a_sign2 = 4'd14; a_sign3 = 4'd5;
b_sign0 = 4'd1; b_sign1 = 4'd6; b_sign2 = 4'd13; b_sign3 = 4'd16;
@(posedge clk_i);
a_mant0 = 8'd253; a_mant1 = 8'd205; a_mant2 = 8'd253; a_mant3 = 8'd94;
b_mant0 = 8'd56; b_mant1 = 8'd91; b_mant2 = 8'd151; b_mant3 = 8'd37;
a_exp0 = 10'd870; a_exp1 = 10'd875; a_exp2 = 10'd747; a_exp3 = 10'd762;
b_exp0 = 10'd691; b_exp1 = 10'd655; b_exp2 = 10'd314; b_exp3 = 10'd904;
a_sign0 = 4'd14; a_sign1 = 4'd11; a_sign2 = 4'd14; a_sign3 = 4'd7;
b_sign0 = 4'd12; b_sign1 = 4'd13; b_sign2 = 4'd12; b_sign3 = 4'd14;
@(posedge clk_i);
a_mant0 = 8'd136; a_mant1 = 8'd152; a_mant2 = 8'd112; a_mant3 = 8'd58;
b_mant0 = 8'd22; b_mant1 = 8'd103; b_mant2 = 8'd106; b_mant3 = 8'd39;
a_exp0 = 10'd736; a_exp1 = 10'd840; a_exp2 = 10'd15; a_exp3 = 10'd886;
b_exp0 = 10'd256; b_exp1 = 10'd678; b_exp2 = 10'd357; b_exp3 = 10'd1006;
a_sign0 = 4'd10; a_sign1 = 4'd5; a_sign2 = 4'd11; a_sign3 = 4'd9;
b_sign0 = 4'd15; b_sign1 = 4'd3; b_sign2 = 4'd12; b_sign3 = 4'd5;
@(posedge clk_i);
a_mant0 = 8'd238; a_mant1 = 8'd111; a_mant2 = 8'd18; a_mant3 = 8'd38;
b_mant0 = 8'd165; b_mant1 = 8'd154; b_mant2 = 8'd17; b_mant3 = 8'd114;
a_exp0 = 10'd398; a_exp1 = 10'd348; a_exp2 = 10'd898; a_exp3 = 10'd626;
b_exp0 = 10'd362; b_exp1 = 10'd889; b_exp2 = 10'd734; b_exp3 = 10'd463;
a_sign0 = 4'd7; a_sign1 = 4'd15; a_sign2 = 4'd8; a_sign3 = 4'd11;
b_sign0 = 4'd12; b_sign1 = 4'd15; b_sign2 = 4'd6; b_sign3 = 4'd7;
@(posedge clk_i);
a_mant0 = 8'd211; a_mant1 = 8'd81; a_mant2 = 8'd252; a_mant3 = 8'd68;
b_mant0 = 8'd114; b_mant1 = 8'd239; b_mant2 = 8'd239; b_mant3 = 8'd131;
a_exp0 = 10'd432; a_exp1 = 10'd784; a_exp2 = 10'd371; a_exp3 = 10'd385;
b_exp0 = 10'd903; b_exp1 = 10'd633; b_exp2 = 10'd126; b_exp3 = 10'd584;
a_sign0 = 4'd16; a_sign1 = 4'd6; a_sign2 = 4'd10; a_sign3 = 4'd2;
b_sign0 = 4'd16; b_sign1 = 4'd10; b_sign2 = 4'd16; b_sign3 = 4'd15;
@(posedge clk_i);
a_mant0 = 8'd53; a_mant1 = 8'd59; a_mant2 = 8'd205; a_mant3 = 8'd246;
b_mant0 = 8'd1; b_mant1 = 8'd169; b_mant2 = 8'd74; b_mant3 = 8'd194;
a_exp0 = 10'd104; a_exp1 = 10'd189; a_exp2 = 10'd573; a_exp3 = 10'd502;
b_exp0 = 10'd211; b_exp1 = 10'd614; b_exp2 = 10'd328; b_exp3 = 10'd160;
a_sign0 = 4'd7; a_sign1 = 4'd15; a_sign2 = 4'd7; a_sign3 = 4'd13;
b_sign0 = 4'd14; b_sign1 = 4'd15; b_sign2 = 4'd4; b_sign3 = 4'd7;
@(posedge clk_i);
a_mant0 = 8'd208; a_mant1 = 8'd24; a_mant2 = 8'd12; a_mant3 = 8'd139;
b_mant0 = 8'd205; b_mant1 = 8'd148; b_mant2 = 8'd232; b_mant3 = 8'd153;
a_exp0 = 10'd985; a_exp1 = 10'd702; a_exp2 = 10'd664; a_exp3 = 10'd672;
b_exp0 = 10'd914; b_exp1 = 10'd573; b_exp2 = 10'd717; b_exp3 = 10'd728;
a_sign0 = 4'd3; a_sign1 = 4'd15; a_sign2 = 4'd6; a_sign3 = 4'd15;
b_sign0 = 4'd5; b_sign1 = 4'd0; b_sign2 = 4'd16; b_sign3 = 4'd3;
@(posedge clk_i);
a_mant0 = 8'd231; a_mant1 = 8'd248; a_mant2 = 8'd21; a_mant3 = 8'd128;
b_mant0 = 8'd255; b_mant1 = 8'd169; b_mant2 = 8'd178; b_mant3 = 8'd165;
a_exp0 = 10'd81; a_exp1 = 10'd922; a_exp2 = 10'd411; a_exp3 = 10'd467;
b_exp0 = 10'd358; b_exp1 = 10'd540; b_exp2 = 10'd708; b_exp3 = 10'd236;
a_sign0 = 4'd0; a_sign1 = 4'd16; a_sign2 = 4'd5; a_sign3 = 4'd13;
b_sign0 = 4'd7; b_sign1 = 4'd2; b_sign2 = 4'd6; b_sign3 = 4'd6;
@(posedge clk_i);
shared_exps0 = 8'd139;
shared_exps1 = 8'd126;
a_mant0 = 8'd248; a_mant1 = 8'd172; a_mant2 = 8'd198; a_mant3 = 8'd156;
b_mant0 = 8'd236; b_mant1 = 8'd242; b_mant2 = 8'd237; b_mant3 = 8'd71;
a_exp0 = 10'd949; a_exp1 = 10'd368; a_exp2 = 10'd697; a_exp3 = 10'd1013;
b_exp0 = 10'd980; b_exp1 = 10'd189; b_exp2 = 10'd622; b_exp3 = 10'd370;
a_sign0 = 4'd11; a_sign1 = 4'd5; a_sign2 = 4'd12; a_sign3 = 4'd14;
b_sign0 = 4'd5; b_sign1 = 4'd1; b_sign2 = 4'd14; b_sign3 = 4'd1;
@(posedge clk_i);
a_mant0 = 8'd251; a_mant1 = 8'd246; a_mant2 = 8'd20; a_mant3 = 8'd61;
b_mant0 = 8'd12; b_mant1 = 8'd116; b_mant2 = 8'd47; b_mant3 = 8'd101;
a_exp0 = 10'd696; a_exp1 = 10'd107; a_exp2 = 10'd256; a_exp3 = 10'd60;
b_exp0 = 10'd562; b_exp1 = 10'd272; b_exp2 = 10'd471; b_exp3 = 10'd385;
a_sign0 = 4'd8; a_sign1 = 4'd15; a_sign2 = 4'd13; a_sign3 = 4'd4;
b_sign0 = 4'd15; b_sign1 = 4'd8; b_sign2 = 4'd0; b_sign3 = 4'd15;
@(posedge clk_i);
a_mant0 = 8'd96; a_mant1 = 8'd101; a_mant2 = 8'd191; a_mant3 = 8'd78;
b_mant0 = 8'd11; b_mant1 = 8'd2; b_mant2 = 8'd174; b_mant3 = 8'd123;
a_exp0 = 10'd207; a_exp1 = 10'd159; a_exp2 = 10'd369; a_exp3 = 10'd916;
b_exp0 = 10'd878; b_exp1 = 10'd901; b_exp2 = 10'd343; b_exp3 = 10'd153;
a_sign0 = 4'd8; a_sign1 = 4'd13; a_sign2 = 4'd16; a_sign3 = 4'd9;
b_sign0 = 4'd2; b_sign1 = 4'd3; b_sign2 = 4'd15; b_sign3 = 4'd1;
@(posedge clk_i);
a_mant0 = 8'd58; a_mant1 = 8'd248; a_mant2 = 8'd16; a_mant3 = 8'd188;
b_mant0 = 8'd55; b_mant1 = 8'd121; b_mant2 = 8'd83; b_mant3 = 8'd225;
a_exp0 = 10'd52; a_exp1 = 10'd813; a_exp2 = 10'd518; a_exp3 = 10'd201;
b_exp0 = 10'd873; b_exp1 = 10'd383; b_exp2 = 10'd830; b_exp3 = 10'd862;
a_sign0 = 4'd4; a_sign1 = 4'd14; a_sign2 = 4'd14; a_sign3 = 4'd6;
b_sign0 = 4'd14; b_sign1 = 4'd5; b_sign2 = 4'd8; b_sign3 = 4'd6;
@(posedge clk_i);
a_mant0 = 8'd174; a_mant1 = 8'd250; a_mant2 = 8'd7; a_mant3 = 8'd188;
b_mant0 = 8'd104; b_mant1 = 8'd50; b_mant2 = 8'd112; b_mant3 = 8'd84;
a_exp0 = 10'd539; a_exp1 = 10'd462; a_exp2 = 10'd60; a_exp3 = 10'd687;
b_exp0 = 10'd951; b_exp1 = 10'd520; b_exp2 = 10'd588; b_exp3 = 10'd592;
a_sign0 = 4'd4; a_sign1 = 4'd12; a_sign2 = 4'd8; a_sign3 = 4'd13;
b_sign0 = 4'd7; b_sign1 = 4'd16; b_sign2 = 4'd14; b_sign3 = 4'd5;
@(posedge clk_i);
a_mant0 = 8'd135; a_mant1 = 8'd201; a_mant2 = 8'd170; a_mant3 = 8'd192;
b_mant0 = 8'd250; b_mant1 = 8'd96; b_mant2 = 8'd199; b_mant3 = 8'd189;
a_exp0 = 10'd72; a_exp1 = 10'd122; a_exp2 = 10'd585; a_exp3 = 10'd799;
b_exp0 = 10'd191; b_exp1 = 10'd80; b_exp2 = 10'd642; b_exp3 = 10'd128;
a_sign0 = 4'd0; a_sign1 = 4'd16; a_sign2 = 4'd12; a_sign3 = 4'd8;
b_sign0 = 4'd15; b_sign1 = 4'd4; b_sign2 = 4'd9; b_sign3 = 4'd5;
@(posedge clk_i);
a_mant0 = 8'd50; a_mant1 = 8'd37; a_mant2 = 8'd232; a_mant3 = 8'd184;
b_mant0 = 8'd202; b_mant1 = 8'd47; b_mant2 = 8'd18; b_mant3 = 8'd104;
a_exp0 = 10'd759; a_exp1 = 10'd348; a_exp2 = 10'd225; a_exp3 = 10'd763;
b_exp0 = 10'd968; b_exp1 = 10'd1006; b_exp2 = 10'd493; b_exp3 = 10'd429;
a_sign0 = 4'd8; a_sign1 = 4'd10; a_sign2 = 4'd10; a_sign3 = 4'd12;
b_sign0 = 4'd7; b_sign1 = 4'd11; b_sign2 = 4'd14; b_sign3 = 4'd16;
@(posedge clk_i);
a_mant0 = 8'd202; a_mant1 = 8'd82; a_mant2 = 8'd175; a_mant3 = 8'd172;
b_mant0 = 8'd91; b_mant1 = 8'd74; b_mant2 = 8'd182; b_mant3 = 8'd37;
a_exp0 = 10'd823; a_exp1 = 10'd352; a_exp2 = 10'd340; a_exp3 = 10'd348;
b_exp0 = 10'd741; b_exp1 = 10'd24; b_exp2 = 10'd270; b_exp3 = 10'd123;
a_sign0 = 4'd4; a_sign1 = 4'd12; a_sign2 = 4'd0; a_sign3 = 4'd1;
b_sign0 = 4'd9; b_sign1 = 4'd1; b_sign2 = 4'd0; b_sign3 = 4'd7;
@(posedge clk_i);
shared_exps0 = 8'd121;
shared_exps1 = 8'd125;
rstn = 0;
@(posedge clk_i);
rstn = 1;
a_mant0 = 8'd166; a_mant1 = 8'd36; a_mant2 = 8'd149; a_mant3 = 8'd115;
b_mant0 = 8'd1; b_mant1 = 8'd81; b_mant2 = 8'd225; b_mant3 = 8'd73;
a_exp0 = 10'd506; a_exp1 = 10'd987; a_exp2 = 10'd612; a_exp3 = 10'd1014;
b_exp0 = 10'd341; b_exp1 = 10'd654; b_exp2 = 10'd657; b_exp3 = 10'd822;
a_sign0 = 4'd0; a_sign1 = 4'd5; a_sign2 = 4'd2; a_sign3 = 4'd10;
b_sign0 = 4'd3; b_sign1 = 4'd9; b_sign2 = 4'd3; b_sign3 = 4'd16;
@(posedge clk_i);
a_mant0 = 8'd148; a_mant1 = 8'd118; a_mant2 = 8'd214; a_mant3 = 8'd76;
b_mant0 = 8'd51; b_mant1 = 8'd110; b_mant2 = 8'd97; b_mant3 = 8'd126;
a_exp0 = 10'd551; a_exp1 = 10'd697; a_exp2 = 10'd178; a_exp3 = 10'd346;
b_exp0 = 10'd292; b_exp1 = 10'd316; b_exp2 = 10'd544; b_exp3 = 10'd452;
a_sign0 = 4'd10; a_sign1 = 4'd10; a_sign2 = 4'd10; a_sign3 = 4'd9;
b_sign0 = 4'd5; b_sign1 = 4'd0; b_sign2 = 4'd10; b_sign3 = 4'd5;
@(posedge clk_i);
a_mant0 = 8'd6; a_mant1 = 8'd163; a_mant2 = 8'd54; a_mant3 = 8'd57;
b_mant0 = 8'd237; b_mant1 = 8'd13; b_mant2 = 8'd40; b_mant3 = 8'd168;
a_exp0 = 10'd461; a_exp1 = 10'd238; a_exp2 = 10'd111; a_exp3 = 10'd22;
b_exp0 = 10'd565; b_exp1 = 10'd774; b_exp2 = 10'd152; b_exp3 = 10'd187;
a_sign0 = 4'd1; a_sign1 = 4'd7; a_sign2 = 4'd5; a_sign3 = 4'd1;
b_sign0 = 4'd13; b_sign1 = 4'd15; b_sign2 = 4'd12; b_sign3 = 4'd8;
@(posedge clk_i);
a_mant0 = 8'd112; a_mant1 = 8'd210; a_mant2 = 8'd78; a_mant3 = 8'd41;
b_mant0 = 8'd133; b_mant1 = 8'd1; b_mant2 = 8'd107; b_mant3 = 8'd249;
a_exp0 = 10'd845; a_exp1 = 10'd851; a_exp2 = 10'd889; a_exp3 = 10'd930;
b_exp0 = 10'd856; b_exp1 = 10'd72; b_exp2 = 10'd762; b_exp3 = 10'd38;
a_sign0 = 4'd6; a_sign1 = 4'd3; a_sign2 = 4'd10; a_sign3 = 4'd5;
b_sign0 = 4'd16; b_sign1 = 4'd13; b_sign2 = 4'd2; b_sign3 = 4'd10;
@(posedge clk_i);
a_mant0 = 8'd116; a_mant1 = 8'd222; a_mant2 = 8'd27; a_mant3 = 8'd44;
b_mant0 = 8'd185; b_mant1 = 8'd238; b_mant2 = 8'd161; b_mant3 = 8'd109;
a_exp0 = 10'd559; a_exp1 = 10'd160; a_exp2 = 10'd7; a_exp3 = 10'd890;
b_exp0 = 10'd138; b_exp1 = 10'd400; b_exp2 = 10'd149; b_exp3 = 10'd3;
a_sign0 = 4'd16; a_sign1 = 4'd15; a_sign2 = 4'd16; a_sign3 = 4'd12;
b_sign0 = 4'd0; b_sign1 = 4'd3; b_sign2 = 4'd4; b_sign3 = 4'd3;
@(posedge clk_i);
a_mant0 = 8'd135; a_mant1 = 8'd72; a_mant2 = 8'd216; a_mant3 = 8'd242;
b_mant0 = 8'd54; b_mant1 = 8'd107; b_mant2 = 8'd112; b_mant3 = 8'd88;
a_exp0 = 10'd797; a_exp1 = 10'd123; a_exp2 = 10'd658; a_exp3 = 10'd302;
b_exp0 = 10'd872; b_exp1 = 10'd219; b_exp2 = 10'd859; b_exp3 = 10'd871;
a_sign0 = 4'd14; a_sign1 = 4'd9; a_sign2 = 4'd12; a_sign3 = 4'd10;
b_sign0 = 4'd11; b_sign1 = 4'd5; b_sign2 = 4'd0; b_sign3 = 4'd11;
@(posedge clk_i);
a_mant0 = 8'd187; a_mant1 = 8'd102; a_mant2 = 8'd202; a_mant3 = 8'd91;
b_mant0 = 8'd164; b_mant1 = 8'd246; b_mant2 = 8'd166; b_mant3 = 8'd165;
a_exp0 = 10'd609; a_exp1 = 10'd436; a_exp2 = 10'd84; a_exp3 = 10'd813;
b_exp0 = 10'd358; b_exp1 = 10'd35; b_exp2 = 10'd1019; b_exp3 = 10'd750;
a_sign0 = 4'd9; a_sign1 = 4'd5; a_sign2 = 4'd1; a_sign3 = 4'd3;
b_sign0 = 4'd0; b_sign1 = 4'd3; b_sign2 = 4'd4; b_sign3 = 4'd14;
@(posedge clk_i);
shared_exps0 = 8'd111;
shared_exps1 = 8'd134;
a_mant0 = 8'd233; a_mant1 = 8'd111; a_mant2 = 8'd155; a_mant3 = 8'd41;
b_mant0 = 8'd53; b_mant1 = 8'd71; b_mant2 = 8'd55; b_mant3 = 8'd222;
a_exp0 = 10'd974; a_exp1 = 10'd755; a_exp2 = 10'd560; a_exp3 = 10'd306;
b_exp0 = 10'd17; b_exp1 = 10'd124; b_exp2 = 10'd341; b_exp3 = 10'd597;
a_sign0 = 4'd7; a_sign1 = 4'd4; a_sign2 = 4'd13; a_sign3 = 4'd7;
b_sign0 = 4'd10; b_sign1 = 4'd4; b_sign2 = 4'd7; b_sign3 = 4'd15;
@(posedge clk_i);
a_mant0 = 8'd201; a_mant1 = 8'd42; a_mant2 = 8'd109; a_mant3 = 8'd52;
b_mant0 = 8'd85; b_mant1 = 8'd47; b_mant2 = 8'd159; b_mant3 = 8'd150;
a_exp0 = 10'd821; a_exp1 = 10'd568; a_exp2 = 10'd138; a_exp3 = 10'd764;
b_exp0 = 10'd349; b_exp1 = 10'd457; b_exp2 = 10'd692; b_exp3 = 10'd147;
a_sign0 = 4'd7; a_sign1 = 4'd5; a_sign2 = 4'd16; a_sign3 = 4'd8;
b_sign0 = 4'd7; b_sign1 = 4'd5; b_sign2 = 4'd0; b_sign3 = 4'd14;
@(posedge clk_i);
a_mant0 = 8'd107; a_mant1 = 8'd102; a_mant2 = 8'd226; a_mant3 = 8'd88;
b_mant0 = 8'd151; b_mant1 = 8'd127; b_mant2 = 8'd149; b_mant3 = 8'd54;
a_exp0 = 10'd205; a_exp1 = 10'd261; a_exp2 = 10'd47; a_exp3 = 10'd39;
b_exp0 = 10'd177; b_exp1 = 10'd231; b_exp2 = 10'd17; b_exp3 = 10'd377;
a_sign0 = 4'd0; a_sign1 = 4'd12; a_sign2 = 4'd5; a_sign3 = 4'd15;
b_sign0 = 4'd3; b_sign1 = 4'd16; b_sign2 = 4'd4; b_sign3 = 4'd10;
@(posedge clk_i);
a_mant0 = 8'd1; a_mant1 = 8'd192; a_mant2 = 8'd67; a_mant3 = 8'd74;
b_mant0 = 8'd116; b_mant1 = 8'd99; b_mant2 = 8'd173; b_mant3 = 8'd76;
a_exp0 = 10'd423; a_exp1 = 10'd466; a_exp2 = 10'd390; a_exp3 = 10'd942;
b_exp0 = 10'd725; b_exp1 = 10'd483; b_exp2 = 10'd654; b_exp3 = 10'd998;
a_sign0 = 4'd2; a_sign1 = 4'd2; a_sign2 = 4'd2; a_sign3 = 4'd14;
b_sign0 = 4'd3; b_sign1 = 4'd8; b_sign2 = 4'd11; b_sign3 = 4'd7;
@(posedge clk_i);
a_mant0 = 8'd62; a_mant1 = 8'd196; a_mant2 = 8'd90; a_mant3 = 8'd23;
b_mant0 = 8'd184; b_mant1 = 8'd14; b_mant2 = 8'd157; b_mant3 = 8'd59;
a_exp0 = 10'd246; a_exp1 = 10'd903; a_exp2 = 10'd42; a_exp3 = 10'd326;
b_exp0 = 10'd239; b_exp1 = 10'd835; b_exp2 = 10'd78; b_exp3 = 10'd28;
a_sign0 = 4'd8; a_sign1 = 4'd1; a_sign2 = 4'd12; a_sign3 = 4'd12;
b_sign0 = 4'd8; b_sign1 = 4'd12; b_sign2 = 4'd13; b_sign3 = 4'd13;
@(posedge clk_i);
a_mant0 = 8'd113; a_mant1 = 8'd164; a_mant2 = 8'd239; a_mant3 = 8'd50;
b_mant0 = 8'd83; b_mant1 = 8'd191; b_mant2 = 8'd61; b_mant3 = 8'd239;
a_exp0 = 10'd130; a_exp1 = 10'd103; a_exp2 = 10'd656; a_exp3 = 10'd72;
b_exp0 = 10'd919; b_exp1 = 10'd740; b_exp2 = 10'd1002; b_exp3 = 10'd437;
a_sign0 = 4'd12; a_sign1 = 4'd3; a_sign2 = 4'd13; a_sign3 = 4'd7;
b_sign0 = 4'd16; b_sign1 = 4'd2; b_sign2 = 4'd6; b_sign3 = 4'd14;
@(posedge clk_i);
a_mant0 = 8'd69; a_mant1 = 8'd113; a_mant2 = 8'd185; a_mant3 = 8'd0;
b_mant0 = 8'd182; b_mant1 = 8'd44; b_mant2 = 8'd61; b_mant3 = 8'd114;
a_exp0 = 10'd372; a_exp1 = 10'd136; a_exp2 = 10'd40; a_exp3 = 10'd773;
b_exp0 = 10'd401; b_exp1 = 10'd49; b_exp2 = 10'd585; b_exp3 = 10'd325;
a_sign0 = 4'd0; a_sign1 = 4'd15; a_sign2 = 4'd6; a_sign3 = 4'd11;
b_sign0 = 4'd3; b_sign1 = 4'd8; b_sign2 = 4'd3; b_sign3 = 4'd15;
@(posedge clk_i);
a_mant0 = 8'd91; a_mant1 = 8'd227; a_mant2 = 8'd244; a_mant3 = 8'd219;
b_mant0 = 8'd211; b_mant1 = 8'd132; b_mant2 = 8'd4; b_mant3 = 8'd175;
a_exp0 = 10'd60; a_exp1 = 10'd857; a_exp2 = 10'd191; a_exp3 = 10'd377;
b_exp0 = 10'd109; b_exp1 = 10'd286; b_exp2 = 10'd774; b_exp3 = 10'd982;
a_sign0 = 4'd6; a_sign1 = 4'd13; a_sign2 = 4'd11; a_sign3 = 4'd2;
b_sign0 = 4'd2; b_sign1 = 4'd12; b_sign2 = 4'd6; b_sign3 = 4'd12;
@(posedge clk_i);
shared_exps0 = 8'd105;
shared_exps1 = 8'd138;
a_mant0 = 8'd20; a_mant1 = 8'd15; a_mant2 = 8'd155; a_mant3 = 8'd89;
b_mant0 = 8'd238; b_mant1 = 8'd79; b_mant2 = 8'd37; b_mant3 = 8'd81;
a_exp0 = 10'd492; a_exp1 = 10'd1016; a_exp2 = 10'd207; a_exp3 = 10'd363;
b_exp0 = 10'd219; b_exp1 = 10'd202; b_exp2 = 10'd199; b_exp3 = 10'd832;
a_sign0 = 4'd11; a_sign1 = 4'd15; a_sign2 = 4'd1; a_sign3 = 4'd2;
b_sign0 = 4'd11; b_sign1 = 4'd13; b_sign2 = 4'd0; b_sign3 = 4'd12;
@(posedge clk_i);
a_mant0 = 8'd106; a_mant1 = 8'd178; a_mant2 = 8'd51; a_mant3 = 8'd126;
b_mant0 = 8'd195; b_mant1 = 8'd128; b_mant2 = 8'd168; b_mant3 = 8'd209;
a_exp0 = 10'd976; a_exp1 = 10'd34; a_exp2 = 10'd186; a_exp3 = 10'd1015;
b_exp0 = 10'd318; b_exp1 = 10'd725; b_exp2 = 10'd1001; b_exp3 = 10'd984;
a_sign0 = 4'd6; a_sign1 = 4'd8; a_sign2 = 4'd8; a_sign3 = 4'd13;
b_sign0 = 4'd5; b_sign1 = 4'd6; b_sign2 = 4'd5; b_sign3 = 4'd16;
@(posedge clk_i);
a_mant0 = 8'd55; a_mant1 = 8'd170; a_mant2 = 8'd63; a_mant3 = 8'd212;
b_mant0 = 8'd253; b_mant1 = 8'd46; b_mant2 = 8'd202; b_mant3 = 8'd153;
a_exp0 = 10'd109; a_exp1 = 10'd738; a_exp2 = 10'd210; a_exp3 = 10'd80;
b_exp0 = 10'd652; b_exp1 = 10'd278; b_exp2 = 10'd818; b_exp3 = 10'd253;
a_sign0 = 4'd11; a_sign1 = 4'd14; a_sign2 = 4'd9; a_sign3 = 4'd4;
b_sign0 = 4'd12; b_sign1 = 4'd3; b_sign2 = 4'd10; b_sign3 = 4'd13;
@(posedge clk_i);
a_mant0 = 8'd210; a_mant1 = 8'd166; a_mant2 = 8'd152; a_mant3 = 8'd238;
b_mant0 = 8'd243; b_mant1 = 8'd135; b_mant2 = 8'd86; b_mant3 = 8'd130;
a_exp0 = 10'd582; a_exp1 = 10'd419; a_exp2 = 10'd591; a_exp3 = 10'd189;
b_exp0 = 10'd463; b_exp1 = 10'd187; b_exp2 = 10'd112; b_exp3 = 10'd308;
a_sign0 = 4'd6; a_sign1 = 4'd14; a_sign2 = 4'd9; a_sign3 = 4'd9;
b_sign0 = 4'd10; b_sign1 = 4'd5; b_sign2 = 4'd15; b_sign3 = 4'd5;
@(posedge clk_i);
a_mant0 = 8'd150; a_mant1 = 8'd83; a_mant2 = 8'd146; a_mant3 = 8'd76;
b_mant0 = 8'd5; b_mant1 = 8'd46; b_mant2 = 8'd30; b_mant3 = 8'd1;
a_exp0 = 10'd281; a_exp1 = 10'd113; a_exp2 = 10'd815; a_exp3 = 10'd298;
b_exp0 = 10'd67; b_exp1 = 10'd104; b_exp2 = 10'd814; b_exp3 = 10'd515;
a_sign0 = 4'd1; a_sign1 = 4'd10; a_sign2 = 4'd10; a_sign3 = 4'd4;
b_sign0 = 4'd16; b_sign1 = 4'd12; b_sign2 = 4'd10; b_sign3 = 4'd2;
@(posedge clk_i);
a_mant0 = 8'd148; a_mant1 = 8'd77; a_mant2 = 8'd68; a_mant3 = 8'd177;
b_mant0 = 8'd64; b_mant1 = 8'd134; b_mant2 = 8'd126; b_mant3 = 8'd222;
a_exp0 = 10'd800; a_exp1 = 10'd827; a_exp2 = 10'd256; a_exp3 = 10'd546;
b_exp0 = 10'd423; b_exp1 = 10'd421; b_exp2 = 10'd976; b_exp3 = 10'd155;
a_sign0 = 4'd15; a_sign1 = 4'd0; a_sign2 = 4'd8; a_sign3 = 4'd7;
b_sign0 = 4'd10; b_sign1 = 4'd8; b_sign2 = 4'd16; b_sign3 = 4'd14;
@(posedge clk_i);
a_mant0 = 8'd137; a_mant1 = 8'd59; a_mant2 = 8'd165; a_mant3 = 8'd144;
b_mant0 = 8'd192; b_mant1 = 8'd23; b_mant2 = 8'd88; b_mant3 = 8'd120;
a_exp0 = 10'd217; a_exp1 = 10'd455; a_exp2 = 10'd996; a_exp3 = 10'd276;
b_exp0 = 10'd182; b_exp1 = 10'd862; b_exp2 = 10'd503; b_exp3 = 10'd741;
a_sign0 = 4'd2; a_sign1 = 4'd15; a_sign2 = 4'd4; a_sign3 = 4'd2;
b_sign0 = 4'd12; b_sign1 = 4'd15; b_sign2 = 4'd13; b_sign3 = 4'd5;
@(posedge clk_i);
a_mant0 = 8'd220; a_mant1 = 8'd44; a_mant2 = 8'd10; a_mant3 = 8'd92;
b_mant0 = 8'd73; b_mant1 = 8'd153; b_mant2 = 8'd61; b_mant3 = 8'd11;
a_exp0 = 10'd701; a_exp1 = 10'd728; a_exp2 = 10'd283; a_exp3 = 10'd662;
b_exp0 = 10'd121; b_exp1 = 10'd617; b_exp2 = 10'd913; b_exp3 = 10'd578;
a_sign0 = 4'd8; a_sign1 = 4'd12; a_sign2 = 4'd3; a_sign3 = 4'd2;
b_sign0 = 4'd5; b_sign1 = 4'd16; b_sign2 = 4'd15; b_sign3 = 4'd14;
@(posedge clk_i);
shared_exps0 = 8'd124;
shared_exps1 = 8'd120;
a_mant0 = 8'd9; a_mant1 = 8'd150; a_mant2 = 8'd10; a_mant3 = 8'd51;
b_mant0 = 8'd78; b_mant1 = 8'd160; b_mant2 = 8'd12; b_mant3 = 8'd24;
a_exp0 = 10'd850; a_exp1 = 10'd824; a_exp2 = 10'd531; a_exp3 = 10'd131;
b_exp0 = 10'd317; b_exp1 = 10'd554; b_exp2 = 10'd864; b_exp3 = 10'd790;
a_sign0 = 4'd4; a_sign1 = 4'd15; a_sign2 = 4'd10; a_sign3 = 4'd8;
b_sign0 = 4'd12; b_sign1 = 4'd12; b_sign2 = 4'd6; b_sign3 = 4'd2;
@(posedge clk_i);
a_mant0 = 8'd41; a_mant1 = 8'd92; a_mant2 = 8'd25; a_mant3 = 8'd149;
b_mant0 = 8'd21; b_mant1 = 8'd194; b_mant2 = 8'd178; b_mant3 = 8'd24;
a_exp0 = 10'd876; a_exp1 = 10'd610; a_exp2 = 10'd846; a_exp3 = 10'd37;
b_exp0 = 10'd60; b_exp1 = 10'd975; b_exp2 = 10'd248; b_exp3 = 10'd353;
a_sign0 = 4'd11; a_sign1 = 4'd15; a_sign2 = 4'd2; a_sign3 = 4'd1;
b_sign0 = 4'd14; b_sign1 = 4'd0; b_sign2 = 4'd5; b_sign3 = 4'd12;
@(posedge clk_i);
a_mant0 = 8'd234; a_mant1 = 8'd71; a_mant2 = 8'd196; a_mant3 = 8'd9;
b_mant0 = 8'd93; b_mant1 = 8'd226; b_mant2 = 8'd252; b_mant3 = 8'd34;
a_exp0 = 10'd764; a_exp1 = 10'd306; a_exp2 = 10'd93; a_exp3 = 10'd134;
b_exp0 = 10'd443; b_exp1 = 10'd869; b_exp2 = 10'd910; b_exp3 = 10'd818;
a_sign0 = 4'd10; a_sign1 = 4'd0; a_sign2 = 4'd1; a_sign3 = 4'd2;
b_sign0 = 4'd13; b_sign1 = 4'd10; b_sign2 = 4'd13; b_sign3 = 4'd11;
@(posedge clk_i);
a_mant0 = 8'd19; a_mant1 = 8'd159; a_mant2 = 8'd198; a_mant3 = 8'd243;
b_mant0 = 8'd163; b_mant1 = 8'd200; b_mant2 = 8'd240; b_mant3 = 8'd152;
a_exp0 = 10'd0; a_exp1 = 10'd627; a_exp2 = 10'd315; a_exp3 = 10'd363;
b_exp0 = 10'd303; b_exp1 = 10'd611; b_exp2 = 10'd664; b_exp3 = 10'd424;
a_sign0 = 4'd1; a_sign1 = 4'd9; a_sign2 = 4'd6; a_sign3 = 4'd13;
b_sign0 = 4'd3; b_sign1 = 4'd1; b_sign2 = 4'd5; b_sign3 = 4'd13;
@(posedge clk_i);
a_mant0 = 8'd100; a_mant1 = 8'd253; a_mant2 = 8'd32; a_mant3 = 8'd53;
b_mant0 = 8'd155; b_mant1 = 8'd204; b_mant2 = 8'd195; b_mant3 = 8'd97;
a_exp0 = 10'd163; a_exp1 = 10'd441; a_exp2 = 10'd658; a_exp3 = 10'd400;
b_exp0 = 10'd841; b_exp1 = 10'd224; b_exp2 = 10'd127; b_exp3 = 10'd393;
a_sign0 = 4'd12; a_sign1 = 4'd4; a_sign2 = 4'd4; a_sign3 = 4'd10;
b_sign0 = 4'd9; b_sign1 = 4'd9; b_sign2 = 4'd5; b_sign3 = 4'd2;
@(posedge clk_i);
a_mant0 = 8'd251; a_mant1 = 8'd34; a_mant2 = 8'd193; a_mant3 = 8'd229;
b_mant0 = 8'd134; b_mant1 = 8'd153; b_mant2 = 8'd174; b_mant3 = 8'd121;
a_exp0 = 10'd742; a_exp1 = 10'd984; a_exp2 = 10'd736; a_exp3 = 10'd564;
b_exp0 = 10'd470; b_exp1 = 10'd28; b_exp2 = 10'd298; b_exp3 = 10'd397;
a_sign0 = 4'd7; a_sign1 = 4'd9; a_sign2 = 4'd8; a_sign3 = 4'd13;
b_sign0 = 4'd0; b_sign1 = 4'd12; b_sign2 = 4'd8; b_sign3 = 4'd12;
@(posedge clk_i);
a_mant0 = 8'd207; a_mant1 = 8'd237; a_mant2 = 8'd197; a_mant3 = 8'd133;
b_mant0 = 8'd228; b_mant1 = 8'd61; b_mant2 = 8'd34; b_mant3 = 8'd198;
a_exp0 = 10'd686; a_exp1 = 10'd465; a_exp2 = 10'd490; a_exp3 = 10'd293;
b_exp0 = 10'd721; b_exp1 = 10'd410; b_exp2 = 10'd336; b_exp3 = 10'd659;
a_sign0 = 4'd16; a_sign1 = 4'd5; a_sign2 = 4'd16; a_sign3 = 4'd12;
b_sign0 = 4'd1; b_sign1 = 4'd6; b_sign2 = 4'd7; b_sign3 = 4'd11;
@(posedge clk_i);
a_mant0 = 8'd72; a_mant1 = 8'd11; a_mant2 = 8'd2; a_mant3 = 8'd169;
b_mant0 = 8'd107; b_mant1 = 8'd228; b_mant2 = 8'd72; b_mant3 = 8'd63;
a_exp0 = 10'd430; a_exp1 = 10'd550; a_exp2 = 10'd981; a_exp3 = 10'd365;
b_exp0 = 10'd531; b_exp1 = 10'd95; b_exp2 = 10'd604; b_exp3 = 10'd73;
a_sign0 = 4'd10; a_sign1 = 4'd2; a_sign2 = 4'd10; a_sign3 = 4'd11;
b_sign0 = 4'd4; b_sign1 = 4'd8; b_sign2 = 4'd12; b_sign3 = 4'd16;
@(posedge clk_i);
shared_exps0 = 8'd144;
shared_exps1 = 8'd141;
rstn = 0;
@(posedge clk_i);
rstn = 1;
a_mant0 = 8'd99; a_mant1 = 8'd153; a_mant2 = 8'd28; a_mant3 = 8'd17;
b_mant0 = 8'd90; b_mant1 = 8'd219; b_mant2 = 8'd154; b_mant3 = 8'd232;
a_exp0 = 10'd948; a_exp1 = 10'd561; a_exp2 = 10'd165; a_exp3 = 10'd45;
b_exp0 = 10'd819; b_exp1 = 10'd702; b_exp2 = 10'd792; b_exp3 = 10'd952;
a_sign0 = 4'd12; a_sign1 = 4'd14; a_sign2 = 4'd3; a_sign3 = 4'd5;
b_sign0 = 4'd3; b_sign1 = 4'd10; b_sign2 = 4'd12; b_sign3 = 4'd13;
@(posedge clk_i);
a_mant0 = 8'd106; a_mant1 = 8'd147; a_mant2 = 8'd226; a_mant3 = 8'd246;
b_mant0 = 8'd121; b_mant1 = 8'd212; b_mant2 = 8'd196; b_mant3 = 8'd65;
a_exp0 = 10'd426; a_exp1 = 10'd441; a_exp2 = 10'd730; a_exp3 = 10'd477;
b_exp0 = 10'd330; b_exp1 = 10'd440; b_exp2 = 10'd591; b_exp3 = 10'd999;
a_sign0 = 4'd13; a_sign1 = 4'd9; a_sign2 = 4'd4; a_sign3 = 4'd15;
b_sign0 = 4'd0; b_sign1 = 4'd6; b_sign2 = 4'd15; b_sign3 = 4'd0;
@(posedge clk_i);
a_mant0 = 8'd164; a_mant1 = 8'd122; a_mant2 = 8'd170; a_mant3 = 8'd130;
b_mant0 = 8'd0; b_mant1 = 8'd244; b_mant2 = 8'd190; b_mant3 = 8'd156;
a_exp0 = 10'd288; a_exp1 = 10'd405; a_exp2 = 10'd45; a_exp3 = 10'd940;
b_exp0 = 10'd291; b_exp1 = 10'd784; b_exp2 = 10'd636; b_exp3 = 10'd429;
a_sign0 = 4'd11; a_sign1 = 4'd10; a_sign2 = 4'd14; a_sign3 = 4'd7;
b_sign0 = 4'd10; b_sign1 = 4'd11; b_sign2 = 4'd16; b_sign3 = 4'd11;
@(posedge clk_i);
a_mant0 = 8'd29; a_mant1 = 8'd95; a_mant2 = 8'd135; a_mant3 = 8'd254;
b_mant0 = 8'd3; b_mant1 = 8'd242; b_mant2 = 8'd32; b_mant3 = 8'd211;
a_exp0 = 10'd273; a_exp1 = 10'd594; a_exp2 = 10'd704; a_exp3 = 10'd671;
b_exp0 = 10'd395; b_exp1 = 10'd426; b_exp2 = 10'd268; b_exp3 = 10'd191;
a_sign0 = 4'd7; a_sign1 = 4'd3; a_sign2 = 4'd11; a_sign3 = 4'd13;
b_sign0 = 4'd7; b_sign1 = 4'd2; b_sign2 = 4'd14; b_sign3 = 4'd5;
@(posedge clk_i);
a_mant0 = 8'd209; a_mant1 = 8'd66; a_mant2 = 8'd212; a_mant3 = 8'd171;
b_mant0 = 8'd253; b_mant1 = 8'd237; b_mant2 = 8'd127; b_mant3 = 8'd51;
a_exp0 = 10'd776; a_exp1 = 10'd862; a_exp2 = 10'd956; a_exp3 = 10'd79;
b_exp0 = 10'd967; b_exp1 = 10'd741; b_exp2 = 10'd69; b_exp3 = 10'd271;
a_sign0 = 4'd1; a_sign1 = 4'd15; a_sign2 = 4'd7; a_sign3 = 4'd5;
b_sign0 = 4'd6; b_sign1 = 4'd8; b_sign2 = 4'd2; b_sign3 = 4'd9;
@(posedge clk_i);
a_mant0 = 8'd31; a_mant1 = 8'd200; a_mant2 = 8'd160; a_mant3 = 8'd173;
b_mant0 = 8'd136; b_mant1 = 8'd55; b_mant2 = 8'd65; b_mant3 = 8'd71;
a_exp0 = 10'd481; a_exp1 = 10'd80; a_exp2 = 10'd483; a_exp3 = 10'd60;
b_exp0 = 10'd832; b_exp1 = 10'd529; b_exp2 = 10'd578; b_exp3 = 10'd241;
a_sign0 = 4'd13; a_sign1 = 4'd0; a_sign2 = 4'd8; a_sign3 = 4'd9;
b_sign0 = 4'd2; b_sign1 = 4'd3; b_sign2 = 4'd7; b_sign3 = 4'd3;
@(posedge clk_i);
a_mant0 = 8'd116; a_mant1 = 8'd122; a_mant2 = 8'd38; a_mant3 = 8'd231;
b_mant0 = 8'd20; b_mant1 = 8'd15; b_mant2 = 8'd77; b_mant3 = 8'd83;
a_exp0 = 10'd342; a_exp1 = 10'd749; a_exp2 = 10'd533; a_exp3 = 10'd774;
b_exp0 = 10'd705; b_exp1 = 10'd923; b_exp2 = 10'd112; b_exp3 = 10'd119;
a_sign0 = 4'd16; a_sign1 = 4'd8; a_sign2 = 4'd6; a_sign3 = 4'd4;
b_sign0 = 4'd3; b_sign1 = 4'd8; b_sign2 = 4'd11; b_sign3 = 4'd8;
@(posedge clk_i);
shared_exps0 = 8'd135;
shared_exps1 = 8'd102;
a_mant0 = 8'd59; a_mant1 = 8'd77; a_mant2 = 8'd10; a_mant3 = 8'd14;
b_mant0 = 8'd170; b_mant1 = 8'd72; b_mant2 = 8'd26; b_mant3 = 8'd182;
a_exp0 = 10'd546; a_exp1 = 10'd353; a_exp2 = 10'd810; a_exp3 = 10'd944;
b_exp0 = 10'd277; b_exp1 = 10'd713; b_exp2 = 10'd468; b_exp3 = 10'd331;
a_sign0 = 4'd10; a_sign1 = 4'd10; a_sign2 = 4'd14; a_sign3 = 4'd4;
b_sign0 = 4'd1; b_sign1 = 4'd8; b_sign2 = 4'd12; b_sign3 = 4'd12;
@(posedge clk_i);
a_mant0 = 8'd52; a_mant1 = 8'd203; a_mant2 = 8'd154; a_mant3 = 8'd97;
b_mant0 = 8'd56; b_mant1 = 8'd16; b_mant2 = 8'd40; b_mant3 = 8'd119;
a_exp0 = 10'd763; a_exp1 = 10'd184; a_exp2 = 10'd419; a_exp3 = 10'd884;
b_exp0 = 10'd526; b_exp1 = 10'd893; b_exp2 = 10'd655; b_exp3 = 10'd787;
a_sign0 = 4'd2; a_sign1 = 4'd14; a_sign2 = 4'd13; a_sign3 = 4'd13;
b_sign0 = 4'd7; b_sign1 = 4'd14; b_sign2 = 4'd4; b_sign3 = 4'd9;
@(posedge clk_i);
a_mant0 = 8'd150; a_mant1 = 8'd231; a_mant2 = 8'd236; a_mant3 = 8'd172;
b_mant0 = 8'd208; b_mant1 = 8'd213; b_mant2 = 8'd51; b_mant3 = 8'd104;
a_exp0 = 10'd802; a_exp1 = 10'd632; a_exp2 = 10'd216; a_exp3 = 10'd451;
b_exp0 = 10'd457; b_exp1 = 10'd390; b_exp2 = 10'd276; b_exp3 = 10'd187;
a_sign0 = 4'd16; a_sign1 = 4'd12; a_sign2 = 4'd11; a_sign3 = 4'd10;
b_sign0 = 4'd11; b_sign1 = 4'd3; b_sign2 = 4'd1; b_sign3 = 4'd5;
@(posedge clk_i);
a_mant0 = 8'd71; a_mant1 = 8'd222; a_mant2 = 8'd235; a_mant3 = 8'd123;
b_mant0 = 8'd74; b_mant1 = 8'd156; b_mant2 = 8'd207; b_mant3 = 8'd71;
a_exp0 = 10'd388; a_exp1 = 10'd170; a_exp2 = 10'd428; a_exp3 = 10'd813;
b_exp0 = 10'd188; b_exp1 = 10'd183; b_exp2 = 10'd868; b_exp3 = 10'd312;
a_sign0 = 4'd14; a_sign1 = 4'd11; a_sign2 = 4'd2; a_sign3 = 4'd8;
b_sign0 = 4'd15; b_sign1 = 4'd1; b_sign2 = 4'd9; b_sign3 = 4'd10;
@(posedge clk_i);
a_mant0 = 8'd117; a_mant1 = 8'd58; a_mant2 = 8'd20; a_mant3 = 8'd207;
b_mant0 = 8'd79; b_mant1 = 8'd68; b_mant2 = 8'd24; b_mant3 = 8'd174;
a_exp0 = 10'd923; a_exp1 = 10'd161; a_exp2 = 10'd72; a_exp3 = 10'd946;
b_exp0 = 10'd329; b_exp1 = 10'd5; b_exp2 = 10'd285; b_exp3 = 10'd101;
a_sign0 = 4'd14; a_sign1 = 4'd5; a_sign2 = 4'd2; a_sign3 = 4'd4;
b_sign0 = 4'd8; b_sign1 = 4'd10; b_sign2 = 4'd8; b_sign3 = 4'd15;
@(posedge clk_i);
a_mant0 = 8'd142; a_mant1 = 8'd22; a_mant2 = 8'd94; a_mant3 = 8'd110;
b_mant0 = 8'd252; b_mant1 = 8'd61; b_mant2 = 8'd78; b_mant3 = 8'd60;
a_exp0 = 10'd452; a_exp1 = 10'd948; a_exp2 = 10'd592; a_exp3 = 10'd918;
b_exp0 = 10'd820; b_exp1 = 10'd770; b_exp2 = 10'd376; b_exp3 = 10'd141;
a_sign0 = 4'd15; a_sign1 = 4'd12; a_sign2 = 4'd2; a_sign3 = 4'd0;
b_sign0 = 4'd8; b_sign1 = 4'd14; b_sign2 = 4'd11; b_sign3 = 4'd4;
@(posedge clk_i);
a_mant0 = 8'd237; a_mant1 = 8'd132; a_mant2 = 8'd165; a_mant3 = 8'd59;
b_mant0 = 8'd72; b_mant1 = 8'd199; b_mant2 = 8'd24; b_mant3 = 8'd200;
a_exp0 = 10'd675; a_exp1 = 10'd238; a_exp2 = 10'd358; a_exp3 = 10'd114;
b_exp0 = 10'd283; b_exp1 = 10'd492; b_exp2 = 10'd335; b_exp3 = 10'd816;
a_sign0 = 4'd5; a_sign1 = 4'd13; a_sign2 = 4'd12; a_sign3 = 4'd1;
b_sign0 = 4'd5; b_sign1 = 4'd8; b_sign2 = 4'd0; b_sign3 = 4'd14;
@(posedge clk_i);
a_mant0 = 8'd16; a_mant1 = 8'd219; a_mant2 = 8'd47; a_mant3 = 8'd163;
b_mant0 = 8'd241; b_mant1 = 8'd53; b_mant2 = 8'd171; b_mant3 = 8'd195;
a_exp0 = 10'd968; a_exp1 = 10'd540; a_exp2 = 10'd281; a_exp3 = 10'd304;
b_exp0 = 10'd589; b_exp1 = 10'd275; b_exp2 = 10'd214; b_exp3 = 10'd667;
a_sign0 = 4'd9; a_sign1 = 4'd8; a_sign2 = 4'd0; a_sign3 = 4'd14;
b_sign0 = 4'd11; b_sign1 = 4'd6; b_sign2 = 4'd3; b_sign3 = 4'd1;
@(posedge clk_i);
shared_exps0 = 8'd131;
shared_exps1 = 8'd129;
a_mant0 = 8'd219; a_mant1 = 8'd177; a_mant2 = 8'd246; a_mant3 = 8'd147;
b_mant0 = 8'd160; b_mant1 = 8'd236; b_mant2 = 8'd233; b_mant3 = 8'd201;
a_exp0 = 10'd285; a_exp1 = 10'd91; a_exp2 = 10'd792; a_exp3 = 10'd6;
b_exp0 = 10'd797; b_exp1 = 10'd155; b_exp2 = 10'd414; b_exp3 = 10'd180;
a_sign0 = 4'd8; a_sign1 = 4'd0; a_sign2 = 4'd12; a_sign3 = 4'd8;
b_sign0 = 4'd14; b_sign1 = 4'd6; b_sign2 = 4'd1; b_sign3 = 4'd8;
@(posedge clk_i);
a_mant0 = 8'd14; a_mant1 = 8'd246; a_mant2 = 8'd18; a_mant3 = 8'd192;
b_mant0 = 8'd16; b_mant1 = 8'd164; b_mant2 = 8'd151; b_mant3 = 8'd198;
a_exp0 = 10'd824; a_exp1 = 10'd903; a_exp2 = 10'd342; a_exp3 = 10'd182;
b_exp0 = 10'd162; b_exp1 = 10'd937; b_exp2 = 10'd220; b_exp3 = 10'd388;
a_sign0 = 4'd14; a_sign1 = 4'd3; a_sign2 = 4'd1; a_sign3 = 4'd9;
b_sign0 = 4'd12; b_sign1 = 4'd2; b_sign2 = 4'd6; b_sign3 = 4'd11;
@(posedge clk_i);
a_mant0 = 8'd61; a_mant1 = 8'd247; a_mant2 = 8'd153; a_mant3 = 8'd19;
b_mant0 = 8'd34; b_mant1 = 8'd142; b_mant2 = 8'd8; b_mant3 = 8'd153;
a_exp0 = 10'd555; a_exp1 = 10'd272; a_exp2 = 10'd180; a_exp3 = 10'd11;
b_exp0 = 10'd408; b_exp1 = 10'd511; b_exp2 = 10'd762; b_exp3 = 10'd589;
a_sign0 = 4'd4; a_sign1 = 4'd11; a_sign2 = 4'd13; a_sign3 = 4'd5;
b_sign0 = 4'd10; b_sign1 = 4'd12; b_sign2 = 4'd7; b_sign3 = 4'd12;
@(posedge clk_i);
a_mant0 = 8'd165; a_mant1 = 8'd215; a_mant2 = 8'd79; a_mant3 = 8'd116;
b_mant0 = 8'd175; b_mant1 = 8'd120; b_mant2 = 8'd206; b_mant3 = 8'd120;
a_exp0 = 10'd966; a_exp1 = 10'd446; a_exp2 = 10'd221; a_exp3 = 10'd10;
b_exp0 = 10'd507; b_exp1 = 10'd559; b_exp2 = 10'd346; b_exp3 = 10'd720;
a_sign0 = 4'd3; a_sign1 = 4'd9; a_sign2 = 4'd9; a_sign3 = 4'd13;
b_sign0 = 4'd7; b_sign1 = 4'd3; b_sign2 = 4'd16; b_sign3 = 4'd12;
@(posedge clk_i);
a_mant0 = 8'd107; a_mant1 = 8'd201; a_mant2 = 8'd0; a_mant3 = 8'd32;
b_mant0 = 8'd55; b_mant1 = 8'd234; b_mant2 = 8'd82; b_mant3 = 8'd92;
a_exp0 = 10'd882; a_exp1 = 10'd868; a_exp2 = 10'd259; a_exp3 = 10'd410;
b_exp0 = 10'd127; b_exp1 = 10'd42; b_exp2 = 10'd663; b_exp3 = 10'd65;
a_sign0 = 4'd13; a_sign1 = 4'd15; a_sign2 = 4'd9; a_sign3 = 4'd4;
b_sign0 = 4'd13; b_sign1 = 4'd3; b_sign2 = 4'd4; b_sign3 = 4'd3;
@(posedge clk_i);
a_mant0 = 8'd197; a_mant1 = 8'd182; a_mant2 = 8'd159; a_mant3 = 8'd45;
b_mant0 = 8'd204; b_mant1 = 8'd108; b_mant2 = 8'd139; b_mant3 = 8'd168;
a_exp0 = 10'd836; a_exp1 = 10'd241; a_exp2 = 10'd789; a_exp3 = 10'd239;
b_exp0 = 10'd124; b_exp1 = 10'd337; b_exp2 = 10'd136; b_exp3 = 10'd12;
a_sign0 = 4'd5; a_sign1 = 4'd12; a_sign2 = 4'd3; a_sign3 = 4'd7;
b_sign0 = 4'd12; b_sign1 = 4'd13; b_sign2 = 4'd4; b_sign3 = 4'd2;
@(posedge clk_i);
a_mant0 = 8'd167; a_mant1 = 8'd146; a_mant2 = 8'd188; a_mant3 = 8'd40;
b_mant0 = 8'd200; b_mant1 = 8'd167; b_mant2 = 8'd18; b_mant3 = 8'd63;
a_exp0 = 10'd952; a_exp1 = 10'd105; a_exp2 = 10'd787; a_exp3 = 10'd697;
b_exp0 = 10'd50; b_exp1 = 10'd767; b_exp2 = 10'd552; b_exp3 = 10'd891;
a_sign0 = 4'd12; a_sign1 = 4'd16; a_sign2 = 4'd15; a_sign3 = 4'd1;
b_sign0 = 4'd0; b_sign1 = 4'd10; b_sign2 = 4'd8; b_sign3 = 4'd3;
@(posedge clk_i);
a_mant0 = 8'd245; a_mant1 = 8'd215; a_mant2 = 8'd213; a_mant3 = 8'd27;
b_mant0 = 8'd193; b_mant1 = 8'd84; b_mant2 = 8'd8; b_mant3 = 8'd174;
a_exp0 = 10'd119; a_exp1 = 10'd270; a_exp2 = 10'd827; a_exp3 = 10'd655;
b_exp0 = 10'd238; b_exp1 = 10'd200; b_exp2 = 10'd536; b_exp3 = 10'd174;
a_sign0 = 4'd5; a_sign1 = 4'd3; a_sign2 = 4'd0; a_sign3 = 4'd7;
b_sign0 = 4'd10; b_sign1 = 4'd12; b_sign2 = 4'd13; b_sign3 = 4'd0;
@(posedge clk_i);
shared_exps0 = 8'd132;
shared_exps1 = 8'd127;
a_mant0 = 8'd250; a_mant1 = 8'd153; a_mant2 = 8'd129; a_mant3 = 8'd163;
b_mant0 = 8'd64; b_mant1 = 8'd18; b_mant2 = 8'd161; b_mant3 = 8'd157;
a_exp0 = 10'd516; a_exp1 = 10'd356; a_exp2 = 10'd278; a_exp3 = 10'd812;
b_exp0 = 10'd301; b_exp1 = 10'd356; b_exp2 = 10'd656; b_exp3 = 10'd834;
a_sign0 = 4'd6; a_sign1 = 4'd9; a_sign2 = 4'd15; a_sign3 = 4'd7;
b_sign0 = 4'd10; b_sign1 = 4'd3; b_sign2 = 4'd4; b_sign3 = 4'd15;
@(posedge clk_i);
a_mant0 = 8'd182; a_mant1 = 8'd166; a_mant2 = 8'd168; a_mant3 = 8'd241;
b_mant0 = 8'd164; b_mant1 = 8'd181; b_mant2 = 8'd76; b_mant3 = 8'd226;
a_exp0 = 10'd324; a_exp1 = 10'd233; a_exp2 = 10'd154; a_exp3 = 10'd434;
b_exp0 = 10'd342; b_exp1 = 10'd465; b_exp2 = 10'd579; b_exp3 = 10'd749;
a_sign0 = 4'd12; a_sign1 = 4'd0; a_sign2 = 4'd6; a_sign3 = 4'd15;
b_sign0 = 4'd10; b_sign1 = 4'd1; b_sign2 = 4'd12; b_sign3 = 4'd2;
@(posedge clk_i);
a_mant0 = 8'd5; a_mant1 = 8'd130; a_mant2 = 8'd120; a_mant3 = 8'd22;
b_mant0 = 8'd150; b_mant1 = 8'd165; b_mant2 = 8'd112; b_mant3 = 8'd142;
a_exp0 = 10'd201; a_exp1 = 10'd56; a_exp2 = 10'd735; a_exp3 = 10'd69;
b_exp0 = 10'd942; b_exp1 = 10'd598; b_exp2 = 10'd138; b_exp3 = 10'd874;
a_sign0 = 4'd4; a_sign1 = 4'd8; a_sign2 = 4'd4; a_sign3 = 4'd5;
b_sign0 = 4'd13; b_sign1 = 4'd16; b_sign2 = 4'd8; b_sign3 = 4'd14;
@(posedge clk_i);
a_mant0 = 8'd205; a_mant1 = 8'd93; a_mant2 = 8'd33; a_mant3 = 8'd192;
b_mant0 = 8'd232; b_mant1 = 8'd195; b_mant2 = 8'd107; b_mant3 = 8'd122;
a_exp0 = 10'd181; a_exp1 = 10'd777; a_exp2 = 10'd872; a_exp3 = 10'd36;
b_exp0 = 10'd549; b_exp1 = 10'd961; b_exp2 = 10'd251; b_exp3 = 10'd558;
a_sign0 = 4'd3; a_sign1 = 4'd6; a_sign2 = 4'd11; a_sign3 = 4'd2;
b_sign0 = 4'd5; b_sign1 = 4'd8; b_sign2 = 4'd2; b_sign3 = 4'd4;
@(posedge clk_i);
a_mant0 = 8'd191; a_mant1 = 8'd251; a_mant2 = 8'd228; a_mant3 = 8'd36;
b_mant0 = 8'd219; b_mant1 = 8'd183; b_mant2 = 8'd151; b_mant3 = 8'd116;
a_exp0 = 10'd504; a_exp1 = 10'd266; a_exp2 = 10'd416; a_exp3 = 10'd889;
b_exp0 = 10'd862; b_exp1 = 10'd997; b_exp2 = 10'd12; b_exp3 = 10'd788;
a_sign0 = 4'd8; a_sign1 = 4'd14; a_sign2 = 4'd2; a_sign3 = 4'd5;
b_sign0 = 4'd4; b_sign1 = 4'd11; b_sign2 = 4'd10; b_sign3 = 4'd16;
@(posedge clk_i);
a_mant0 = 8'd168; a_mant1 = 8'd234; a_mant2 = 8'd120; a_mant3 = 8'd244;
b_mant0 = 8'd47; b_mant1 = 8'd16; b_mant2 = 8'd176; b_mant3 = 8'd157;
a_exp0 = 10'd250; a_exp1 = 10'd245; a_exp2 = 10'd131; a_exp3 = 10'd87;
b_exp0 = 10'd473; b_exp1 = 10'd234; b_exp2 = 10'd947; b_exp3 = 10'd103;
a_sign0 = 4'd11; a_sign1 = 4'd10; a_sign2 = 4'd3; a_sign3 = 4'd5;
b_sign0 = 4'd15; b_sign1 = 4'd7; b_sign2 = 4'd1; b_sign3 = 4'd5;
@(posedge clk_i);
a_mant0 = 8'd20; a_mant1 = 8'd145; a_mant2 = 8'd126; a_mant3 = 8'd121;
b_mant0 = 8'd185; b_mant1 = 8'd176; b_mant2 = 8'd173; b_mant3 = 8'd194;
a_exp0 = 10'd765; a_exp1 = 10'd471; a_exp2 = 10'd448; a_exp3 = 10'd506;
b_exp0 = 10'd995; b_exp1 = 10'd186; b_exp2 = 10'd173; b_exp3 = 10'd888;
a_sign0 = 4'd9; a_sign1 = 4'd0; a_sign2 = 4'd6; a_sign3 = 4'd9;
b_sign0 = 4'd4; b_sign1 = 4'd7; b_sign2 = 4'd7; b_sign3 = 4'd12;
@(posedge clk_i);
a_mant0 = 8'd254; a_mant1 = 8'd18; a_mant2 = 8'd91; a_mant3 = 8'd185;
b_mant0 = 8'd144; b_mant1 = 8'd250; b_mant2 = 8'd228; b_mant3 = 8'd36;
a_exp0 = 10'd708; a_exp1 = 10'd19; a_exp2 = 10'd262; a_exp3 = 10'd964;
b_exp0 = 10'd535; b_exp1 = 10'd163; b_exp2 = 10'd944; b_exp3 = 10'd401;
a_sign0 = 4'd15; a_sign1 = 4'd2; a_sign2 = 4'd2; a_sign3 = 4'd13;
b_sign0 = 4'd1; b_sign1 = 4'd14; b_sign2 = 4'd9; b_sign3 = 4'd16;
@(posedge clk_i);
shared_exps0 = 8'd131;
shared_exps1 = 8'd153;
rstn = 0;
@(posedge clk_i);
rstn = 1;
a_mant0 = 8'd158; a_mant1 = 8'd63; a_mant2 = 8'd17; a_mant3 = 8'd172;
b_mant0 = 8'd61; b_mant1 = 8'd54; b_mant2 = 8'd229; b_mant3 = 8'd212;
a_exp0 = 10'd873; a_exp1 = 10'd474; a_exp2 = 10'd932; a_exp3 = 10'd683;
b_exp0 = 10'd863; b_exp1 = 10'd961; b_exp2 = 10'd457; b_exp3 = 10'd310;
a_sign0 = 4'd6; a_sign1 = 4'd3; a_sign2 = 4'd7; a_sign3 = 4'd2;
b_sign0 = 4'd7; b_sign1 = 4'd7; b_sign2 = 4'd14; b_sign3 = 4'd12;
@(posedge clk_i);
a_mant0 = 8'd15; a_mant1 = 8'd1; a_mant2 = 8'd134; a_mant3 = 8'd76;
b_mant0 = 8'd39; b_mant1 = 8'd204; b_mant2 = 8'd251; b_mant3 = 8'd156;
a_exp0 = 10'd975; a_exp1 = 10'd993; a_exp2 = 10'd949; a_exp3 = 10'd608;
b_exp0 = 10'd488; b_exp1 = 10'd770; b_exp2 = 10'd878; b_exp3 = 10'd480;
a_sign0 = 4'd12; a_sign1 = 4'd6; a_sign2 = 4'd2; a_sign3 = 4'd8;
b_sign0 = 4'd7; b_sign1 = 4'd12; b_sign2 = 4'd15; b_sign3 = 4'd8;
@(posedge clk_i);
a_mant0 = 8'd75; a_mant1 = 8'd254; a_mant2 = 8'd136; a_mant3 = 8'd199;
b_mant0 = 8'd90; b_mant1 = 8'd84; b_mant2 = 8'd130; b_mant3 = 8'd75;
a_exp0 = 10'd769; a_exp1 = 10'd844; a_exp2 = 10'd196; a_exp3 = 10'd102;
b_exp0 = 10'd68; b_exp1 = 10'd996; b_exp2 = 10'd311; b_exp3 = 10'd533;
a_sign0 = 4'd1; a_sign1 = 4'd6; a_sign2 = 4'd5; a_sign3 = 4'd14;
b_sign0 = 4'd3; b_sign1 = 4'd13; b_sign2 = 4'd12; b_sign3 = 4'd13;
@(posedge clk_i);
a_mant0 = 8'd195; a_mant1 = 8'd132; a_mant2 = 8'd103; a_mant3 = 8'd75;
b_mant0 = 8'd173; b_mant1 = 8'd23; b_mant2 = 8'd196; b_mant3 = 8'd234;
a_exp0 = 10'd1022; a_exp1 = 10'd708; a_exp2 = 10'd986; a_exp3 = 10'd405;
b_exp0 = 10'd525; b_exp1 = 10'd804; b_exp2 = 10'd704; b_exp3 = 10'd131;
a_sign0 = 4'd11; a_sign1 = 4'd10; a_sign2 = 4'd16; a_sign3 = 4'd16;
b_sign0 = 4'd5; b_sign1 = 4'd6; b_sign2 = 4'd13; b_sign3 = 4'd10;
@(posedge clk_i);
a_mant0 = 8'd68; a_mant1 = 8'd243; a_mant2 = 8'd35; a_mant3 = 8'd141;
b_mant0 = 8'd19; b_mant1 = 8'd91; b_mant2 = 8'd89; b_mant3 = 8'd179;
a_exp0 = 10'd990; a_exp1 = 10'd116; a_exp2 = 10'd739; a_exp3 = 10'd791;
b_exp0 = 10'd742; b_exp1 = 10'd906; b_exp2 = 10'd988; b_exp3 = 10'd43;
a_sign0 = 4'd16; a_sign1 = 4'd5; a_sign2 = 4'd6; a_sign3 = 4'd8;
b_sign0 = 4'd16; b_sign1 = 4'd2; b_sign2 = 4'd14; b_sign3 = 4'd10;
@(posedge clk_i);
a_mant0 = 8'd255; a_mant1 = 8'd20; a_mant2 = 8'd86; a_mant3 = 8'd202;
b_mant0 = 8'd113; b_mant1 = 8'd234; b_mant2 = 8'd99; b_mant3 = 8'd227;
a_exp0 = 10'd913; a_exp1 = 10'd816; a_exp2 = 10'd762; a_exp3 = 10'd242;
b_exp0 = 10'd982; b_exp1 = 10'd152; b_exp2 = 10'd864; b_exp3 = 10'd400;
a_sign0 = 4'd2; a_sign1 = 4'd8; a_sign2 = 4'd5; a_sign3 = 4'd1;
b_sign0 = 4'd8; b_sign1 = 4'd4; b_sign2 = 4'd6; b_sign3 = 4'd3;
@(posedge clk_i);
a_mant0 = 8'd71; a_mant1 = 8'd26; a_mant2 = 8'd166; a_mant3 = 8'd11;
b_mant0 = 8'd184; b_mant1 = 8'd63; b_mant2 = 8'd53; b_mant3 = 8'd57;
a_exp0 = 10'd272; a_exp1 = 10'd39; a_exp2 = 10'd900; a_exp3 = 10'd477;
b_exp0 = 10'd462; b_exp1 = 10'd127; b_exp2 = 10'd415; b_exp3 = 10'd196;
a_sign0 = 4'd5; a_sign1 = 4'd4; a_sign2 = 4'd15; a_sign3 = 4'd8;
b_sign0 = 4'd16; b_sign1 = 4'd9; b_sign2 = 4'd3; b_sign3 = 4'd4;
@(posedge clk_i);
shared_exps0 = 8'd154;
shared_exps1 = 8'd149;
a_mant0 = 8'd87; a_mant1 = 8'd21; a_mant2 = 8'd107; a_mant3 = 8'd177;
b_mant0 = 8'd102; b_mant1 = 8'd35; b_mant2 = 8'd166; b_mant3 = 8'd11;
a_exp0 = 10'd921; a_exp1 = 10'd109; a_exp2 = 10'd135; a_exp3 = 10'd154;
b_exp0 = 10'd202; b_exp1 = 10'd20; b_exp2 = 10'd686; b_exp3 = 10'd578;
a_sign0 = 4'd6; a_sign1 = 4'd11; a_sign2 = 4'd8; a_sign3 = 4'd15;
b_sign0 = 4'd15; b_sign1 = 4'd12; b_sign2 = 4'd5; b_sign3 = 4'd12;
@(posedge clk_i);
a_mant0 = 8'd23; a_mant1 = 8'd214; a_mant2 = 8'd210; a_mant3 = 8'd48;
b_mant0 = 8'd127; b_mant1 = 8'd225; b_mant2 = 8'd48; b_mant3 = 8'd146;
a_exp0 = 10'd526; a_exp1 = 10'd661; a_exp2 = 10'd20; a_exp3 = 10'd166;
b_exp0 = 10'd850; b_exp1 = 10'd765; b_exp2 = 10'd437; b_exp3 = 10'd684;
a_sign0 = 4'd14; a_sign1 = 4'd10; a_sign2 = 4'd12; a_sign3 = 4'd9;
b_sign0 = 4'd7; b_sign1 = 4'd2; b_sign2 = 4'd6; b_sign3 = 4'd14;
@(posedge clk_i);
a_mant0 = 8'd113; a_mant1 = 8'd123; a_mant2 = 8'd72; a_mant3 = 8'd223;
b_mant0 = 8'd246; b_mant1 = 8'd22; b_mant2 = 8'd60; b_mant3 = 8'd96;
a_exp0 = 10'd474; a_exp1 = 10'd167; a_exp2 = 10'd450; a_exp3 = 10'd57;
b_exp0 = 10'd515; b_exp1 = 10'd892; b_exp2 = 10'd207; b_exp3 = 10'd294;
a_sign0 = 4'd7; a_sign1 = 4'd8; a_sign2 = 4'd5; a_sign3 = 4'd14;
b_sign0 = 4'd10; b_sign1 = 4'd9; b_sign2 = 4'd11; b_sign3 = 4'd9;
@(posedge clk_i);
a_mant0 = 8'd217; a_mant1 = 8'd151; a_mant2 = 8'd204; a_mant3 = 8'd195;
b_mant0 = 8'd9; b_mant1 = 8'd0; b_mant2 = 8'd1; b_mant3 = 8'd255;
a_exp0 = 10'd647; a_exp1 = 10'd306; a_exp2 = 10'd250; a_exp3 = 10'd535;
b_exp0 = 10'd974; b_exp1 = 10'd880; b_exp2 = 10'd834; b_exp3 = 10'd982;
a_sign0 = 4'd8; a_sign1 = 4'd4; a_sign2 = 4'd8; a_sign3 = 4'd14;
b_sign0 = 4'd0; b_sign1 = 4'd2; b_sign2 = 4'd2; b_sign3 = 4'd13;
@(posedge clk_i);
a_mant0 = 8'd208; a_mant1 = 8'd137; a_mant2 = 8'd106; a_mant3 = 8'd22;
b_mant0 = 8'd145; b_mant1 = 8'd34; b_mant2 = 8'd32; b_mant3 = 8'd86;
a_exp0 = 10'd327; a_exp1 = 10'd352; a_exp2 = 10'd44; a_exp3 = 10'd902;
b_exp0 = 10'd278; b_exp1 = 10'd380; b_exp2 = 10'd686; b_exp3 = 10'd605;
a_sign0 = 4'd9; a_sign1 = 4'd1; a_sign2 = 4'd16; a_sign3 = 4'd9;
b_sign0 = 4'd6; b_sign1 = 4'd4; b_sign2 = 4'd4; b_sign3 = 4'd11;
@(posedge clk_i);
a_mant0 = 8'd94; a_mant1 = 8'd72; a_mant2 = 8'd203; a_mant3 = 8'd238;
b_mant0 = 8'd106; b_mant1 = 8'd66; b_mant2 = 8'd178; b_mant3 = 8'd153;
a_exp0 = 10'd877; a_exp1 = 10'd497; a_exp2 = 10'd290; a_exp3 = 10'd264;
b_exp0 = 10'd930; b_exp1 = 10'd694; b_exp2 = 10'd419; b_exp3 = 10'd967;
a_sign0 = 4'd0; a_sign1 = 4'd16; a_sign2 = 4'd15; a_sign3 = 4'd15;
b_sign0 = 4'd14; b_sign1 = 4'd7; b_sign2 = 4'd16; b_sign3 = 4'd8;
@(posedge clk_i);
a_mant0 = 8'd93; a_mant1 = 8'd165; a_mant2 = 8'd180; a_mant3 = 8'd56;
b_mant0 = 8'd5; b_mant1 = 8'd244; b_mant2 = 8'd147; b_mant3 = 8'd75;
a_exp0 = 10'd453; a_exp1 = 10'd439; a_exp2 = 10'd530; a_exp3 = 10'd195;
b_exp0 = 10'd324; b_exp1 = 10'd39; b_exp2 = 10'd827; b_exp3 = 10'd39;
a_sign0 = 4'd16; a_sign1 = 4'd8; a_sign2 = 4'd5; a_sign3 = 4'd0;
b_sign0 = 4'd7; b_sign1 = 4'd0; b_sign2 = 4'd11; b_sign3 = 4'd14;
@(posedge clk_i);
a_mant0 = 8'd171; a_mant1 = 8'd75; a_mant2 = 8'd87; a_mant3 = 8'd85;
b_mant0 = 8'd254; b_mant1 = 8'd134; b_mant2 = 8'd201; b_mant3 = 8'd87;
a_exp0 = 10'd749; a_exp1 = 10'd506; a_exp2 = 10'd943; a_exp3 = 10'd163;
b_exp0 = 10'd752; b_exp1 = 10'd993; b_exp2 = 10'd904; b_exp3 = 10'd820;
a_sign0 = 4'd6; a_sign1 = 4'd8; a_sign2 = 4'd16; a_sign3 = 4'd6;
b_sign0 = 4'd12; b_sign1 = 4'd0; b_sign2 = 4'd14; b_sign3 = 4'd12;
@(posedge clk_i);
shared_exps0 = 8'd125;
shared_exps1 = 8'd134;
a_mant0 = 8'd93; a_mant1 = 8'd249; a_mant2 = 8'd198; a_mant3 = 8'd155;
b_mant0 = 8'd159; b_mant1 = 8'd60; b_mant2 = 8'd97; b_mant3 = 8'd145;
a_exp0 = 10'd983; a_exp1 = 10'd119; a_exp2 = 10'd708; a_exp3 = 10'd68;
b_exp0 = 10'd33; b_exp1 = 10'd228; b_exp2 = 10'd795; b_exp3 = 10'd520;
a_sign0 = 4'd7; a_sign1 = 4'd6; a_sign2 = 4'd11; a_sign3 = 4'd13;
b_sign0 = 4'd0; b_sign1 = 4'd13; b_sign2 = 4'd4; b_sign3 = 4'd15;
@(posedge clk_i);
a_mant0 = 8'd51; a_mant1 = 8'd137; a_mant2 = 8'd248; a_mant3 = 8'd178;
b_mant0 = 8'd28; b_mant1 = 8'd220; b_mant2 = 8'd235; b_mant3 = 8'd221;
a_exp0 = 10'd16; a_exp1 = 10'd7; a_exp2 = 10'd420; a_exp3 = 10'd462;
b_exp0 = 10'd683; b_exp1 = 10'd558; b_exp2 = 10'd878; b_exp3 = 10'd983;
a_sign0 = 4'd15; a_sign1 = 4'd1; a_sign2 = 4'd0; a_sign3 = 4'd0;
b_sign0 = 4'd10; b_sign1 = 4'd12; b_sign2 = 4'd0; b_sign3 = 4'd16;
@(posedge clk_i);
a_mant0 = 8'd118; a_mant1 = 8'd115; a_mant2 = 8'd244; a_mant3 = 8'd63;
b_mant0 = 8'd254; b_mant1 = 8'd55; b_mant2 = 8'd119; b_mant3 = 8'd227;
a_exp0 = 10'd444; a_exp1 = 10'd421; a_exp2 = 10'd64; a_exp3 = 10'd835;
b_exp0 = 10'd777; b_exp1 = 10'd543; b_exp2 = 10'd116; b_exp3 = 10'd197;
a_sign0 = 4'd6; a_sign1 = 4'd1; a_sign2 = 4'd11; a_sign3 = 4'd10;
b_sign0 = 4'd8; b_sign1 = 4'd7; b_sign2 = 4'd4; b_sign3 = 4'd4;
@(posedge clk_i);
a_mant0 = 8'd153; a_mant1 = 8'd19; a_mant2 = 8'd167; a_mant3 = 8'd9;
b_mant0 = 8'd35; b_mant1 = 8'd70; b_mant2 = 8'd91; b_mant3 = 8'd50;
a_exp0 = 10'd678; a_exp1 = 10'd368; a_exp2 = 10'd239; a_exp3 = 10'd916;
b_exp0 = 10'd932; b_exp1 = 10'd812; b_exp2 = 10'd196; b_exp3 = 10'd141;
a_sign0 = 4'd1; a_sign1 = 4'd8; a_sign2 = 4'd16; a_sign3 = 4'd10;
b_sign0 = 4'd5; b_sign1 = 4'd5; b_sign2 = 4'd7; b_sign3 = 4'd5;
@(posedge clk_i);
a_mant0 = 8'd23; a_mant1 = 8'd34; a_mant2 = 8'd37; a_mant3 = 8'd86;
b_mant0 = 8'd15; b_mant1 = 8'd42; b_mant2 = 8'd5; b_mant3 = 8'd80;
a_exp0 = 10'd321; a_exp1 = 10'd662; a_exp2 = 10'd299; a_exp3 = 10'd640;
b_exp0 = 10'd845; b_exp1 = 10'd338; b_exp2 = 10'd30; b_exp3 = 10'd643;
a_sign0 = 4'd10; a_sign1 = 4'd10; a_sign2 = 4'd14; a_sign3 = 4'd9;
b_sign0 = 4'd3; b_sign1 = 4'd4; b_sign2 = 4'd1; b_sign3 = 4'd11;
@(posedge clk_i);
a_mant0 = 8'd90; a_mant1 = 8'd59; a_mant2 = 8'd172; a_mant3 = 8'd170;
b_mant0 = 8'd210; b_mant1 = 8'd99; b_mant2 = 8'd153; b_mant3 = 8'd77;
a_exp0 = 10'd514; a_exp1 = 10'd89; a_exp2 = 10'd311; a_exp3 = 10'd532;
b_exp0 = 10'd500; b_exp1 = 10'd744; b_exp2 = 10'd882; b_exp3 = 10'd191;
a_sign0 = 4'd10; a_sign1 = 4'd3; a_sign2 = 4'd16; a_sign3 = 4'd11;
b_sign0 = 4'd15; b_sign1 = 4'd1; b_sign2 = 4'd7; b_sign3 = 4'd9;
@(posedge clk_i);
a_mant0 = 8'd223; a_mant1 = 8'd238; a_mant2 = 8'd86; a_mant3 = 8'd30;
b_mant0 = 8'd65; b_mant1 = 8'd23; b_mant2 = 8'd119; b_mant3 = 8'd148;
a_exp0 = 10'd723; a_exp1 = 10'd225; a_exp2 = 10'd384; a_exp3 = 10'd897;
b_exp0 = 10'd699; b_exp1 = 10'd298; b_exp2 = 10'd175; b_exp3 = 10'd129;
a_sign0 = 4'd12; a_sign1 = 4'd9; a_sign2 = 4'd13; a_sign3 = 4'd6;
b_sign0 = 4'd11; b_sign1 = 4'd11; b_sign2 = 4'd14; b_sign3 = 4'd12;
@(posedge clk_i);
a_mant0 = 8'd38; a_mant1 = 8'd254; a_mant2 = 8'd21; a_mant3 = 8'd136;
b_mant0 = 8'd181; b_mant1 = 8'd63; b_mant2 = 8'd77; b_mant3 = 8'd38;
a_exp0 = 10'd844; a_exp1 = 10'd167; a_exp2 = 10'd226; a_exp3 = 10'd899;
b_exp0 = 10'd179; b_exp1 = 10'd715; b_exp2 = 10'd777; b_exp3 = 10'd1021;
a_sign0 = 4'd15; a_sign1 = 4'd9; a_sign2 = 4'd4; a_sign3 = 4'd15;
b_sign0 = 4'd16; b_sign1 = 4'd12; b_sign2 = 4'd10; b_sign3 = 4'd5;
@(posedge clk_i);
shared_exps0 = 8'd104;
shared_exps1 = 8'd105;
a_mant0 = 8'd193; a_mant1 = 8'd72; a_mant2 = 8'd44; a_mant3 = 8'd212;
b_mant0 = 8'd66; b_mant1 = 8'd95; b_mant2 = 8'd33; b_mant3 = 8'd120;
a_exp0 = 10'd261; a_exp1 = 10'd679; a_exp2 = 10'd416; a_exp3 = 10'd862;
b_exp0 = 10'd740; b_exp1 = 10'd998; b_exp2 = 10'd1018; b_exp3 = 10'd155;
a_sign0 = 4'd1; a_sign1 = 4'd3; a_sign2 = 4'd2; a_sign3 = 4'd7;
b_sign0 = 4'd6; b_sign1 = 4'd11; b_sign2 = 4'd2; b_sign3 = 4'd1;
@(posedge clk_i);
a_mant0 = 8'd249; a_mant1 = 8'd152; a_mant2 = 8'd161; a_mant3 = 8'd186;
b_mant0 = 8'd167; b_mant1 = 8'd151; b_mant2 = 8'd44; b_mant3 = 8'd214;
a_exp0 = 10'd671; a_exp1 = 10'd764; a_exp2 = 10'd421; a_exp3 = 10'd286;
b_exp0 = 10'd920; b_exp1 = 10'd631; b_exp2 = 10'd203; b_exp3 = 10'd630;
a_sign0 = 4'd10; a_sign1 = 4'd1; a_sign2 = 4'd3; a_sign3 = 4'd3;
b_sign0 = 4'd13; b_sign1 = 4'd13; b_sign2 = 4'd8; b_sign3 = 4'd6;
@(posedge clk_i);
a_mant0 = 8'd94; a_mant1 = 8'd82; a_mant2 = 8'd98; a_mant3 = 8'd116;
b_mant0 = 8'd219; b_mant1 = 8'd242; b_mant2 = 8'd67; b_mant3 = 8'd37;
a_exp0 = 10'd486; a_exp1 = 10'd253; a_exp2 = 10'd523; a_exp3 = 10'd70;
b_exp0 = 10'd750; b_exp1 = 10'd591; b_exp2 = 10'd384; b_exp3 = 10'd160;
a_sign0 = 4'd4; a_sign1 = 4'd7; a_sign2 = 4'd1; a_sign3 = 4'd12;
b_sign0 = 4'd5; b_sign1 = 4'd0; b_sign2 = 4'd16; b_sign3 = 4'd11;
@(posedge clk_i);
a_mant0 = 8'd148; a_mant1 = 8'd156; a_mant2 = 8'd35; a_mant3 = 8'd71;
b_mant0 = 8'd177; b_mant1 = 8'd56; b_mant2 = 8'd143; b_mant3 = 8'd164;
a_exp0 = 10'd843; a_exp1 = 10'd65; a_exp2 = 10'd532; a_exp3 = 10'd498;
b_exp0 = 10'd983; b_exp1 = 10'd160; b_exp2 = 10'd904; b_exp3 = 10'd701;
a_sign0 = 4'd4; a_sign1 = 4'd8; a_sign2 = 4'd12; a_sign3 = 4'd5;
b_sign0 = 4'd9; b_sign1 = 4'd1; b_sign2 = 4'd14; b_sign3 = 4'd6;
@(posedge clk_i);
a_mant0 = 8'd51; a_mant1 = 8'd95; a_mant2 = 8'd253; a_mant3 = 8'd32;
b_mant0 = 8'd96; b_mant1 = 8'd171; b_mant2 = 8'd229; b_mant3 = 8'd105;
a_exp0 = 10'd442; a_exp1 = 10'd611; a_exp2 = 10'd859; a_exp3 = 10'd197;
b_exp0 = 10'd793; b_exp1 = 10'd659; b_exp2 = 10'd1011; b_exp3 = 10'd542;
a_sign0 = 4'd14; a_sign1 = 4'd12; a_sign2 = 4'd10; a_sign3 = 4'd7;
b_sign0 = 4'd11; b_sign1 = 4'd16; b_sign2 = 4'd2; b_sign3 = 4'd6;
@(posedge clk_i);
a_mant0 = 8'd230; a_mant1 = 8'd16; a_mant2 = 8'd201; a_mant3 = 8'd176;
b_mant0 = 8'd184; b_mant1 = 8'd255; b_mant2 = 8'd3; b_mant3 = 8'd209;
a_exp0 = 10'd540; a_exp1 = 10'd788; a_exp2 = 10'd597; a_exp3 = 10'd255;
b_exp0 = 10'd543; b_exp1 = 10'd876; b_exp2 = 10'd886; b_exp3 = 10'd771;
a_sign0 = 4'd4; a_sign1 = 4'd14; a_sign2 = 4'd13; a_sign3 = 4'd15;
b_sign0 = 4'd3; b_sign1 = 4'd9; b_sign2 = 4'd15; b_sign3 = 4'd6;
@(posedge clk_i);
a_mant0 = 8'd240; a_mant1 = 8'd167; a_mant2 = 8'd149; a_mant3 = 8'd171;
b_mant0 = 8'd4; b_mant1 = 8'd13; b_mant2 = 8'd54; b_mant3 = 8'd221;
a_exp0 = 10'd521; a_exp1 = 10'd957; a_exp2 = 10'd570; a_exp3 = 10'd905;
b_exp0 = 10'd117; b_exp1 = 10'd15; b_exp2 = 10'd210; b_exp3 = 10'd900;
a_sign0 = 4'd1; a_sign1 = 4'd7; a_sign2 = 4'd2; a_sign3 = 4'd8;
b_sign0 = 4'd15; b_sign1 = 4'd10; b_sign2 = 4'd16; b_sign3 = 4'd15;
@(posedge clk_i);
a_mant0 = 8'd226; a_mant1 = 8'd114; a_mant2 = 8'd243; a_mant3 = 8'd127;
b_mant0 = 8'd194; b_mant1 = 8'd239; b_mant2 = 8'd89; b_mant3 = 8'd173;
a_exp0 = 10'd377; a_exp1 = 10'd7; a_exp2 = 10'd105; a_exp3 = 10'd604;
b_exp0 = 10'd784; b_exp1 = 10'd948; b_exp2 = 10'd796; b_exp3 = 10'd196;
a_sign0 = 4'd15; a_sign1 = 4'd9; a_sign2 = 4'd7; a_sign3 = 4'd0;
b_sign0 = 4'd0; b_sign1 = 4'd9; b_sign2 = 4'd11; b_sign3 = 4'd7;
@(posedge clk_i);
shared_exps0 = 8'd128;
shared_exps1 = 8'd111;
rstn = 0;
@(posedge clk_i);
rstn = 1;
a_mant0 = 8'd114; a_mant1 = 8'd180; a_mant2 = 8'd152; a_mant3 = 8'd41;
b_mant0 = 8'd106; b_mant1 = 8'd241; b_mant2 = 8'd204; b_mant3 = 8'd88;
a_exp0 = 10'd13; a_exp1 = 10'd214; a_exp2 = 10'd621; a_exp3 = 10'd506;
b_exp0 = 10'd201; b_exp1 = 10'd170; b_exp2 = 10'd493; b_exp3 = 10'd239;
a_sign0 = 4'd11; a_sign1 = 4'd16; a_sign2 = 4'd1; a_sign3 = 4'd15;
b_sign0 = 4'd1; b_sign1 = 4'd8; b_sign2 = 4'd16; b_sign3 = 4'd11;
@(posedge clk_i);
a_mant0 = 8'd172; a_mant1 = 8'd201; a_mant2 = 8'd97; a_mant3 = 8'd104;
b_mant0 = 8'd177; b_mant1 = 8'd213; b_mant2 = 8'd80; b_mant3 = 8'd135;
a_exp0 = 10'd765; a_exp1 = 10'd832; a_exp2 = 10'd313; a_exp3 = 10'd103;
b_exp0 = 10'd690; b_exp1 = 10'd348; b_exp2 = 10'd264; b_exp3 = 10'd44;
a_sign0 = 4'd13; a_sign1 = 4'd14; a_sign2 = 4'd6; a_sign3 = 4'd16;
b_sign0 = 4'd10; b_sign1 = 4'd13; b_sign2 = 4'd1; b_sign3 = 4'd7;
@(posedge clk_i);
a_mant0 = 8'd241; a_mant1 = 8'd242; a_mant2 = 8'd91; a_mant3 = 8'd191;
b_mant0 = 8'd240; b_mant1 = 8'd44; b_mant2 = 8'd46; b_mant3 = 8'd39;
a_exp0 = 10'd883; a_exp1 = 10'd423; a_exp2 = 10'd386; a_exp3 = 10'd787;
b_exp0 = 10'd6; b_exp1 = 10'd753; b_exp2 = 10'd746; b_exp3 = 10'd140;
a_sign0 = 4'd15; a_sign1 = 4'd14; a_sign2 = 4'd14; a_sign3 = 4'd8;
b_sign0 = 4'd12; b_sign1 = 4'd6; b_sign2 = 4'd10; b_sign3 = 4'd0;
@(posedge clk_i);
a_mant0 = 8'd232; a_mant1 = 8'd90; a_mant2 = 8'd151; a_mant3 = 8'd16;
b_mant0 = 8'd143; b_mant1 = 8'd182; b_mant2 = 8'd3; b_mant3 = 8'd153;
a_exp0 = 10'd253; a_exp1 = 10'd174; a_exp2 = 10'd424; a_exp3 = 10'd661;
b_exp0 = 10'd1023; b_exp1 = 10'd636; b_exp2 = 10'd760; b_exp3 = 10'd147;
a_sign0 = 4'd12; a_sign1 = 4'd5; a_sign2 = 4'd14; a_sign3 = 4'd4;
b_sign0 = 4'd14; b_sign1 = 4'd15; b_sign2 = 4'd15; b_sign3 = 4'd14;
@(posedge clk_i);
a_mant0 = 8'd219; a_mant1 = 8'd234; a_mant2 = 8'd108; a_mant3 = 8'd191;
b_mant0 = 8'd71; b_mant1 = 8'd144; b_mant2 = 8'd112; b_mant3 = 8'd86;
a_exp0 = 10'd122; a_exp1 = 10'd9; a_exp2 = 10'd251; a_exp3 = 10'd676;
b_exp0 = 10'd791; b_exp1 = 10'd738; b_exp2 = 10'd495; b_exp3 = 10'd915;
a_sign0 = 4'd6; a_sign1 = 4'd14; a_sign2 = 4'd15; a_sign3 = 4'd10;
b_sign0 = 4'd3; b_sign1 = 4'd15; b_sign2 = 4'd5; b_sign3 = 4'd5;
@(posedge clk_i);
a_mant0 = 8'd169; a_mant1 = 8'd131; a_mant2 = 8'd224; a_mant3 = 8'd138;
b_mant0 = 8'd83; b_mant1 = 8'd189; b_mant2 = 8'd222; b_mant3 = 8'd151;
a_exp0 = 10'd301; a_exp1 = 10'd66; a_exp2 = 10'd959; a_exp3 = 10'd873;
b_exp0 = 10'd549; b_exp1 = 10'd46; b_exp2 = 10'd292; b_exp3 = 10'd568;
a_sign0 = 4'd11; a_sign1 = 4'd16; a_sign2 = 4'd6; a_sign3 = 4'd8;
b_sign0 = 4'd4; b_sign1 = 4'd13; b_sign2 = 4'd8; b_sign3 = 4'd1;
@(posedge clk_i);
a_mant0 = 8'd96; a_mant1 = 8'd101; a_mant2 = 8'd198; a_mant3 = 8'd5;
b_mant0 = 8'd33; b_mant1 = 8'd125; b_mant2 = 8'd11; b_mant3 = 8'd114;
a_exp0 = 10'd980; a_exp1 = 10'd659; a_exp2 = 10'd102; a_exp3 = 10'd592;
b_exp0 = 10'd590; b_exp1 = 10'd156; b_exp2 = 10'd515; b_exp3 = 10'd351;
a_sign0 = 4'd10; a_sign1 = 4'd0; a_sign2 = 4'd2; a_sign3 = 4'd3;
b_sign0 = 4'd3; b_sign1 = 4'd3; b_sign2 = 4'd6; b_sign3 = 4'd15;
@(posedge clk_i);
shared_exps0 = 8'd135;
shared_exps1 = 8'd100;
a_mant0 = 8'd107; a_mant1 = 8'd242; a_mant2 = 8'd96; a_mant3 = 8'd137;
b_mant0 = 8'd117; b_mant1 = 8'd7; b_mant2 = 8'd49; b_mant3 = 8'd167;
a_exp0 = 10'd46; a_exp1 = 10'd1021; a_exp2 = 10'd899; a_exp3 = 10'd631;
b_exp0 = 10'd694; b_exp1 = 10'd66; b_exp2 = 10'd57; b_exp3 = 10'd508;
a_sign0 = 4'd8; a_sign1 = 4'd9; a_sign2 = 4'd0; a_sign3 = 4'd14;
b_sign0 = 4'd14; b_sign1 = 4'd8; b_sign2 = 4'd0; b_sign3 = 4'd7;
@(posedge clk_i);
a_mant0 = 8'd52; a_mant1 = 8'd99; a_mant2 = 8'd147; a_mant3 = 8'd191;
b_mant0 = 8'd191; b_mant1 = 8'd152; b_mant2 = 8'd62; b_mant3 = 8'd126;
a_exp0 = 10'd518; a_exp1 = 10'd675; a_exp2 = 10'd702; a_exp3 = 10'd837;
b_exp0 = 10'd609; b_exp1 = 10'd339; b_exp2 = 10'd154; b_exp3 = 10'd358;
a_sign0 = 4'd9; a_sign1 = 4'd15; a_sign2 = 4'd1; a_sign3 = 4'd12;
b_sign0 = 4'd8; b_sign1 = 4'd3; b_sign2 = 4'd2; b_sign3 = 4'd12;
@(posedge clk_i);
a_mant0 = 8'd137; a_mant1 = 8'd4; a_mant2 = 8'd116; a_mant3 = 8'd210;
b_mant0 = 8'd221; b_mant1 = 8'd251; b_mant2 = 8'd5; b_mant3 = 8'd81;
a_exp0 = 10'd1007; a_exp1 = 10'd143; a_exp2 = 10'd890; a_exp3 = 10'd561;
b_exp0 = 10'd251; b_exp1 = 10'd52; b_exp2 = 10'd559; b_exp3 = 10'd170;
a_sign0 = 4'd6; a_sign1 = 4'd2; a_sign2 = 4'd6; a_sign3 = 4'd6;
b_sign0 = 4'd9; b_sign1 = 4'd5; b_sign2 = 4'd9; b_sign3 = 4'd12;
@(posedge clk_i);
a_mant0 = 8'd17; a_mant1 = 8'd4; a_mant2 = 8'd30; a_mant3 = 8'd181;
b_mant0 = 8'd99; b_mant1 = 8'd202; b_mant2 = 8'd38; b_mant3 = 8'd125;
a_exp0 = 10'd186; a_exp1 = 10'd493; a_exp2 = 10'd627; a_exp3 = 10'd209;
b_exp0 = 10'd754; b_exp1 = 10'd224; b_exp2 = 10'd972; b_exp3 = 10'd943;
a_sign0 = 4'd16; a_sign1 = 4'd15; a_sign2 = 4'd14; a_sign3 = 4'd10;
b_sign0 = 4'd5; b_sign1 = 4'd14; b_sign2 = 4'd0; b_sign3 = 4'd15;
@(posedge clk_i);
a_mant0 = 8'd181; a_mant1 = 8'd131; a_mant2 = 8'd142; a_mant3 = 8'd83;
b_mant0 = 8'd89; b_mant1 = 8'd86; b_mant2 = 8'd161; b_mant3 = 8'd109;
a_exp0 = 10'd50; a_exp1 = 10'd748; a_exp2 = 10'd910; a_exp3 = 10'd712;
b_exp0 = 10'd711; b_exp1 = 10'd907; b_exp2 = 10'd504; b_exp3 = 10'd298;
a_sign0 = 4'd0; a_sign1 = 4'd6; a_sign2 = 4'd6; a_sign3 = 4'd0;
b_sign0 = 4'd4; b_sign1 = 4'd11; b_sign2 = 4'd0; b_sign3 = 4'd16;
@(posedge clk_i);
a_mant0 = 8'd80; a_mant1 = 8'd6; a_mant2 = 8'd24; a_mant3 = 8'd24;
b_mant0 = 8'd85; b_mant1 = 8'd63; b_mant2 = 8'd31; b_mant3 = 8'd197;
a_exp0 = 10'd574; a_exp1 = 10'd631; a_exp2 = 10'd770; a_exp3 = 10'd548;
b_exp0 = 10'd771; b_exp1 = 10'd278; b_exp2 = 10'd666; b_exp3 = 10'd493;
a_sign0 = 4'd16; a_sign1 = 4'd7; a_sign2 = 4'd5; a_sign3 = 4'd10;
b_sign0 = 4'd1; b_sign1 = 4'd12; b_sign2 = 4'd10; b_sign3 = 4'd11;
@(posedge clk_i);
a_mant0 = 8'd161; a_mant1 = 8'd1; a_mant2 = 8'd125; a_mant3 = 8'd99;
b_mant0 = 8'd191; b_mant1 = 8'd76; b_mant2 = 8'd132; b_mant3 = 8'd101;
a_exp0 = 10'd517; a_exp1 = 10'd752; a_exp2 = 10'd845; a_exp3 = 10'd950;
b_exp0 = 10'd1023; b_exp1 = 10'd684; b_exp2 = 10'd840; b_exp3 = 10'd312;
a_sign0 = 4'd2; a_sign1 = 4'd4; a_sign2 = 4'd7; a_sign3 = 4'd13;
b_sign0 = 4'd11; b_sign1 = 4'd8; b_sign2 = 4'd11; b_sign3 = 4'd6;
@(posedge clk_i);
a_mant0 = 8'd100; a_mant1 = 8'd162; a_mant2 = 8'd203; a_mant3 = 8'd244;
b_mant0 = 8'd75; b_mant1 = 8'd186; b_mant2 = 8'd140; b_mant3 = 8'd152;
a_exp0 = 10'd746; a_exp1 = 10'd663; a_exp2 = 10'd118; a_exp3 = 10'd802;
b_exp0 = 10'd344; b_exp1 = 10'd590; b_exp2 = 10'd280; b_exp3 = 10'd600;
a_sign0 = 4'd16; a_sign1 = 4'd5; a_sign2 = 4'd15; a_sign3 = 4'd6;
b_sign0 = 4'd14; b_sign1 = 4'd10; b_sign2 = 4'd6; b_sign3 = 4'd6;
@(posedge clk_i);
shared_exps0 = 8'd129;
shared_exps1 = 8'd102;
a_mant0 = 8'd188; a_mant1 = 8'd222; a_mant2 = 8'd3; a_mant3 = 8'd169;
b_mant0 = 8'd227; b_mant1 = 8'd158; b_mant2 = 8'd204; b_mant3 = 8'd191;
a_exp0 = 10'd172; a_exp1 = 10'd619; a_exp2 = 10'd638; a_exp3 = 10'd191;
b_exp0 = 10'd299; b_exp1 = 10'd191; b_exp2 = 10'd370; b_exp3 = 10'd154;
a_sign0 = 4'd13; a_sign1 = 4'd4; a_sign2 = 4'd14; a_sign3 = 4'd2;
b_sign0 = 4'd7; b_sign1 = 4'd10; b_sign2 = 4'd7; b_sign3 = 4'd5;
@(posedge clk_i);
a_mant0 = 8'd163; a_mant1 = 8'd238; a_mant2 = 8'd135; a_mant3 = 8'd19;
b_mant0 = 8'd247; b_mant1 = 8'd168; b_mant2 = 8'd103; b_mant3 = 8'd124;
a_exp0 = 10'd101; a_exp1 = 10'd614; a_exp2 = 10'd202; a_exp3 = 10'd98;
b_exp0 = 10'd137; b_exp1 = 10'd532; b_exp2 = 10'd405; b_exp3 = 10'd181;
a_sign0 = 4'd3; a_sign1 = 4'd6; a_sign2 = 4'd10; a_sign3 = 4'd15;
b_sign0 = 4'd13; b_sign1 = 4'd16; b_sign2 = 4'd15; b_sign3 = 4'd14;
@(posedge clk_i);
a_mant0 = 8'd12; a_mant1 = 8'd76; a_mant2 = 8'd221; a_mant3 = 8'd80;
b_mant0 = 8'd218; b_mant1 = 8'd99; b_mant2 = 8'd47; b_mant3 = 8'd19;
a_exp0 = 10'd211; a_exp1 = 10'd319; a_exp2 = 10'd836; a_exp3 = 10'd725;
b_exp0 = 10'd500; b_exp1 = 10'd961; b_exp2 = 10'd122; b_exp3 = 10'd847;
a_sign0 = 4'd5; a_sign1 = 4'd3; a_sign2 = 4'd5; a_sign3 = 4'd15;
b_sign0 = 4'd11; b_sign1 = 4'd9; b_sign2 = 4'd1; b_sign3 = 4'd5;
@(posedge clk_i);
a_mant0 = 8'd229; a_mant1 = 8'd99; a_mant2 = 8'd29; a_mant3 = 8'd200;
b_mant0 = 8'd21; b_mant1 = 8'd107; b_mant2 = 8'd75; b_mant3 = 8'd159;
a_exp0 = 10'd622; a_exp1 = 10'd463; a_exp2 = 10'd574; a_exp3 = 10'd723;
b_exp0 = 10'd625; b_exp1 = 10'd1021; b_exp2 = 10'd59; b_exp3 = 10'd428;
a_sign0 = 4'd4; a_sign1 = 4'd15; a_sign2 = 4'd0; a_sign3 = 4'd1;
b_sign0 = 4'd9; b_sign1 = 4'd11; b_sign2 = 4'd4; b_sign3 = 4'd7;
@(posedge clk_i);
a_mant0 = 8'd145; a_mant1 = 8'd128; a_mant2 = 8'd133; a_mant3 = 8'd50;
b_mant0 = 8'd102; b_mant1 = 8'd39; b_mant2 = 8'd33; b_mant3 = 8'd0;
a_exp0 = 10'd839; a_exp1 = 10'd270; a_exp2 = 10'd361; a_exp3 = 10'd108;
b_exp0 = 10'd776; b_exp1 = 10'd181; b_exp2 = 10'd1005; b_exp3 = 10'd57;
a_sign0 = 4'd6; a_sign1 = 4'd7; a_sign2 = 4'd10; a_sign3 = 4'd5;
b_sign0 = 4'd9; b_sign1 = 4'd0; b_sign2 = 4'd16; b_sign3 = 4'd1;
@(posedge clk_i);
a_mant0 = 8'd160; a_mant1 = 8'd126; a_mant2 = 8'd146; a_mant3 = 8'd21;
b_mant0 = 8'd157; b_mant1 = 8'd136; b_mant2 = 8'd243; b_mant3 = 8'd110;
a_exp0 = 10'd887; a_exp1 = 10'd122; a_exp2 = 10'd767; a_exp3 = 10'd846;
b_exp0 = 10'd104; b_exp1 = 10'd827; b_exp2 = 10'd109; b_exp3 = 10'd524;
a_sign0 = 4'd15; a_sign1 = 4'd4; a_sign2 = 4'd11; a_sign3 = 4'd2;
b_sign0 = 4'd13; b_sign1 = 4'd3; b_sign2 = 4'd2; b_sign3 = 4'd7;
@(posedge clk_i);
a_mant0 = 8'd57; a_mant1 = 8'd92; a_mant2 = 8'd146; a_mant3 = 8'd192;
b_mant0 = 8'd6; b_mant1 = 8'd155; b_mant2 = 8'd11; b_mant3 = 8'd18;
a_exp0 = 10'd74; a_exp1 = 10'd988; a_exp2 = 10'd10; a_exp3 = 10'd361;
b_exp0 = 10'd703; b_exp1 = 10'd671; b_exp2 = 10'd292; b_exp3 = 10'd966;
a_sign0 = 4'd8; a_sign1 = 4'd6; a_sign2 = 4'd12; a_sign3 = 4'd2;
b_sign0 = 4'd5; b_sign1 = 4'd9; b_sign2 = 4'd16; b_sign3 = 4'd16;
@(posedge clk_i);
a_mant0 = 8'd7; a_mant1 = 8'd211; a_mant2 = 8'd24; a_mant3 = 8'd83;
b_mant0 = 8'd0; b_mant1 = 8'd114; b_mant2 = 8'd93; b_mant3 = 8'd48;
a_exp0 = 10'd844; a_exp1 = 10'd861; a_exp2 = 10'd568; a_exp3 = 10'd939;
b_exp0 = 10'd577; b_exp1 = 10'd837; b_exp2 = 10'd356; b_exp3 = 10'd939;
a_sign0 = 4'd6; a_sign1 = 4'd4; a_sign2 = 4'd14; a_sign3 = 4'd13;
b_sign0 = 4'd5; b_sign1 = 4'd5; b_sign2 = 4'd2; b_sign3 = 4'd1;
@(posedge clk_i);
shared_exps0 = 8'd144;
shared_exps1 = 8'd103;
a_mant0 = 8'd60; a_mant1 = 8'd62; a_mant2 = 8'd31; a_mant3 = 8'd87;
b_mant0 = 8'd99; b_mant1 = 8'd89; b_mant2 = 8'd190; b_mant3 = 8'd1;
a_exp0 = 10'd602; a_exp1 = 10'd677; a_exp2 = 10'd982; a_exp3 = 10'd143;
b_exp0 = 10'd651; b_exp1 = 10'd420; b_exp2 = 10'd578; b_exp3 = 10'd1008;
a_sign0 = 4'd8; a_sign1 = 4'd4; a_sign2 = 4'd6; a_sign3 = 4'd0;
b_sign0 = 4'd11; b_sign1 = 4'd11; b_sign2 = 4'd12; b_sign3 = 4'd8;
@(posedge clk_i);
a_mant0 = 8'd120; a_mant1 = 8'd247; a_mant2 = 8'd210; a_mant3 = 8'd238;
b_mant0 = 8'd109; b_mant1 = 8'd87; b_mant2 = 8'd167; b_mant3 = 8'd230;
a_exp0 = 10'd415; a_exp1 = 10'd588; a_exp2 = 10'd923; a_exp3 = 10'd365;
b_exp0 = 10'd219; b_exp1 = 10'd629; b_exp2 = 10'd833; b_exp3 = 10'd878;
a_sign0 = 4'd0; a_sign1 = 4'd1; a_sign2 = 4'd15; a_sign3 = 4'd6;
b_sign0 = 4'd10; b_sign1 = 4'd11; b_sign2 = 4'd7; b_sign3 = 4'd6;
@(posedge clk_i);
a_mant0 = 8'd151; a_mant1 = 8'd102; a_mant2 = 8'd181; a_mant3 = 8'd70;
b_mant0 = 8'd56; b_mant1 = 8'd200; b_mant2 = 8'd222; b_mant3 = 8'd110;
a_exp0 = 10'd185; a_exp1 = 10'd1011; a_exp2 = 10'd444; a_exp3 = 10'd986;
b_exp0 = 10'd525; b_exp1 = 10'd974; b_exp2 = 10'd678; b_exp3 = 10'd974;
a_sign0 = 4'd16; a_sign1 = 4'd4; a_sign2 = 4'd8; a_sign3 = 4'd0;
b_sign0 = 4'd12; b_sign1 = 4'd16; b_sign2 = 4'd7; b_sign3 = 4'd8;
@(posedge clk_i);
a_mant0 = 8'd132; a_mant1 = 8'd113; a_mant2 = 8'd235; a_mant3 = 8'd157;
b_mant0 = 8'd81; b_mant1 = 8'd186; b_mant2 = 8'd38; b_mant3 = 8'd103;
a_exp0 = 10'd626; a_exp1 = 10'd122; a_exp2 = 10'd26; a_exp3 = 10'd385;
b_exp0 = 10'd669; b_exp1 = 10'd237; b_exp2 = 10'd696; b_exp3 = 10'd946;
a_sign0 = 4'd13; a_sign1 = 4'd9; a_sign2 = 4'd16; a_sign3 = 4'd8;
b_sign0 = 4'd0; b_sign1 = 4'd9; b_sign2 = 4'd10; b_sign3 = 4'd10;
@(posedge clk_i);
a_mant0 = 8'd28; a_mant1 = 8'd246; a_mant2 = 8'd220; a_mant3 = 8'd92;
b_mant0 = 8'd1; b_mant1 = 8'd86; b_mant2 = 8'd232; b_mant3 = 8'd81;
a_exp0 = 10'd816; a_exp1 = 10'd861; a_exp2 = 10'd357; a_exp3 = 10'd959;
b_exp0 = 10'd421; b_exp1 = 10'd769; b_exp2 = 10'd319; b_exp3 = 10'd180;
a_sign0 = 4'd2; a_sign1 = 4'd12; a_sign2 = 4'd10; a_sign3 = 4'd1;
b_sign0 = 4'd0; b_sign1 = 4'd11; b_sign2 = 4'd8; b_sign3 = 4'd5;
@(posedge clk_i);
a_mant0 = 8'd152; a_mant1 = 8'd96; a_mant2 = 8'd44; a_mant3 = 8'd13;
b_mant0 = 8'd225; b_mant1 = 8'd22; b_mant2 = 8'd92; b_mant3 = 8'd164;
a_exp0 = 10'd756; a_exp1 = 10'd258; a_exp2 = 10'd654; a_exp3 = 10'd245;
b_exp0 = 10'd163; b_exp1 = 10'd524; b_exp2 = 10'd836; b_exp3 = 10'd746;
a_sign0 = 4'd6; a_sign1 = 4'd10; a_sign2 = 4'd16; a_sign3 = 4'd1;
b_sign0 = 4'd5; b_sign1 = 4'd2; b_sign2 = 4'd13; b_sign3 = 4'd10;
@(posedge clk_i);
a_mant0 = 8'd133; a_mant1 = 8'd95; a_mant2 = 8'd44; a_mant3 = 8'd18;
b_mant0 = 8'd89; b_mant1 = 8'd161; b_mant2 = 8'd219; b_mant3 = 8'd219;
a_exp0 = 10'd812; a_exp1 = 10'd441; a_exp2 = 10'd97; a_exp3 = 10'd489;
b_exp0 = 10'd979; b_exp1 = 10'd783; b_exp2 = 10'd995; b_exp3 = 10'd176;
a_sign0 = 4'd12; a_sign1 = 4'd14; a_sign2 = 4'd5; a_sign3 = 4'd14;
b_sign0 = 4'd12; b_sign1 = 4'd4; b_sign2 = 4'd7; b_sign3 = 4'd11;
@(posedge clk_i);
a_mant0 = 8'd16; a_mant1 = 8'd87; a_mant2 = 8'd228; a_mant3 = 8'd182;
b_mant0 = 8'd223; b_mant1 = 8'd95; b_mant2 = 8'd149; b_mant3 = 8'd101;
a_exp0 = 10'd569; a_exp1 = 10'd629; a_exp2 = 10'd56; a_exp3 = 10'd316;
b_exp0 = 10'd159; b_exp1 = 10'd269; b_exp2 = 10'd522; b_exp3 = 10'd723;
a_sign0 = 4'd10; a_sign1 = 4'd7; a_sign2 = 4'd16; a_sign3 = 4'd5;
b_sign0 = 4'd2; b_sign1 = 4'd9; b_sign2 = 4'd3; b_sign3 = 4'd14;
@(posedge clk_i);
shared_exps0 = 8'd114;
shared_exps1 = 8'd150;
rstn = 0;
@(posedge clk_i);
rstn = 1;
a_mant0 = 8'd53; a_mant1 = 8'd73; a_mant2 = 8'd228; a_mant3 = 8'd15;
b_mant0 = 8'd224; b_mant1 = 8'd81; b_mant2 = 8'd126; b_mant3 = 8'd28;
a_exp0 = 10'd625; a_exp1 = 10'd552; a_exp2 = 10'd995; a_exp3 = 10'd509;
b_exp0 = 10'd342; b_exp1 = 10'd710; b_exp2 = 10'd136; b_exp3 = 10'd484;
a_sign0 = 4'd3; a_sign1 = 4'd4; a_sign2 = 4'd15; a_sign3 = 4'd16;
b_sign0 = 4'd7; b_sign1 = 4'd0; b_sign2 = 4'd14; b_sign3 = 4'd7;
@(posedge clk_i);
a_mant0 = 8'd132; a_mant1 = 8'd153; a_mant2 = 8'd35; a_mant3 = 8'd82;
b_mant0 = 8'd13; b_mant1 = 8'd222; b_mant2 = 8'd158; b_mant3 = 8'd20;
a_exp0 = 10'd325; a_exp1 = 10'd302; a_exp2 = 10'd635; a_exp3 = 10'd857;
b_exp0 = 10'd957; b_exp1 = 10'd38; b_exp2 = 10'd633; b_exp3 = 10'd62;
a_sign0 = 4'd16; a_sign1 = 4'd10; a_sign2 = 4'd12; a_sign3 = 4'd0;
b_sign0 = 4'd16; b_sign1 = 4'd2; b_sign2 = 4'd2; b_sign3 = 4'd5;
@(posedge clk_i);
a_mant0 = 8'd189; a_mant1 = 8'd132; a_mant2 = 8'd229; a_mant3 = 8'd185;
b_mant0 = 8'd47; b_mant1 = 8'd56; b_mant2 = 8'd124; b_mant3 = 8'd177;
a_exp0 = 10'd843; a_exp1 = 10'd638; a_exp2 = 10'd1020; a_exp3 = 10'd963;
b_exp0 = 10'd445; b_exp1 = 10'd715; b_exp2 = 10'd575; b_exp3 = 10'd129;
a_sign0 = 4'd3; a_sign1 = 4'd14; a_sign2 = 4'd7; a_sign3 = 4'd8;
b_sign0 = 4'd6; b_sign1 = 4'd9; b_sign2 = 4'd12; b_sign3 = 4'd10;
@(posedge clk_i);
a_mant0 = 8'd39; a_mant1 = 8'd182; a_mant2 = 8'd126; a_mant3 = 8'd1;
b_mant0 = 8'd125; b_mant1 = 8'd164; b_mant2 = 8'd205; b_mant3 = 8'd147;
a_exp0 = 10'd13; a_exp1 = 10'd658; a_exp2 = 10'd933; a_exp3 = 10'd588;
b_exp0 = 10'd743; b_exp1 = 10'd241; b_exp2 = 10'd123; b_exp3 = 10'd543;
a_sign0 = 4'd9; a_sign1 = 4'd2; a_sign2 = 4'd10; a_sign3 = 4'd3;
b_sign0 = 4'd12; b_sign1 = 4'd10; b_sign2 = 4'd15; b_sign3 = 4'd12;
@(posedge clk_i);
a_mant0 = 8'd60; a_mant1 = 8'd165; a_mant2 = 8'd242; a_mant3 = 8'd128;
b_mant0 = 8'd88; b_mant1 = 8'd251; b_mant2 = 8'd238; b_mant3 = 8'd64;
a_exp0 = 10'd355; a_exp1 = 10'd695; a_exp2 = 10'd540; a_exp3 = 10'd613;
b_exp0 = 10'd273; b_exp1 = 10'd627; b_exp2 = 10'd388; b_exp3 = 10'd209;
a_sign0 = 4'd15; a_sign1 = 4'd16; a_sign2 = 4'd5; a_sign3 = 4'd12;
b_sign0 = 4'd16; b_sign1 = 4'd11; b_sign2 = 4'd14; b_sign3 = 4'd3;
@(posedge clk_i);
a_mant0 = 8'd8; a_mant1 = 8'd121; a_mant2 = 8'd253; a_mant3 = 8'd165;
b_mant0 = 8'd244; b_mant1 = 8'd116; b_mant2 = 8'd233; b_mant3 = 8'd168;
a_exp0 = 10'd759; a_exp1 = 10'd677; a_exp2 = 10'd815; a_exp3 = 10'd501;
b_exp0 = 10'd854; b_exp1 = 10'd493; b_exp2 = 10'd556; b_exp3 = 10'd638;
a_sign0 = 4'd10; a_sign1 = 4'd12; a_sign2 = 4'd15; a_sign3 = 4'd14;
b_sign0 = 4'd16; b_sign1 = 4'd6; b_sign2 = 4'd16; b_sign3 = 4'd9;
@(posedge clk_i);
a_mant0 = 8'd201; a_mant1 = 8'd212; a_mant2 = 8'd99; a_mant3 = 8'd61;
b_mant0 = 8'd85; b_mant1 = 8'd57; b_mant2 = 8'd110; b_mant3 = 8'd0;
a_exp0 = 10'd711; a_exp1 = 10'd752; a_exp2 = 10'd109; a_exp3 = 10'd118;
b_exp0 = 10'd82; b_exp1 = 10'd759; b_exp2 = 10'd231; b_exp3 = 10'd962;
a_sign0 = 4'd0; a_sign1 = 4'd10; a_sign2 = 4'd10; a_sign3 = 4'd7;
b_sign0 = 4'd10; b_sign1 = 4'd4; b_sign2 = 4'd5; b_sign3 = 4'd6;
@(posedge clk_i);
shared_exps0 = 8'd117;
shared_exps1 = 8'd101;
a_mant0 = 8'd115; a_mant1 = 8'd66; a_mant2 = 8'd80; a_mant3 = 8'd133;
b_mant0 = 8'd211; b_mant1 = 8'd93; b_mant2 = 8'd54; b_mant3 = 8'd208;
a_exp0 = 10'd172; a_exp1 = 10'd893; a_exp2 = 10'd694; a_exp3 = 10'd32;
b_exp0 = 10'd287; b_exp1 = 10'd737; b_exp2 = 10'd279; b_exp3 = 10'd501;
a_sign0 = 4'd14; a_sign1 = 4'd12; a_sign2 = 4'd2; a_sign3 = 4'd6;
b_sign0 = 4'd6; b_sign1 = 4'd7; b_sign2 = 4'd8; b_sign3 = 4'd11;
@(posedge clk_i);
a_mant0 = 8'd236; a_mant1 = 8'd28; a_mant2 = 8'd237; a_mant3 = 8'd26;
b_mant0 = 8'd18; b_mant1 = 8'd30; b_mant2 = 8'd91; b_mant3 = 8'd8;
a_exp0 = 10'd347; a_exp1 = 10'd376; a_exp2 = 10'd1017; a_exp3 = 10'd68;
b_exp0 = 10'd302; b_exp1 = 10'd920; b_exp2 = 10'd411; b_exp3 = 10'd895;
a_sign0 = 4'd16; a_sign1 = 4'd8; a_sign2 = 4'd6; a_sign3 = 4'd15;
b_sign0 = 4'd1; b_sign1 = 4'd10; b_sign2 = 4'd15; b_sign3 = 4'd8;
@(posedge clk_i);
a_mant0 = 8'd44; a_mant1 = 8'd193; a_mant2 = 8'd54; a_mant3 = 8'd97;
b_mant0 = 8'd206; b_mant1 = 8'd101; b_mant2 = 8'd168; b_mant3 = 8'd159;
a_exp0 = 10'd122; a_exp1 = 10'd782; a_exp2 = 10'd435; a_exp3 = 10'd991;
b_exp0 = 10'd291; b_exp1 = 10'd998; b_exp2 = 10'd693; b_exp3 = 10'd378;
a_sign0 = 4'd10; a_sign1 = 4'd7; a_sign2 = 4'd14; a_sign3 = 4'd5;
b_sign0 = 4'd10; b_sign1 = 4'd6; b_sign2 = 4'd0; b_sign3 = 4'd11;
@(posedge clk_i);
a_mant0 = 8'd47; a_mant1 = 8'd19; a_mant2 = 8'd84; a_mant3 = 8'd215;
b_mant0 = 8'd129; b_mant1 = 8'd123; b_mant2 = 8'd239; b_mant3 = 8'd0;
a_exp0 = 10'd315; a_exp1 = 10'd409; a_exp2 = 10'd752; a_exp3 = 10'd634;
b_exp0 = 10'd538; b_exp1 = 10'd711; b_exp2 = 10'd234; b_exp3 = 10'd792;
a_sign0 = 4'd6; a_sign1 = 4'd7; a_sign2 = 4'd15; a_sign3 = 4'd8;
b_sign0 = 4'd16; b_sign1 = 4'd1; b_sign2 = 4'd16; b_sign3 = 4'd3;
@(posedge clk_i);
a_mant0 = 8'd145; a_mant1 = 8'd173; a_mant2 = 8'd149; a_mant3 = 8'd166;
b_mant0 = 8'd192; b_mant1 = 8'd12; b_mant2 = 8'd159; b_mant3 = 8'd211;
a_exp0 = 10'd969; a_exp1 = 10'd16; a_exp2 = 10'd560; a_exp3 = 10'd235;
b_exp0 = 10'd40; b_exp1 = 10'd1019; b_exp2 = 10'd253; b_exp3 = 10'd325;
a_sign0 = 4'd16; a_sign1 = 4'd3; a_sign2 = 4'd5; a_sign3 = 4'd15;
b_sign0 = 4'd9; b_sign1 = 4'd13; b_sign2 = 4'd0; b_sign3 = 4'd15;
@(posedge clk_i);
a_mant0 = 8'd229; a_mant1 = 8'd37; a_mant2 = 8'd227; a_mant3 = 8'd67;
b_mant0 = 8'd172; b_mant1 = 8'd57; b_mant2 = 8'd199; b_mant3 = 8'd160;
a_exp0 = 10'd311; a_exp1 = 10'd956; a_exp2 = 10'd89; a_exp3 = 10'd810;
b_exp0 = 10'd1016; b_exp1 = 10'd876; b_exp2 = 10'd133; b_exp3 = 10'd980;
a_sign0 = 4'd8; a_sign1 = 4'd1; a_sign2 = 4'd1; a_sign3 = 4'd3;
b_sign0 = 4'd6; b_sign1 = 4'd0; b_sign2 = 4'd15; b_sign3 = 4'd6;
@(posedge clk_i);
a_mant0 = 8'd240; a_mant1 = 8'd221; a_mant2 = 8'd32; a_mant3 = 8'd205;
b_mant0 = 8'd123; b_mant1 = 8'd151; b_mant2 = 8'd233; b_mant3 = 8'd72;
a_exp0 = 10'd377; a_exp1 = 10'd62; a_exp2 = 10'd154; a_exp3 = 10'd749;
b_exp0 = 10'd282; b_exp1 = 10'd415; b_exp2 = 10'd624; b_exp3 = 10'd153;
a_sign0 = 4'd5; a_sign1 = 4'd12; a_sign2 = 4'd7; a_sign3 = 4'd5;
b_sign0 = 4'd12; b_sign1 = 4'd16; b_sign2 = 4'd13; b_sign3 = 4'd12;
@(posedge clk_i);
a_mant0 = 8'd187; a_mant1 = 8'd225; a_mant2 = 8'd69; a_mant3 = 8'd76;
b_mant0 = 8'd155; b_mant1 = 8'd229; b_mant2 = 8'd162; b_mant3 = 8'd20;
a_exp0 = 10'd16; a_exp1 = 10'd792; a_exp2 = 10'd939; a_exp3 = 10'd777;
b_exp0 = 10'd333; b_exp1 = 10'd596; b_exp2 = 10'd130; b_exp3 = 10'd831;
a_sign0 = 4'd6; a_sign1 = 4'd16; a_sign2 = 4'd16; a_sign3 = 4'd2;
b_sign0 = 4'd4; b_sign1 = 4'd7; b_sign2 = 4'd9; b_sign3 = 4'd11;
@(posedge clk_i);
shared_exps0 = 8'd130;
shared_exps1 = 8'd115;
a_mant0 = 8'd30; a_mant1 = 8'd107; a_mant2 = 8'd204; a_mant3 = 8'd148;
b_mant0 = 8'd152; b_mant1 = 8'd103; b_mant2 = 8'd208; b_mant3 = 8'd237;
a_exp0 = 10'd464; a_exp1 = 10'd344; a_exp2 = 10'd844; a_exp3 = 10'd427;
b_exp0 = 10'd684; b_exp1 = 10'd98; b_exp2 = 10'd233; b_exp3 = 10'd348;
a_sign0 = 4'd6; a_sign1 = 4'd5; a_sign2 = 4'd8; a_sign3 = 4'd4;
b_sign0 = 4'd11; b_sign1 = 4'd6; b_sign2 = 4'd6; b_sign3 = 4'd7;
@(posedge clk_i);
a_mant0 = 8'd116; a_mant1 = 8'd134; a_mant2 = 8'd68; a_mant3 = 8'd104;
b_mant0 = 8'd236; b_mant1 = 8'd177; b_mant2 = 8'd16; b_mant3 = 8'd19;
a_exp0 = 10'd623; a_exp1 = 10'd420; a_exp2 = 10'd756; a_exp3 = 10'd51;
b_exp0 = 10'd1011; b_exp1 = 10'd548; b_exp2 = 10'd605; b_exp3 = 10'd1010;
a_sign0 = 4'd14; a_sign1 = 4'd16; a_sign2 = 4'd14; a_sign3 = 4'd15;
b_sign0 = 4'd14; b_sign1 = 4'd11; b_sign2 = 4'd8; b_sign3 = 4'd12;
@(posedge clk_i);
a_mant0 = 8'd137; a_mant1 = 8'd184; a_mant2 = 8'd214; a_mant3 = 8'd250;
b_mant0 = 8'd79; b_mant1 = 8'd168; b_mant2 = 8'd82; b_mant3 = 8'd20;
a_exp0 = 10'd365; a_exp1 = 10'd395; a_exp2 = 10'd13; a_exp3 = 10'd294;
b_exp0 = 10'd56; b_exp1 = 10'd842; b_exp2 = 10'd384; b_exp3 = 10'd12;
a_sign0 = 4'd9; a_sign1 = 4'd1; a_sign2 = 4'd12; a_sign3 = 4'd6;
b_sign0 = 4'd8; b_sign1 = 4'd6; b_sign2 = 4'd7; b_sign3 = 4'd4;
@(posedge clk_i);
a_mant0 = 8'd85; a_mant1 = 8'd240; a_mant2 = 8'd99; a_mant3 = 8'd93;
b_mant0 = 8'd177; b_mant1 = 8'd43; b_mant2 = 8'd76; b_mant3 = 8'd60;
a_exp0 = 10'd856; a_exp1 = 10'd739; a_exp2 = 10'd352; a_exp3 = 10'd695;
b_exp0 = 10'd155; b_exp1 = 10'd591; b_exp2 = 10'd275; b_exp3 = 10'd635;
a_sign0 = 4'd5; a_sign1 = 4'd4; a_sign2 = 4'd3; a_sign3 = 4'd16;
b_sign0 = 4'd12; b_sign1 = 4'd15; b_sign2 = 4'd13; b_sign3 = 4'd9;
@(posedge clk_i);
a_mant0 = 8'd241; a_mant1 = 8'd48; a_mant2 = 8'd36; a_mant3 = 8'd23;
b_mant0 = 8'd87; b_mant1 = 8'd249; b_mant2 = 8'd198; b_mant3 = 8'd166;
a_exp0 = 10'd454; a_exp1 = 10'd288; a_exp2 = 10'd692; a_exp3 = 10'd933;
b_exp0 = 10'd585; b_exp1 = 10'd393; b_exp2 = 10'd1017; b_exp3 = 10'd380;
a_sign0 = 4'd14; a_sign1 = 4'd2; a_sign2 = 4'd9; a_sign3 = 4'd11;
b_sign0 = 4'd16; b_sign1 = 4'd11; b_sign2 = 4'd8; b_sign3 = 4'd6;
@(posedge clk_i);
a_mant0 = 8'd180; a_mant1 = 8'd134; a_mant2 = 8'd20; a_mant3 = 8'd119;
b_mant0 = 8'd185; b_mant1 = 8'd61; b_mant2 = 8'd210; b_mant3 = 8'd164;
a_exp0 = 10'd42; a_exp1 = 10'd577; a_exp2 = 10'd419; a_exp3 = 10'd757;
b_exp0 = 10'd237; b_exp1 = 10'd203; b_exp2 = 10'd86; b_exp3 = 10'd106;
a_sign0 = 4'd10; a_sign1 = 4'd13; a_sign2 = 4'd9; a_sign3 = 4'd0;
b_sign0 = 4'd9; b_sign1 = 4'd1; b_sign2 = 4'd9; b_sign3 = 4'd9;
@(posedge clk_i);
a_mant0 = 8'd30; a_mant1 = 8'd151; a_mant2 = 8'd132; a_mant3 = 8'd236;
b_mant0 = 8'd50; b_mant1 = 8'd128; b_mant2 = 8'd201; b_mant3 = 8'd82;
a_exp0 = 10'd113; a_exp1 = 10'd357; a_exp2 = 10'd540; a_exp3 = 10'd981;
b_exp0 = 10'd461; b_exp1 = 10'd677; b_exp2 = 10'd804; b_exp3 = 10'd131;
a_sign0 = 4'd14; a_sign1 = 4'd1; a_sign2 = 4'd14; a_sign3 = 4'd5;
b_sign0 = 4'd8; b_sign1 = 4'd7; b_sign2 = 4'd11; b_sign3 = 4'd15;
@(posedge clk_i);
a_mant0 = 8'd229; a_mant1 = 8'd164; a_mant2 = 8'd43; a_mant3 = 8'd170;
b_mant0 = 8'd94; b_mant1 = 8'd200; b_mant2 = 8'd167; b_mant3 = 8'd177;
a_exp0 = 10'd152; a_exp1 = 10'd821; a_exp2 = 10'd434; a_exp3 = 10'd709;
b_exp0 = 10'd90; b_exp1 = 10'd645; b_exp2 = 10'd166; b_exp3 = 10'd961;
a_sign0 = 4'd12; a_sign1 = 4'd4; a_sign2 = 4'd1; a_sign3 = 4'd3;
b_sign0 = 4'd10; b_sign1 = 4'd0; b_sign2 = 4'd3; b_sign3 = 4'd1;
@(posedge clk_i);
shared_exps0 = 8'd149;
shared_exps1 = 8'd118;
a_mant0 = 8'd43; a_mant1 = 8'd249; a_mant2 = 8'd224; a_mant3 = 8'd127;
b_mant0 = 8'd183; b_mant1 = 8'd156; b_mant2 = 8'd113; b_mant3 = 8'd36;
a_exp0 = 10'd289; a_exp1 = 10'd332; a_exp2 = 10'd872; a_exp3 = 10'd420;
b_exp0 = 10'd453; b_exp1 = 10'd41; b_exp2 = 10'd13; b_exp3 = 10'd514;
a_sign0 = 4'd9; a_sign1 = 4'd16; a_sign2 = 4'd1; a_sign3 = 4'd15;
b_sign0 = 4'd1; b_sign1 = 4'd5; b_sign2 = 4'd6; b_sign3 = 4'd5;
@(posedge clk_i);
a_mant0 = 8'd104; a_mant1 = 8'd133; a_mant2 = 8'd178; a_mant3 = 8'd124;
b_mant0 = 8'd96; b_mant1 = 8'd226; b_mant2 = 8'd46; b_mant3 = 8'd240;
a_exp0 = 10'd428; a_exp1 = 10'd489; a_exp2 = 10'd766; a_exp3 = 10'd785;
b_exp0 = 10'd12; b_exp1 = 10'd690; b_exp2 = 10'd483; b_exp3 = 10'd783;
a_sign0 = 4'd10; a_sign1 = 4'd5; a_sign2 = 4'd6; a_sign3 = 4'd15;
b_sign0 = 4'd9; b_sign1 = 4'd8; b_sign2 = 4'd3; b_sign3 = 4'd10;
@(posedge clk_i);
a_mant0 = 8'd105; a_mant1 = 8'd231; a_mant2 = 8'd243; a_mant3 = 8'd227;
b_mant0 = 8'd106; b_mant1 = 8'd254; b_mant2 = 8'd29; b_mant3 = 8'd2;
a_exp0 = 10'd919; a_exp1 = 10'd443; a_exp2 = 10'd119; a_exp3 = 10'd112;
b_exp0 = 10'd718; b_exp1 = 10'd235; b_exp2 = 10'd61; b_exp3 = 10'd313;
a_sign0 = 4'd10; a_sign1 = 4'd3; a_sign2 = 4'd16; a_sign3 = 4'd1;
b_sign0 = 4'd0; b_sign1 = 4'd8; b_sign2 = 4'd8; b_sign3 = 4'd16;
@(posedge clk_i);
a_mant0 = 8'd169; a_mant1 = 8'd220; a_mant2 = 8'd253; a_mant3 = 8'd13;
b_mant0 = 8'd22; b_mant1 = 8'd81; b_mant2 = 8'd173; b_mant3 = 8'd115;
a_exp0 = 10'd207; a_exp1 = 10'd756; a_exp2 = 10'd740; a_exp3 = 10'd703;
b_exp0 = 10'd534; b_exp1 = 10'd304; b_exp2 = 10'd55; b_exp3 = 10'd859;
a_sign0 = 4'd2; a_sign1 = 4'd15; a_sign2 = 4'd6; a_sign3 = 4'd14;
b_sign0 = 4'd10; b_sign1 = 4'd1; b_sign2 = 4'd11; b_sign3 = 4'd5;
@(posedge clk_i);
a_mant0 = 8'd68; a_mant1 = 8'd18; a_mant2 = 8'd63; a_mant3 = 8'd2;
b_mant0 = 8'd127; b_mant1 = 8'd128; b_mant2 = 8'd221; b_mant3 = 8'd65;
a_exp0 = 10'd343; a_exp1 = 10'd231; a_exp2 = 10'd378; a_exp3 = 10'd155;
b_exp0 = 10'd666; b_exp1 = 10'd829; b_exp2 = 10'd871; b_exp3 = 10'd683;
a_sign0 = 4'd14; a_sign1 = 4'd15; a_sign2 = 4'd1; a_sign3 = 4'd5;
b_sign0 = 4'd4; b_sign1 = 4'd3; b_sign2 = 4'd4; b_sign3 = 4'd8;
@(posedge clk_i);
a_mant0 = 8'd181; a_mant1 = 8'd6; a_mant2 = 8'd79; a_mant3 = 8'd210;
b_mant0 = 8'd76; b_mant1 = 8'd12; b_mant2 = 8'd156; b_mant3 = 8'd143;
a_exp0 = 10'd370; a_exp1 = 10'd487; a_exp2 = 10'd472; a_exp3 = 10'd118;
b_exp0 = 10'd719; b_exp1 = 10'd57; b_exp2 = 10'd570; b_exp3 = 10'd330;
a_sign0 = 4'd0; a_sign1 = 4'd13; a_sign2 = 4'd4; a_sign3 = 4'd8;
b_sign0 = 4'd0; b_sign1 = 4'd9; b_sign2 = 4'd16; b_sign3 = 4'd1;
@(posedge clk_i);
a_mant0 = 8'd88; a_mant1 = 8'd64; a_mant2 = 8'd224; a_mant3 = 8'd197;
b_mant0 = 8'd115; b_mant1 = 8'd90; b_mant2 = 8'd114; b_mant3 = 8'd170;
a_exp0 = 10'd285; a_exp1 = 10'd602; a_exp2 = 10'd949; a_exp3 = 10'd828;
b_exp0 = 10'd755; b_exp1 = 10'd374; b_exp2 = 10'd54; b_exp3 = 10'd742;
a_sign0 = 4'd0; a_sign1 = 4'd3; a_sign2 = 4'd16; a_sign3 = 4'd5;
b_sign0 = 4'd3; b_sign1 = 4'd5; b_sign2 = 4'd2; b_sign3 = 4'd16;
@(posedge clk_i);
a_mant0 = 8'd82; a_mant1 = 8'd64; a_mant2 = 8'd117; a_mant3 = 8'd3;
b_mant0 = 8'd132; b_mant1 = 8'd246; b_mant2 = 8'd30; b_mant3 = 8'd49;
a_exp0 = 10'd221; a_exp1 = 10'd320; a_exp2 = 10'd710; a_exp3 = 10'd538;
b_exp0 = 10'd899; b_exp1 = 10'd363; b_exp2 = 10'd800; b_exp3 = 10'd84;
a_sign0 = 4'd4; a_sign1 = 4'd15; a_sign2 = 4'd16; a_sign3 = 4'd15;
b_sign0 = 4'd3; b_sign1 = 4'd4; b_sign2 = 4'd2; b_sign3 = 4'd15;
@(posedge clk_i);
shared_exps0 = 8'd111;
shared_exps1 = 8'd110;
rstn = 0;
@(posedge clk_i);
rstn = 1;
a_mant0 = 8'd16; a_mant1 = 8'd84; a_mant2 = 8'd89; a_mant3 = 8'd176;
b_mant0 = 8'd158; b_mant1 = 8'd85; b_mant2 = 8'd251; b_mant3 = 8'd220;
a_exp0 = 10'd236; a_exp1 = 10'd141; a_exp2 = 10'd760; a_exp3 = 10'd704;
b_exp0 = 10'd922; b_exp1 = 10'd449; b_exp2 = 10'd21; b_exp3 = 10'd981;
a_sign0 = 4'd14; a_sign1 = 4'd6; a_sign2 = 4'd11; a_sign3 = 4'd15;
b_sign0 = 4'd12; b_sign1 = 4'd15; b_sign2 = 4'd3; b_sign3 = 4'd4;
@(posedge clk_i);
a_mant0 = 8'd3; a_mant1 = 8'd1; a_mant2 = 8'd168; a_mant3 = 8'd228;
b_mant0 = 8'd165; b_mant1 = 8'd91; b_mant2 = 8'd209; b_mant3 = 8'd27;
a_exp0 = 10'd141; a_exp1 = 10'd820; a_exp2 = 10'd272; a_exp3 = 10'd324;
b_exp0 = 10'd265; b_exp1 = 10'd432; b_exp2 = 10'd500; b_exp3 = 10'd337;
a_sign0 = 4'd15; a_sign1 = 4'd0; a_sign2 = 4'd9; a_sign3 = 4'd5;
b_sign0 = 4'd0; b_sign1 = 4'd13; b_sign2 = 4'd10; b_sign3 = 4'd3;
@(posedge clk_i);
a_mant0 = 8'd14; a_mant1 = 8'd36; a_mant2 = 8'd172; a_mant3 = 8'd105;
b_mant0 = 8'd17; b_mant1 = 8'd2; b_mant2 = 8'd190; b_mant3 = 8'd6;
a_exp0 = 10'd538; a_exp1 = 10'd211; a_exp2 = 10'd146; a_exp3 = 10'd545;
b_exp0 = 10'd950; b_exp1 = 10'd886; b_exp2 = 10'd896; b_exp3 = 10'd601;
a_sign0 = 4'd8; a_sign1 = 4'd11; a_sign2 = 4'd5; a_sign3 = 4'd11;
b_sign0 = 4'd3; b_sign1 = 4'd9; b_sign2 = 4'd9; b_sign3 = 4'd0;
@(posedge clk_i);
a_mant0 = 8'd247; a_mant1 = 8'd108; a_mant2 = 8'd97; a_mant3 = 8'd224;
b_mant0 = 8'd45; b_mant1 = 8'd215; b_mant2 = 8'd189; b_mant3 = 8'd94;
a_exp0 = 10'd429; a_exp1 = 10'd81; a_exp2 = 10'd487; a_exp3 = 10'd554;
b_exp0 = 10'd191; b_exp1 = 10'd162; b_exp2 = 10'd15; b_exp3 = 10'd1017;
a_sign0 = 4'd5; a_sign1 = 4'd12; a_sign2 = 4'd7; a_sign3 = 4'd7;
b_sign0 = 4'd0; b_sign1 = 4'd11; b_sign2 = 4'd8; b_sign3 = 4'd10;
@(posedge clk_i);
a_mant0 = 8'd39; a_mant1 = 8'd112; a_mant2 = 8'd111; a_mant3 = 8'd36;
b_mant0 = 8'd111; b_mant1 = 8'd246; b_mant2 = 8'd64; b_mant3 = 8'd120;
a_exp0 = 10'd17; a_exp1 = 10'd241; a_exp2 = 10'd623; a_exp3 = 10'd356;
b_exp0 = 10'd151; b_exp1 = 10'd886; b_exp2 = 10'd95; b_exp3 = 10'd73;
a_sign0 = 4'd7; a_sign1 = 4'd1; a_sign2 = 4'd9; a_sign3 = 4'd9;
b_sign0 = 4'd13; b_sign1 = 4'd4; b_sign2 = 4'd2; b_sign3 = 4'd1;
@(posedge clk_i);
a_mant0 = 8'd166; a_mant1 = 8'd96; a_mant2 = 8'd161; a_mant3 = 8'd131;
b_mant0 = 8'd63; b_mant1 = 8'd207; b_mant2 = 8'd11; b_mant3 = 8'd76;
a_exp0 = 10'd186; a_exp1 = 10'd715; a_exp2 = 10'd402; a_exp3 = 10'd593;
b_exp0 = 10'd947; b_exp1 = 10'd559; b_exp2 = 10'd264; b_exp3 = 10'd629;
a_sign0 = 4'd2; a_sign1 = 4'd12; a_sign2 = 4'd9; a_sign3 = 4'd0;
b_sign0 = 4'd3; b_sign1 = 4'd6; b_sign2 = 4'd5; b_sign3 = 4'd3;
@(posedge clk_i);
a_mant0 = 8'd170; a_mant1 = 8'd193; a_mant2 = 8'd11; a_mant3 = 8'd36;
b_mant0 = 8'd110; b_mant1 = 8'd208; b_mant2 = 8'd234; b_mant3 = 8'd21;
a_exp0 = 10'd829; a_exp1 = 10'd975; a_exp2 = 10'd43; a_exp3 = 10'd666;
b_exp0 = 10'd419; b_exp1 = 10'd442; b_exp2 = 10'd208; b_exp3 = 10'd77;
a_sign0 = 4'd2; a_sign1 = 4'd3; a_sign2 = 4'd8; a_sign3 = 4'd7;
b_sign0 = 4'd0; b_sign1 = 4'd11; b_sign2 = 4'd12; b_sign3 = 4'd7;
@(posedge clk_i);
shared_exps0 = 8'd135;
shared_exps1 = 8'd131;
a_mant0 = 8'd245; a_mant1 = 8'd232; a_mant2 = 8'd92; a_mant3 = 8'd34;
b_mant0 = 8'd177; b_mant1 = 8'd117; b_mant2 = 8'd168; b_mant3 = 8'd22;
a_exp0 = 10'd347; a_exp1 = 10'd1016; a_exp2 = 10'd14; a_exp3 = 10'd843;
b_exp0 = 10'd508; b_exp1 = 10'd294; b_exp2 = 10'd126; b_exp3 = 10'd611;
a_sign0 = 4'd12; a_sign1 = 4'd16; a_sign2 = 4'd0; a_sign3 = 4'd15;
b_sign0 = 4'd13; b_sign1 = 4'd16; b_sign2 = 4'd8; b_sign3 = 4'd0;
@(posedge clk_i);
a_mant0 = 8'd155; a_mant1 = 8'd233; a_mant2 = 8'd94; a_mant3 = 8'd58;
b_mant0 = 8'd1; b_mant1 = 8'd118; b_mant2 = 8'd188; b_mant3 = 8'd210;
a_exp0 = 10'd953; a_exp1 = 10'd801; a_exp2 = 10'd466; a_exp3 = 10'd229;
b_exp0 = 10'd289; b_exp1 = 10'd872; b_exp2 = 10'd146; b_exp3 = 10'd200;
a_sign0 = 4'd6; a_sign1 = 4'd13; a_sign2 = 4'd0; a_sign3 = 4'd9;
b_sign0 = 4'd9; b_sign1 = 4'd8; b_sign2 = 4'd2; b_sign3 = 4'd3;
@(posedge clk_i);
a_mant0 = 8'd255; a_mant1 = 8'd13; a_mant2 = 8'd245; a_mant3 = 8'd230;
b_mant0 = 8'd212; b_mant1 = 8'd126; b_mant2 = 8'd231; b_mant3 = 8'd31;
a_exp0 = 10'd306; a_exp1 = 10'd623; a_exp2 = 10'd374; a_exp3 = 10'd488;
b_exp0 = 10'd401; b_exp1 = 10'd286; b_exp2 = 10'd864; b_exp3 = 10'd748;
a_sign0 = 4'd13; a_sign1 = 4'd8; a_sign2 = 4'd14; a_sign3 = 4'd10;
b_sign0 = 4'd15; b_sign1 = 4'd5; b_sign2 = 4'd12; b_sign3 = 4'd1;
@(posedge clk_i);
a_mant0 = 8'd30; a_mant1 = 8'd92; a_mant2 = 8'd83; a_mant3 = 8'd126;
b_mant0 = 8'd183; b_mant1 = 8'd65; b_mant2 = 8'd201; b_mant3 = 8'd185;
a_exp0 = 10'd72; a_exp1 = 10'd969; a_exp2 = 10'd724; a_exp3 = 10'd284;
b_exp0 = 10'd307; b_exp1 = 10'd370; b_exp2 = 10'd986; b_exp3 = 10'd222;
a_sign0 = 4'd8; a_sign1 = 4'd13; a_sign2 = 4'd4; a_sign3 = 4'd1;
b_sign0 = 4'd5; b_sign1 = 4'd8; b_sign2 = 4'd9; b_sign3 = 4'd3;
@(posedge clk_i);
a_mant0 = 8'd88; a_mant1 = 8'd163; a_mant2 = 8'd35; a_mant3 = 8'd150;
b_mant0 = 8'd4; b_mant1 = 8'd164; b_mant2 = 8'd48; b_mant3 = 8'd7;
a_exp0 = 10'd347; a_exp1 = 10'd332; a_exp2 = 10'd155; a_exp3 = 10'd656;
b_exp0 = 10'd76; b_exp1 = 10'd793; b_exp2 = 10'd181; b_exp3 = 10'd760;
a_sign0 = 4'd0; a_sign1 = 4'd16; a_sign2 = 4'd8; a_sign3 = 4'd3;
b_sign0 = 4'd13; b_sign1 = 4'd7; b_sign2 = 4'd9; b_sign3 = 4'd8;
@(posedge clk_i);
a_mant0 = 8'd80; a_mant1 = 8'd156; a_mant2 = 8'd239; a_mant3 = 8'd48;
b_mant0 = 8'd166; b_mant1 = 8'd165; b_mant2 = 8'd164; b_mant3 = 8'd84;
a_exp0 = 10'd257; a_exp1 = 10'd852; a_exp2 = 10'd744; a_exp3 = 10'd283;
b_exp0 = 10'd137; b_exp1 = 10'd812; b_exp2 = 10'd344; b_exp3 = 10'd94;
a_sign0 = 4'd1; a_sign1 = 4'd3; a_sign2 = 4'd3; a_sign3 = 4'd5;
b_sign0 = 4'd0; b_sign1 = 4'd15; b_sign2 = 4'd2; b_sign3 = 4'd0;
@(posedge clk_i);
a_mant0 = 8'd24; a_mant1 = 8'd36; a_mant2 = 8'd29; a_mant3 = 8'd112;
b_mant0 = 8'd119; b_mant1 = 8'd61; b_mant2 = 8'd219; b_mant3 = 8'd208;
a_exp0 = 10'd100; a_exp1 = 10'd21; a_exp2 = 10'd456; a_exp3 = 10'd122;
b_exp0 = 10'd581; b_exp1 = 10'd670; b_exp2 = 10'd808; b_exp3 = 10'd894;
a_sign0 = 4'd14; a_sign1 = 4'd2; a_sign2 = 4'd4; a_sign3 = 4'd5;
b_sign0 = 4'd0; b_sign1 = 4'd0; b_sign2 = 4'd3; b_sign3 = 4'd3;
@(posedge clk_i);
a_mant0 = 8'd44; a_mant1 = 8'd122; a_mant2 = 8'd77; a_mant3 = 8'd6;
b_mant0 = 8'd209; b_mant1 = 8'd137; b_mant2 = 8'd156; b_mant3 = 8'd39;
a_exp0 = 10'd924; a_exp1 = 10'd447; a_exp2 = 10'd110; a_exp3 = 10'd152;
b_exp0 = 10'd974; b_exp1 = 10'd919; b_exp2 = 10'd366; b_exp3 = 10'd620;
a_sign0 = 4'd11; a_sign1 = 4'd3; a_sign2 = 4'd15; a_sign3 = 4'd6;
b_sign0 = 4'd12; b_sign1 = 4'd13; b_sign2 = 4'd14; b_sign3 = 4'd4;
@(posedge clk_i);
shared_exps0 = 8'd129;
shared_exps1 = 8'd111;
a_mant0 = 8'd206; a_mant1 = 8'd13; a_mant2 = 8'd129; a_mant3 = 8'd217;
b_mant0 = 8'd113; b_mant1 = 8'd27; b_mant2 = 8'd5; b_mant3 = 8'd186;
a_exp0 = 10'd584; a_exp1 = 10'd436; a_exp2 = 10'd738; a_exp3 = 10'd271;
b_exp0 = 10'd539; b_exp1 = 10'd242; b_exp2 = 10'd507; b_exp3 = 10'd932;
a_sign0 = 4'd16; a_sign1 = 4'd0; a_sign2 = 4'd0; a_sign3 = 4'd16;
b_sign0 = 4'd5; b_sign1 = 4'd10; b_sign2 = 4'd9; b_sign3 = 4'd0;
@(posedge clk_i);
a_mant0 = 8'd1; a_mant1 = 8'd224; a_mant2 = 8'd44; a_mant3 = 8'd137;
b_mant0 = 8'd69; b_mant1 = 8'd244; b_mant2 = 8'd111; b_mant3 = 8'd0;
a_exp0 = 10'd900; a_exp1 = 10'd601; a_exp2 = 10'd650; a_exp3 = 10'd991;
b_exp0 = 10'd110; b_exp1 = 10'd454; b_exp2 = 10'd632; b_exp3 = 10'd305;
a_sign0 = 4'd11; a_sign1 = 4'd15; a_sign2 = 4'd11; a_sign3 = 4'd15;
b_sign0 = 4'd16; b_sign1 = 4'd12; b_sign2 = 4'd2; b_sign3 = 4'd11;
@(posedge clk_i);
a_mant0 = 8'd86; a_mant1 = 8'd228; a_mant2 = 8'd69; a_mant3 = 8'd136;
b_mant0 = 8'd95; b_mant1 = 8'd75; b_mant2 = 8'd235; b_mant3 = 8'd58;
a_exp0 = 10'd603; a_exp1 = 10'd322; a_exp2 = 10'd531; a_exp3 = 10'd731;
b_exp0 = 10'd949; b_exp1 = 10'd434; b_exp2 = 10'd134; b_exp3 = 10'd980;
a_sign0 = 4'd0; a_sign1 = 4'd13; a_sign2 = 4'd3; a_sign3 = 4'd7;
b_sign0 = 4'd0; b_sign1 = 4'd16; b_sign2 = 4'd11; b_sign3 = 4'd11;
@(posedge clk_i);
a_mant0 = 8'd12; a_mant1 = 8'd127; a_mant2 = 8'd44; a_mant3 = 8'd199;
b_mant0 = 8'd223; b_mant1 = 8'd90; b_mant2 = 8'd59; b_mant3 = 8'd215;
a_exp0 = 10'd568; a_exp1 = 10'd620; a_exp2 = 10'd398; a_exp3 = 10'd540;
b_exp0 = 10'd505; b_exp1 = 10'd695; b_exp2 = 10'd37; b_exp3 = 10'd884;
a_sign0 = 4'd8; a_sign1 = 4'd16; a_sign2 = 4'd1; a_sign3 = 4'd16;
b_sign0 = 4'd14; b_sign1 = 4'd4; b_sign2 = 4'd3; b_sign3 = 4'd8;
@(posedge clk_i);
a_mant0 = 8'd78; a_mant1 = 8'd192; a_mant2 = 8'd242; a_mant3 = 8'd115;
b_mant0 = 8'd119; b_mant1 = 8'd109; b_mant2 = 8'd103; b_mant3 = 8'd174;
a_exp0 = 10'd180; a_exp1 = 10'd393; a_exp2 = 10'd329; a_exp3 = 10'd748;
b_exp0 = 10'd55; b_exp1 = 10'd244; b_exp2 = 10'd556; b_exp3 = 10'd204;
a_sign0 = 4'd4; a_sign1 = 4'd8; a_sign2 = 4'd12; a_sign3 = 4'd9;
b_sign0 = 4'd13; b_sign1 = 4'd10; b_sign2 = 4'd0; b_sign3 = 4'd13;
@(posedge clk_i);
a_mant0 = 8'd251; a_mant1 = 8'd165; a_mant2 = 8'd251; a_mant3 = 8'd151;
b_mant0 = 8'd6; b_mant1 = 8'd85; b_mant2 = 8'd28; b_mant3 = 8'd133;
a_exp0 = 10'd399; a_exp1 = 10'd1009; a_exp2 = 10'd713; a_exp3 = 10'd628;
b_exp0 = 10'd579; b_exp1 = 10'd986; b_exp2 = 10'd262; b_exp3 = 10'd19;
a_sign0 = 4'd8; a_sign1 = 4'd5; a_sign2 = 4'd12; a_sign3 = 4'd4;
b_sign0 = 4'd16; b_sign1 = 4'd16; b_sign2 = 4'd16; b_sign3 = 4'd9;
@(posedge clk_i);
a_mant0 = 8'd249; a_mant1 = 8'd104; a_mant2 = 8'd87; a_mant3 = 8'd239;
b_mant0 = 8'd106; b_mant1 = 8'd238; b_mant2 = 8'd246; b_mant3 = 8'd163;
a_exp0 = 10'd430; a_exp1 = 10'd17; a_exp2 = 10'd559; a_exp3 = 10'd784;
b_exp0 = 10'd60; b_exp1 = 10'd160; b_exp2 = 10'd1009; b_exp3 = 10'd940;
a_sign0 = 4'd2; a_sign1 = 4'd15; a_sign2 = 4'd7; a_sign3 = 4'd12;
b_sign0 = 4'd1; b_sign1 = 4'd8; b_sign2 = 4'd0; b_sign3 = 4'd12;
@(posedge clk_i);
a_mant0 = 8'd106; a_mant1 = 8'd196; a_mant2 = 8'd120; a_mant3 = 8'd187;
b_mant0 = 8'd247; b_mant1 = 8'd154; b_mant2 = 8'd40; b_mant3 = 8'd116;
a_exp0 = 10'd531; a_exp1 = 10'd819; a_exp2 = 10'd270; a_exp3 = 10'd232;
b_exp0 = 10'd623; b_exp1 = 10'd725; b_exp2 = 10'd419; b_exp3 = 10'd472;
a_sign0 = 4'd9; a_sign1 = 4'd15; a_sign2 = 4'd8; a_sign3 = 4'd15;
b_sign0 = 4'd1; b_sign1 = 4'd0; b_sign2 = 4'd2; b_sign3 = 4'd3;
@(posedge clk_i);
shared_exps0 = 8'd155;
shared_exps1 = 8'd126;
a_mant0 = 8'd177; a_mant1 = 8'd22; a_mant2 = 8'd246; a_mant3 = 8'd241;
b_mant0 = 8'd254; b_mant1 = 8'd186; b_mant2 = 8'd121; b_mant3 = 8'd163;
a_exp0 = 10'd944; a_exp1 = 10'd502; a_exp2 = 10'd658; a_exp3 = 10'd260;
b_exp0 = 10'd415; b_exp1 = 10'd664; b_exp2 = 10'd978; b_exp3 = 10'd675;
a_sign0 = 4'd9; a_sign1 = 4'd1; a_sign2 = 4'd10; a_sign3 = 4'd6;
b_sign0 = 4'd2; b_sign1 = 4'd10; b_sign2 = 4'd3; b_sign3 = 4'd2;
@(posedge clk_i);
a_mant0 = 8'd73; a_mant1 = 8'd210; a_mant2 = 8'd216; a_mant3 = 8'd46;
b_mant0 = 8'd179; b_mant1 = 8'd28; b_mant2 = 8'd198; b_mant3 = 8'd4;
a_exp0 = 10'd489; a_exp1 = 10'd299; a_exp2 = 10'd398; a_exp3 = 10'd209;
b_exp0 = 10'd156; b_exp1 = 10'd148; b_exp2 = 10'd294; b_exp3 = 10'd422;
a_sign0 = 4'd6; a_sign1 = 4'd9; a_sign2 = 4'd12; a_sign3 = 4'd14;
b_sign0 = 4'd0; b_sign1 = 4'd7; b_sign2 = 4'd16; b_sign3 = 4'd0;
@(posedge clk_i);
a_mant0 = 8'd142; a_mant1 = 8'd45; a_mant2 = 8'd112; a_mant3 = 8'd236;
b_mant0 = 8'd163; b_mant1 = 8'd114; b_mant2 = 8'd84; b_mant3 = 8'd118;
a_exp0 = 10'd508; a_exp1 = 10'd177; a_exp2 = 10'd225; a_exp3 = 10'd68;
b_exp0 = 10'd136; b_exp1 = 10'd420; b_exp2 = 10'd530; b_exp3 = 10'd721;
a_sign0 = 4'd15; a_sign1 = 4'd4; a_sign2 = 4'd2; a_sign3 = 4'd7;
b_sign0 = 4'd14; b_sign1 = 4'd10; b_sign2 = 4'd15; b_sign3 = 4'd4;
@(posedge clk_i);
a_mant0 = 8'd246; a_mant1 = 8'd20; a_mant2 = 8'd83; a_mant3 = 8'd57;
b_mant0 = 8'd209; b_mant1 = 8'd153; b_mant2 = 8'd235; b_mant3 = 8'd111;
a_exp0 = 10'd114; a_exp1 = 10'd282; a_exp2 = 10'd151; a_exp3 = 10'd620;
b_exp0 = 10'd716; b_exp1 = 10'd567; b_exp2 = 10'd534; b_exp3 = 10'd420;
a_sign0 = 4'd8; a_sign1 = 4'd9; a_sign2 = 4'd9; a_sign3 = 4'd6;
b_sign0 = 4'd8; b_sign1 = 4'd5; b_sign2 = 4'd3; b_sign3 = 4'd11;
@(posedge clk_i);
a_mant0 = 8'd128; a_mant1 = 8'd142; a_mant2 = 8'd199; a_mant3 = 8'd0;
b_mant0 = 8'd202; b_mant1 = 8'd101; b_mant2 = 8'd63; b_mant3 = 8'd19;
a_exp0 = 10'd158; a_exp1 = 10'd634; a_exp2 = 10'd651; a_exp3 = 10'd482;
b_exp0 = 10'd305; b_exp1 = 10'd449; b_exp2 = 10'd890; b_exp3 = 10'd139;
a_sign0 = 4'd4; a_sign1 = 4'd7; a_sign2 = 4'd1; a_sign3 = 4'd10;
b_sign0 = 4'd5; b_sign1 = 4'd14; b_sign2 = 4'd3; b_sign3 = 4'd2;
@(posedge clk_i);
a_mant0 = 8'd38; a_mant1 = 8'd134; a_mant2 = 8'd124; a_mant3 = 8'd25;
b_mant0 = 8'd156; b_mant1 = 8'd122; b_mant2 = 8'd99; b_mant3 = 8'd2;
a_exp0 = 10'd127; a_exp1 = 10'd101; a_exp2 = 10'd682; a_exp3 = 10'd150;
b_exp0 = 10'd508; b_exp1 = 10'd86; b_exp2 = 10'd714; b_exp3 = 10'd814;
a_sign0 = 4'd5; a_sign1 = 4'd3; a_sign2 = 4'd7; a_sign3 = 4'd5;
b_sign0 = 4'd8; b_sign1 = 4'd10; b_sign2 = 4'd11; b_sign3 = 4'd12;
@(posedge clk_i);
a_mant0 = 8'd79; a_mant1 = 8'd233; a_mant2 = 8'd1; a_mant3 = 8'd214;
b_mant0 = 8'd49; b_mant1 = 8'd117; b_mant2 = 8'd141; b_mant3 = 8'd185;
a_exp0 = 10'd545; a_exp1 = 10'd0; a_exp2 = 10'd409; a_exp3 = 10'd390;
b_exp0 = 10'd598; b_exp1 = 10'd228; b_exp2 = 10'd821; b_exp3 = 10'd674;
a_sign0 = 4'd3; a_sign1 = 4'd5; a_sign2 = 4'd6; a_sign3 = 4'd5;
b_sign0 = 4'd6; b_sign1 = 4'd3; b_sign2 = 4'd1; b_sign3 = 4'd4;
@(posedge clk_i);
a_mant0 = 8'd135; a_mant1 = 8'd235; a_mant2 = 8'd64; a_mant3 = 8'd21;
b_mant0 = 8'd227; b_mant1 = 8'd12; b_mant2 = 8'd38; b_mant3 = 8'd234;
a_exp0 = 10'd89; a_exp1 = 10'd987; a_exp2 = 10'd951; a_exp3 = 10'd320;
b_exp0 = 10'd408; b_exp1 = 10'd187; b_exp2 = 10'd657; b_exp3 = 10'd170;
a_sign0 = 4'd12; a_sign1 = 4'd14; a_sign2 = 4'd11; a_sign3 = 4'd12;
b_sign0 = 4'd5; b_sign1 = 4'd14; b_sign2 = 4'd12; b_sign3 = 4'd3;
@(posedge clk_i);
shared_exps0 = 8'd108;
shared_exps1 = 8'd105;
rstn = 0;
@(posedge clk_i);
rstn = 1;
a_mant0 = 8'd160; a_mant1 = 8'd167; a_mant2 = 8'd251; a_mant3 = 8'd176;
b_mant0 = 8'd13; b_mant1 = 8'd52; b_mant2 = 8'd234; b_mant3 = 8'd166;
a_exp0 = 10'd652; a_exp1 = 10'd298; a_exp2 = 10'd530; a_exp3 = 10'd438;
b_exp0 = 10'd955; b_exp1 = 10'd288; b_exp2 = 10'd507; b_exp3 = 10'd793;
a_sign0 = 4'd6; a_sign1 = 4'd2; a_sign2 = 4'd10; a_sign3 = 4'd15;
b_sign0 = 4'd3; b_sign1 = 4'd13; b_sign2 = 4'd3; b_sign3 = 4'd8;
@(posedge clk_i);
a_mant0 = 8'd238; a_mant1 = 8'd180; a_mant2 = 8'd64; a_mant3 = 8'd198;
b_mant0 = 8'd43; b_mant1 = 8'd144; b_mant2 = 8'd71; b_mant3 = 8'd230;
a_exp0 = 10'd757; a_exp1 = 10'd34; a_exp2 = 10'd542; a_exp3 = 10'd709;
b_exp0 = 10'd2; b_exp1 = 10'd430; b_exp2 = 10'd731; b_exp3 = 10'd850;
a_sign0 = 4'd2; a_sign1 = 4'd1; a_sign2 = 4'd13; a_sign3 = 4'd8;
b_sign0 = 4'd3; b_sign1 = 4'd6; b_sign2 = 4'd3; b_sign3 = 4'd5;
@(posedge clk_i);
a_mant0 = 8'd231; a_mant1 = 8'd230; a_mant2 = 8'd180; a_mant3 = 8'd80;
b_mant0 = 8'd117; b_mant1 = 8'd71; b_mant2 = 8'd97; b_mant3 = 8'd226;
a_exp0 = 10'd258; a_exp1 = 10'd758; a_exp2 = 10'd424; a_exp3 = 10'd357;
b_exp0 = 10'd889; b_exp1 = 10'd607; b_exp2 = 10'd33; b_exp3 = 10'd607;
a_sign0 = 4'd16; a_sign1 = 4'd15; a_sign2 = 4'd10; a_sign3 = 4'd1;
b_sign0 = 4'd9; b_sign1 = 4'd4; b_sign2 = 4'd8; b_sign3 = 4'd3;
@(posedge clk_i);
a_mant0 = 8'd246; a_mant1 = 8'd181; a_mant2 = 8'd163; a_mant3 = 8'd121;
b_mant0 = 8'd108; b_mant1 = 8'd101; b_mant2 = 8'd62; b_mant3 = 8'd139;
a_exp0 = 10'd456; a_exp1 = 10'd628; a_exp2 = 10'd313; a_exp3 = 10'd302;
b_exp0 = 10'd371; b_exp1 = 10'd769; b_exp2 = 10'd391; b_exp3 = 10'd749;
a_sign0 = 4'd1; a_sign1 = 4'd12; a_sign2 = 4'd10; a_sign3 = 4'd13;
b_sign0 = 4'd8; b_sign1 = 4'd2; b_sign2 = 4'd1; b_sign3 = 4'd15;
@(posedge clk_i);
a_mant0 = 8'd232; a_mant1 = 8'd247; a_mant2 = 8'd56; a_mant3 = 8'd202;
b_mant0 = 8'd190; b_mant1 = 8'd31; b_mant2 = 8'd152; b_mant3 = 8'd125;
a_exp0 = 10'd982; a_exp1 = 10'd163; a_exp2 = 10'd84; a_exp3 = 10'd283;
b_exp0 = 10'd908; b_exp1 = 10'd270; b_exp2 = 10'd786; b_exp3 = 10'd929;
a_sign0 = 4'd12; a_sign1 = 4'd10; a_sign2 = 4'd1; a_sign3 = 4'd5;
b_sign0 = 4'd2; b_sign1 = 4'd12; b_sign2 = 4'd11; b_sign3 = 4'd1;
@(posedge clk_i);
a_mant0 = 8'd50; a_mant1 = 8'd209; a_mant2 = 8'd152; a_mant3 = 8'd76;
b_mant0 = 8'd113; b_mant1 = 8'd225; b_mant2 = 8'd60; b_mant3 = 8'd22;
a_exp0 = 10'd585; a_exp1 = 10'd104; a_exp2 = 10'd456; a_exp3 = 10'd72;
b_exp0 = 10'd341; b_exp1 = 10'd359; b_exp2 = 10'd636; b_exp3 = 10'd777;
a_sign0 = 4'd9; a_sign1 = 4'd6; a_sign2 = 4'd7; a_sign3 = 4'd1;
b_sign0 = 4'd4; b_sign1 = 4'd15; b_sign2 = 4'd1; b_sign3 = 4'd15;
@(posedge clk_i);
a_mant0 = 8'd82; a_mant1 = 8'd154; a_mant2 = 8'd33; a_mant3 = 8'd51;
b_mant0 = 8'd160; b_mant1 = 8'd197; b_mant2 = 8'd26; b_mant3 = 8'd24;
a_exp0 = 10'd978; a_exp1 = 10'd195; a_exp2 = 10'd701; a_exp3 = 10'd560;
b_exp0 = 10'd495; b_exp1 = 10'd1; b_exp2 = 10'd768; b_exp3 = 10'd618;
a_sign0 = 4'd14; a_sign1 = 4'd1; a_sign2 = 4'd9; a_sign3 = 4'd10;
b_sign0 = 4'd4; b_sign1 = 4'd11; b_sign2 = 4'd3; b_sign3 = 4'd0;
@(posedge clk_i);
shared_exps0 = 8'd130;
shared_exps1 = 8'd116;
a_mant0 = 8'd166; a_mant1 = 8'd162; a_mant2 = 8'd25; a_mant3 = 8'd189;
b_mant0 = 8'd25; b_mant1 = 8'd226; b_mant2 = 8'd147; b_mant3 = 8'd3;
a_exp0 = 10'd78; a_exp1 = 10'd295; a_exp2 = 10'd716; a_exp3 = 10'd395;
b_exp0 = 10'd767; b_exp1 = 10'd86; b_exp2 = 10'd311; b_exp3 = 10'd619;
a_sign0 = 4'd0; a_sign1 = 4'd3; a_sign2 = 4'd8; a_sign3 = 4'd15;
b_sign0 = 4'd3; b_sign1 = 4'd5; b_sign2 = 4'd12; b_sign3 = 4'd13;
@(posedge clk_i);
a_mant0 = 8'd218; a_mant1 = 8'd226; a_mant2 = 8'd82; a_mant3 = 8'd57;
b_mant0 = 8'd82; b_mant1 = 8'd48; b_mant2 = 8'd237; b_mant3 = 8'd56;
a_exp0 = 10'd485; a_exp1 = 10'd736; a_exp2 = 10'd510; a_exp3 = 10'd518;
b_exp0 = 10'd336; b_exp1 = 10'd387; b_exp2 = 10'd691; b_exp3 = 10'd56;
a_sign0 = 4'd7; a_sign1 = 4'd6; a_sign2 = 4'd5; a_sign3 = 4'd9;
b_sign0 = 4'd16; b_sign1 = 4'd10; b_sign2 = 4'd16; b_sign3 = 4'd2;
@(posedge clk_i);
a_mant0 = 8'd138; a_mant1 = 8'd80; a_mant2 = 8'd133; a_mant3 = 8'd188;
b_mant0 = 8'd81; b_mant1 = 8'd146; b_mant2 = 8'd31; b_mant3 = 8'd158;
a_exp0 = 10'd226; a_exp1 = 10'd350; a_exp2 = 10'd679; a_exp3 = 10'd712;
b_exp0 = 10'd705; b_exp1 = 10'd714; b_exp2 = 10'd746; b_exp3 = 10'd25;
a_sign0 = 4'd14; a_sign1 = 4'd16; a_sign2 = 4'd0; a_sign3 = 4'd4;
b_sign0 = 4'd3; b_sign1 = 4'd7; b_sign2 = 4'd2; b_sign3 = 4'd14;
@(posedge clk_i);
a_mant0 = 8'd54; a_mant1 = 8'd77; a_mant2 = 8'd60; a_mant3 = 8'd229;
b_mant0 = 8'd230; b_mant1 = 8'd31; b_mant2 = 8'd62; b_mant3 = 8'd207;
a_exp0 = 10'd377; a_exp1 = 10'd835; a_exp2 = 10'd184; a_exp3 = 10'd531;
b_exp0 = 10'd608; b_exp1 = 10'd660; b_exp2 = 10'd337; b_exp3 = 10'd572;
a_sign0 = 4'd11; a_sign1 = 4'd4; a_sign2 = 4'd13; a_sign3 = 4'd5;
b_sign0 = 4'd12; b_sign1 = 4'd6; b_sign2 = 4'd2; b_sign3 = 4'd13;
@(posedge clk_i);
a_mant0 = 8'd21; a_mant1 = 8'd114; a_mant2 = 8'd100; a_mant3 = 8'd49;
b_mant0 = 8'd221; b_mant1 = 8'd92; b_mant2 = 8'd10; b_mant3 = 8'd82;
a_exp0 = 10'd672; a_exp1 = 10'd311; a_exp2 = 10'd182; a_exp3 = 10'd761;
b_exp0 = 10'd768; b_exp1 = 10'd757; b_exp2 = 10'd714; b_exp3 = 10'd129;
a_sign0 = 4'd14; a_sign1 = 4'd3; a_sign2 = 4'd11; a_sign3 = 4'd5;
b_sign0 = 4'd12; b_sign1 = 4'd0; b_sign2 = 4'd1; b_sign3 = 4'd11;
@(posedge clk_i);
a_mant0 = 8'd129; a_mant1 = 8'd169; a_mant2 = 8'd93; a_mant3 = 8'd243;
b_mant0 = 8'd30; b_mant1 = 8'd38; b_mant2 = 8'd15; b_mant3 = 8'd176;
a_exp0 = 10'd692; a_exp1 = 10'd349; a_exp2 = 10'd434; a_exp3 = 10'd721;
b_exp0 = 10'd210; b_exp1 = 10'd491; b_exp2 = 10'd214; b_exp3 = 10'd262;
a_sign0 = 4'd9; a_sign1 = 4'd10; a_sign2 = 4'd15; a_sign3 = 4'd4;
b_sign0 = 4'd2; b_sign1 = 4'd10; b_sign2 = 4'd3; b_sign3 = 4'd15;
@(posedge clk_i);
a_mant0 = 8'd160; a_mant1 = 8'd123; a_mant2 = 8'd160; a_mant3 = 8'd68;
b_mant0 = 8'd222; b_mant1 = 8'd156; b_mant2 = 8'd233; b_mant3 = 8'd12;
a_exp0 = 10'd444; a_exp1 = 10'd997; a_exp2 = 10'd854; a_exp3 = 10'd803;
b_exp0 = 10'd434; b_exp1 = 10'd296; b_exp2 = 10'd681; b_exp3 = 10'd39;
a_sign0 = 4'd12; a_sign1 = 4'd16; a_sign2 = 4'd13; a_sign3 = 4'd0;
b_sign0 = 4'd14; b_sign1 = 4'd10; b_sign2 = 4'd0; b_sign3 = 4'd12;
@(posedge clk_i);
a_mant0 = 8'd21; a_mant1 = 8'd57; a_mant2 = 8'd135; a_mant3 = 8'd253;
b_mant0 = 8'd20; b_mant1 = 8'd217; b_mant2 = 8'd161; b_mant3 = 8'd227;
a_exp0 = 10'd733; a_exp1 = 10'd833; a_exp2 = 10'd407; a_exp3 = 10'd27;
b_exp0 = 10'd887; b_exp1 = 10'd874; b_exp2 = 10'd666; b_exp3 = 10'd791;
a_sign0 = 4'd15; a_sign1 = 4'd15; a_sign2 = 4'd16; a_sign3 = 4'd15;
b_sign0 = 4'd7; b_sign1 = 4'd15; b_sign2 = 4'd13; b_sign3 = 4'd0;
@(posedge clk_i);
shared_exps0 = 8'd131;
shared_exps1 = 8'd118;
a_mant0 = 8'd162; a_mant1 = 8'd38; a_mant2 = 8'd246; a_mant3 = 8'd102;
b_mant0 = 8'd9; b_mant1 = 8'd171; b_mant2 = 8'd55; b_mant3 = 8'd74;
a_exp0 = 10'd510; a_exp1 = 10'd165; a_exp2 = 10'd12; a_exp3 = 10'd339;
b_exp0 = 10'd736; b_exp1 = 10'd303; b_exp2 = 10'd523; b_exp3 = 10'd371;
a_sign0 = 4'd1; a_sign1 = 4'd7; a_sign2 = 4'd5; a_sign3 = 4'd4;
b_sign0 = 4'd10; b_sign1 = 4'd9; b_sign2 = 4'd8; b_sign3 = 4'd10;
@(posedge clk_i);
a_mant0 = 8'd103; a_mant1 = 8'd145; a_mant2 = 8'd153; a_mant3 = 8'd209;
b_mant0 = 8'd8; b_mant1 = 8'd133; b_mant2 = 8'd212; b_mant3 = 8'd84;
a_exp0 = 10'd169; a_exp1 = 10'd321; a_exp2 = 10'd307; a_exp3 = 10'd106;
b_exp0 = 10'd851; b_exp1 = 10'd645; b_exp2 = 10'd939; b_exp3 = 10'd410;
a_sign0 = 4'd6; a_sign1 = 4'd3; a_sign2 = 4'd12; a_sign3 = 4'd5;
b_sign0 = 4'd13; b_sign1 = 4'd3; b_sign2 = 4'd2; b_sign3 = 4'd10;
@(posedge clk_i);
a_mant0 = 8'd171; a_mant1 = 8'd196; a_mant2 = 8'd82; a_mant3 = 8'd224;
b_mant0 = 8'd6; b_mant1 = 8'd110; b_mant2 = 8'd220; b_mant3 = 8'd36;
a_exp0 = 10'd89; a_exp1 = 10'd446; a_exp2 = 10'd694; a_exp3 = 10'd872;
b_exp0 = 10'd418; b_exp1 = 10'd148; b_exp2 = 10'd315; b_exp3 = 10'd730;
a_sign0 = 4'd14; a_sign1 = 4'd8; a_sign2 = 4'd0; a_sign3 = 4'd5;
b_sign0 = 4'd1; b_sign1 = 4'd8; b_sign2 = 4'd2; b_sign3 = 4'd9;
@(posedge clk_i);
a_mant0 = 8'd238; a_mant1 = 8'd167; a_mant2 = 8'd13; a_mant3 = 8'd85;
b_mant0 = 8'd37; b_mant1 = 8'd238; b_mant2 = 8'd204; b_mant3 = 8'd198;
a_exp0 = 10'd674; a_exp1 = 10'd272; a_exp2 = 10'd741; a_exp3 = 10'd1022;
b_exp0 = 10'd134; b_exp1 = 10'd175; b_exp2 = 10'd371; b_exp3 = 10'd815;
a_sign0 = 4'd7; a_sign1 = 4'd2; a_sign2 = 4'd3; a_sign3 = 4'd1;
b_sign0 = 4'd7; b_sign1 = 4'd7; b_sign2 = 4'd10; b_sign3 = 4'd12;
@(posedge clk_i);
a_mant0 = 8'd66; a_mant1 = 8'd219; a_mant2 = 8'd85; a_mant3 = 8'd247;
b_mant0 = 8'd60; b_mant1 = 8'd53; b_mant2 = 8'd91; b_mant3 = 8'd239;
a_exp0 = 10'd943; a_exp1 = 10'd728; a_exp2 = 10'd943; a_exp3 = 10'd24;
b_exp0 = 10'd449; b_exp1 = 10'd748; b_exp2 = 10'd469; b_exp3 = 10'd787;
a_sign0 = 4'd3; a_sign1 = 4'd15; a_sign2 = 4'd15; a_sign3 = 4'd12;
b_sign0 = 4'd6; b_sign1 = 4'd11; b_sign2 = 4'd8; b_sign3 = 4'd3;
@(posedge clk_i);
a_mant0 = 8'd151; a_mant1 = 8'd143; a_mant2 = 8'd85; a_mant3 = 8'd60;
b_mant0 = 8'd126; b_mant1 = 8'd157; b_mant2 = 8'd188; b_mant3 = 8'd152;
a_exp0 = 10'd901; a_exp1 = 10'd186; a_exp2 = 10'd937; a_exp3 = 10'd777;
b_exp0 = 10'd982; b_exp1 = 10'd346; b_exp2 = 10'd505; b_exp3 = 10'd325;
a_sign0 = 4'd3; a_sign1 = 4'd6; a_sign2 = 4'd4; a_sign3 = 4'd16;
b_sign0 = 4'd15; b_sign1 = 4'd8; b_sign2 = 4'd4; b_sign3 = 4'd8;
@(posedge clk_i);
a_mant0 = 8'd2; a_mant1 = 8'd59; a_mant2 = 8'd99; a_mant3 = 8'd184;
b_mant0 = 8'd122; b_mant1 = 8'd60; b_mant2 = 8'd114; b_mant3 = 8'd119;
a_exp0 = 10'd659; a_exp1 = 10'd892; a_exp2 = 10'd370; a_exp3 = 10'd909;
b_exp0 = 10'd24; b_exp1 = 10'd421; b_exp2 = 10'd80; b_exp3 = 10'd193;
a_sign0 = 4'd15; a_sign1 = 4'd5; a_sign2 = 4'd8; a_sign3 = 4'd6;
b_sign0 = 4'd12; b_sign1 = 4'd16; b_sign2 = 4'd4; b_sign3 = 4'd0;
@(posedge clk_i);
a_mant0 = 8'd84; a_mant1 = 8'd84; a_mant2 = 8'd110; a_mant3 = 8'd46;
b_mant0 = 8'd252; b_mant1 = 8'd236; b_mant2 = 8'd157; b_mant3 = 8'd158;
a_exp0 = 10'd80; a_exp1 = 10'd63; a_exp2 = 10'd732; a_exp3 = 10'd883;
b_exp0 = 10'd369; b_exp1 = 10'd292; b_exp2 = 10'd584; b_exp3 = 10'd224;
a_sign0 = 4'd4; a_sign1 = 4'd7; a_sign2 = 4'd14; a_sign3 = 4'd1;
b_sign0 = 4'd11; b_sign1 = 4'd16; b_sign2 = 4'd2; b_sign3 = 4'd13;
@(posedge clk_i);
shared_exps0 = 8'd116;
shared_exps1 = 8'd161;
a_mant0 = 8'd14; a_mant1 = 8'd119; a_mant2 = 8'd145; a_mant3 = 8'd118;
b_mant0 = 8'd253; b_mant1 = 8'd9; b_mant2 = 8'd97; b_mant3 = 8'd201;
a_exp0 = 10'd920; a_exp1 = 10'd810; a_exp2 = 10'd675; a_exp3 = 10'd318;
b_exp0 = 10'd402; b_exp1 = 10'd174; b_exp2 = 10'd472; b_exp3 = 10'd16;
a_sign0 = 4'd6; a_sign1 = 4'd6; a_sign2 = 4'd4; a_sign3 = 4'd16;
b_sign0 = 4'd5; b_sign1 = 4'd13; b_sign2 = 4'd11; b_sign3 = 4'd13;
@(posedge clk_i);
a_mant0 = 8'd244; a_mant1 = 8'd212; a_mant2 = 8'd25; a_mant3 = 8'd134;
b_mant0 = 8'd217; b_mant1 = 8'd190; b_mant2 = 8'd253; b_mant3 = 8'd198;
a_exp0 = 10'd621; a_exp1 = 10'd1012; a_exp2 = 10'd639; a_exp3 = 10'd23;
b_exp0 = 10'd59; b_exp1 = 10'd443; b_exp2 = 10'd929; b_exp3 = 10'd156;
a_sign0 = 4'd12; a_sign1 = 4'd2; a_sign2 = 4'd0; a_sign3 = 4'd0;
b_sign0 = 4'd4; b_sign1 = 4'd8; b_sign2 = 4'd3; b_sign3 = 4'd3;
@(posedge clk_i);
a_mant0 = 8'd222; a_mant1 = 8'd141; a_mant2 = 8'd155; a_mant3 = 8'd247;
b_mant0 = 8'd241; b_mant1 = 8'd105; b_mant2 = 8'd81; b_mant3 = 8'd132;
a_exp0 = 10'd40; a_exp1 = 10'd67; a_exp2 = 10'd170; a_exp3 = 10'd15;
b_exp0 = 10'd204; b_exp1 = 10'd231; b_exp2 = 10'd724; b_exp3 = 10'd567;
a_sign0 = 4'd5; a_sign1 = 4'd0; a_sign2 = 4'd12; a_sign3 = 4'd10;
b_sign0 = 4'd12; b_sign1 = 4'd1; b_sign2 = 4'd14; b_sign3 = 4'd14;
@(posedge clk_i);
a_mant0 = 8'd147; a_mant1 = 8'd85; a_mant2 = 8'd232; a_mant3 = 8'd48;
b_mant0 = 8'd152; b_mant1 = 8'd122; b_mant2 = 8'd116; b_mant3 = 8'd26;
a_exp0 = 10'd968; a_exp1 = 10'd888; a_exp2 = 10'd93; a_exp3 = 10'd635;
b_exp0 = 10'd624; b_exp1 = 10'd570; b_exp2 = 10'd979; b_exp3 = 10'd645;
a_sign0 = 4'd4; a_sign1 = 4'd4; a_sign2 = 4'd0; a_sign3 = 4'd4;
b_sign0 = 4'd15; b_sign1 = 4'd14; b_sign2 = 4'd4; b_sign3 = 4'd6;
@(posedge clk_i);
a_mant0 = 8'd129; a_mant1 = 8'd168; a_mant2 = 8'd195; a_mant3 = 8'd44;
b_mant0 = 8'd97; b_mant1 = 8'd185; b_mant2 = 8'd213; b_mant3 = 8'd5;
a_exp0 = 10'd423; a_exp1 = 10'd922; a_exp2 = 10'd135; a_exp3 = 10'd792;
b_exp0 = 10'd242; b_exp1 = 10'd36; b_exp2 = 10'd586; b_exp3 = 10'd829;
a_sign0 = 4'd12; a_sign1 = 4'd0; a_sign2 = 4'd3; a_sign3 = 4'd13;
b_sign0 = 4'd15; b_sign1 = 4'd10; b_sign2 = 4'd1; b_sign3 = 4'd8;
@(posedge clk_i);
a_mant0 = 8'd121; a_mant1 = 8'd106; a_mant2 = 8'd40; a_mant3 = 8'd62;
b_mant0 = 8'd50; b_mant1 = 8'd212; b_mant2 = 8'd113; b_mant3 = 8'd251;
a_exp0 = 10'd938; a_exp1 = 10'd350; a_exp2 = 10'd901; a_exp3 = 10'd26;
b_exp0 = 10'd140; b_exp1 = 10'd459; b_exp2 = 10'd219; b_exp3 = 10'd700;
a_sign0 = 4'd14; a_sign1 = 4'd10; a_sign2 = 4'd12; a_sign3 = 4'd11;
b_sign0 = 4'd14; b_sign1 = 4'd12; b_sign2 = 4'd11; b_sign3 = 4'd4;
@(posedge clk_i);
a_mant0 = 8'd250; a_mant1 = 8'd56; a_mant2 = 8'd225; a_mant3 = 8'd116;
b_mant0 = 8'd155; b_mant1 = 8'd104; b_mant2 = 8'd178; b_mant3 = 8'd60;
a_exp0 = 10'd238; a_exp1 = 10'd8; a_exp2 = 10'd555; a_exp3 = 10'd440;
b_exp0 = 10'd859; b_exp1 = 10'd308; b_exp2 = 10'd616; b_exp3 = 10'd987;
a_sign0 = 4'd11; a_sign1 = 4'd3; a_sign2 = 4'd7; a_sign3 = 4'd7;
b_sign0 = 4'd16; b_sign1 = 4'd12; b_sign2 = 4'd13; b_sign3 = 4'd12;
@(posedge clk_i);
a_mant0 = 8'd159; a_mant1 = 8'd111; a_mant2 = 8'd249; a_mant3 = 8'd39;
b_mant0 = 8'd16; b_mant1 = 8'd106; b_mant2 = 8'd216; b_mant3 = 8'd151;
a_exp0 = 10'd712; a_exp1 = 10'd377; a_exp2 = 10'd540; a_exp3 = 10'd184;
b_exp0 = 10'd359; b_exp1 = 10'd431; b_exp2 = 10'd186; b_exp3 = 10'd568;
a_sign0 = 4'd5; a_sign1 = 4'd7; a_sign2 = 4'd2; a_sign3 = 4'd1;
b_sign0 = 4'd4; b_sign1 = 4'd11; b_sign2 = 4'd8; b_sign3 = 4'd12;
@(posedge clk_i);
shared_exps0 = 8'd127;
shared_exps1 = 8'd129;
rstn = 0;
@(posedge clk_i);
rstn = 1;
a_mant0 = 8'd17; a_mant1 = 8'd131; a_mant2 = 8'd169; a_mant3 = 8'd19;
b_mant0 = 8'd61; b_mant1 = 8'd179; b_mant2 = 8'd170; b_mant3 = 8'd115;
a_exp0 = 10'd594; a_exp1 = 10'd260; a_exp2 = 10'd305; a_exp3 = 10'd561;
b_exp0 = 10'd783; b_exp1 = 10'd566; b_exp2 = 10'd170; b_exp3 = 10'd429;
a_sign0 = 4'd6; a_sign1 = 4'd8; a_sign2 = 4'd13; a_sign3 = 4'd1;
b_sign0 = 4'd4; b_sign1 = 4'd10; b_sign2 = 4'd10; b_sign3 = 4'd10;
@(posedge clk_i);
a_mant0 = 8'd68; a_mant1 = 8'd136; a_mant2 = 8'd191; a_mant3 = 8'd26;
b_mant0 = 8'd129; b_mant1 = 8'd224; b_mant2 = 8'd95; b_mant3 = 8'd115;
a_exp0 = 10'd807; a_exp1 = 10'd526; a_exp2 = 10'd674; a_exp3 = 10'd742;
b_exp0 = 10'd104; b_exp1 = 10'd727; b_exp2 = 10'd775; b_exp3 = 10'd347;
a_sign0 = 4'd6; a_sign1 = 4'd5; a_sign2 = 4'd6; a_sign3 = 4'd2;
b_sign0 = 4'd11; b_sign1 = 4'd10; b_sign2 = 4'd8; b_sign3 = 4'd5;
@(posedge clk_i);
a_mant0 = 8'd130; a_mant1 = 8'd190; a_mant2 = 8'd187; a_mant3 = 8'd227;
b_mant0 = 8'd234; b_mant1 = 8'd151; b_mant2 = 8'd111; b_mant3 = 8'd66;
a_exp0 = 10'd546; a_exp1 = 10'd500; a_exp2 = 10'd855; a_exp3 = 10'd707;
b_exp0 = 10'd165; b_exp1 = 10'd325; b_exp2 = 10'd804; b_exp3 = 10'd781;
a_sign0 = 4'd4; a_sign1 = 4'd10; a_sign2 = 4'd15; a_sign3 = 4'd2;
b_sign0 = 4'd9; b_sign1 = 4'd8; b_sign2 = 4'd10; b_sign3 = 4'd11;
@(posedge clk_i);
a_mant0 = 8'd137; a_mant1 = 8'd109; a_mant2 = 8'd129; a_mant3 = 8'd42;
b_mant0 = 8'd10; b_mant1 = 8'd167; b_mant2 = 8'd146; b_mant3 = 8'd51;
a_exp0 = 10'd17; a_exp1 = 10'd248; a_exp2 = 10'd186; a_exp3 = 10'd401;
b_exp0 = 10'd93; b_exp1 = 10'd296; b_exp2 = 10'd436; b_exp3 = 10'd251;
a_sign0 = 4'd11; a_sign1 = 4'd1; a_sign2 = 4'd9; a_sign3 = 4'd8;
b_sign0 = 4'd7; b_sign1 = 4'd10; b_sign2 = 4'd16; b_sign3 = 4'd4;
@(posedge clk_i);
a_mant0 = 8'd3; a_mant1 = 8'd141; a_mant2 = 8'd96; a_mant3 = 8'd183;
b_mant0 = 8'd129; b_mant1 = 8'd229; b_mant2 = 8'd124; b_mant3 = 8'd155;
a_exp0 = 10'd680; a_exp1 = 10'd998; a_exp2 = 10'd211; a_exp3 = 10'd892;
b_exp0 = 10'd579; b_exp1 = 10'd411; b_exp2 = 10'd895; b_exp3 = 10'd23;
a_sign0 = 4'd13; a_sign1 = 4'd15; a_sign2 = 4'd2; a_sign3 = 4'd9;
b_sign0 = 4'd10; b_sign1 = 4'd13; b_sign2 = 4'd7; b_sign3 = 4'd16;
@(posedge clk_i);
a_mant0 = 8'd189; a_mant1 = 8'd32; a_mant2 = 8'd248; a_mant3 = 8'd75;
b_mant0 = 8'd224; b_mant1 = 8'd77; b_mant2 = 8'd182; b_mant3 = 8'd159;
a_exp0 = 10'd875; a_exp1 = 10'd428; a_exp2 = 10'd705; a_exp3 = 10'd684;
b_exp0 = 10'd254; b_exp1 = 10'd741; b_exp2 = 10'd599; b_exp3 = 10'd238;
a_sign0 = 4'd7; a_sign1 = 4'd5; a_sign2 = 4'd5; a_sign3 = 4'd5;
b_sign0 = 4'd0; b_sign1 = 4'd13; b_sign2 = 4'd0; b_sign3 = 4'd5;
@(posedge clk_i);
a_mant0 = 8'd186; a_mant1 = 8'd10; a_mant2 = 8'd181; a_mant3 = 8'd176;
b_mant0 = 8'd97; b_mant1 = 8'd250; b_mant2 = 8'd162; b_mant3 = 8'd88;
a_exp0 = 10'd144; a_exp1 = 10'd1013; a_exp2 = 10'd795; a_exp3 = 10'd966;
b_exp0 = 10'd503; b_exp1 = 10'd1021; b_exp2 = 10'd158; b_exp3 = 10'd454;
a_sign0 = 4'd4; a_sign1 = 4'd8; a_sign2 = 4'd8; a_sign3 = 4'd1;
b_sign0 = 4'd13; b_sign1 = 4'd12; b_sign2 = 4'd7; b_sign3 = 4'd15;
@(posedge clk_i);
shared_exps0 = 8'd106;
shared_exps1 = 8'd132;
a_mant0 = 8'd162; a_mant1 = 8'd140; a_mant2 = 8'd29; a_mant3 = 8'd84;
b_mant0 = 8'd22; b_mant1 = 8'd158; b_mant2 = 8'd201; b_mant3 = 8'd179;
a_exp0 = 10'd144; a_exp1 = 10'd343; a_exp2 = 10'd723; a_exp3 = 10'd416;
b_exp0 = 10'd977; b_exp1 = 10'd579; b_exp2 = 10'd659; b_exp3 = 10'd180;
a_sign0 = 4'd4; a_sign1 = 4'd3; a_sign2 = 4'd3; a_sign3 = 4'd16;
b_sign0 = 4'd14; b_sign1 = 4'd2; b_sign2 = 4'd16; b_sign3 = 4'd3;
@(posedge clk_i);
a_mant0 = 8'd246; a_mant1 = 8'd122; a_mant2 = 8'd62; a_mant3 = 8'd164;
b_mant0 = 8'd86; b_mant1 = 8'd220; b_mant2 = 8'd35; b_mant3 = 8'd205;
a_exp0 = 10'd376; a_exp1 = 10'd47; a_exp2 = 10'd991; a_exp3 = 10'd40;
b_exp0 = 10'd348; b_exp1 = 10'd411; b_exp2 = 10'd210; b_exp3 = 10'd735;
a_sign0 = 4'd15; a_sign1 = 4'd14; a_sign2 = 4'd14; a_sign3 = 4'd13;
b_sign0 = 4'd16; b_sign1 = 4'd2; b_sign2 = 4'd3; b_sign3 = 4'd3;
@(posedge clk_i);
a_mant0 = 8'd15; a_mant1 = 8'd41; a_mant2 = 8'd234; a_mant3 = 8'd38;
b_mant0 = 8'd112; b_mant1 = 8'd164; b_mant2 = 8'd155; b_mant3 = 8'd70;
a_exp0 = 10'd140; a_exp1 = 10'd211; a_exp2 = 10'd845; a_exp3 = 10'd879;
b_exp0 = 10'd235; b_exp1 = 10'd520; b_exp2 = 10'd494; b_exp3 = 10'd703;
a_sign0 = 4'd15; a_sign1 = 4'd4; a_sign2 = 4'd14; a_sign3 = 4'd3;
b_sign0 = 4'd16; b_sign1 = 4'd10; b_sign2 = 4'd14; b_sign3 = 4'd15;
@(posedge clk_i);
a_mant0 = 8'd103; a_mant1 = 8'd244; a_mant2 = 8'd219; a_mant3 = 8'd209;
b_mant0 = 8'd251; b_mant1 = 8'd149; b_mant2 = 8'd51; b_mant3 = 8'd147;
a_exp0 = 10'd367; a_exp1 = 10'd520; a_exp2 = 10'd388; a_exp3 = 10'd169;
b_exp0 = 10'd431; b_exp1 = 10'd420; b_exp2 = 10'd719; b_exp3 = 10'd862;
a_sign0 = 4'd6; a_sign1 = 4'd10; a_sign2 = 4'd6; a_sign3 = 4'd3;
b_sign0 = 4'd9; b_sign1 = 4'd10; b_sign2 = 4'd2; b_sign3 = 4'd12;
@(posedge clk_i);
a_mant0 = 8'd17; a_mant1 = 8'd185; a_mant2 = 8'd54; a_mant3 = 8'd196;
b_mant0 = 8'd215; b_mant1 = 8'd53; b_mant2 = 8'd34; b_mant3 = 8'd146;
a_exp0 = 10'd81; a_exp1 = 10'd522; a_exp2 = 10'd334; a_exp3 = 10'd173;
b_exp0 = 10'd508; b_exp1 = 10'd744; b_exp2 = 10'd716; b_exp3 = 10'd619;
a_sign0 = 4'd14; a_sign1 = 4'd14; a_sign2 = 4'd11; a_sign3 = 4'd13;
b_sign0 = 4'd0; b_sign1 = 4'd15; b_sign2 = 4'd8; b_sign3 = 4'd4;
@(posedge clk_i);
a_mant0 = 8'd38; a_mant1 = 8'd169; a_mant2 = 8'd119; a_mant3 = 8'd51;
b_mant0 = 8'd118; b_mant1 = 8'd75; b_mant2 = 8'd143; b_mant3 = 8'd181;
a_exp0 = 10'd529; a_exp1 = 10'd574; a_exp2 = 10'd347; a_exp3 = 10'd950;
b_exp0 = 10'd667; b_exp1 = 10'd180; b_exp2 = 10'd693; b_exp3 = 10'd366;
a_sign0 = 4'd12; a_sign1 = 4'd5; a_sign2 = 4'd2; a_sign3 = 4'd8;
b_sign0 = 4'd4; b_sign1 = 4'd8; b_sign2 = 4'd6; b_sign3 = 4'd11;
@(posedge clk_i);
a_mant0 = 8'd75; a_mant1 = 8'd232; a_mant2 = 8'd190; a_mant3 = 8'd201;
b_mant0 = 8'd196; b_mant1 = 8'd174; b_mant2 = 8'd225; b_mant3 = 8'd211;
a_exp0 = 10'd935; a_exp1 = 10'd236; a_exp2 = 10'd413; a_exp3 = 10'd877;
b_exp0 = 10'd17; b_exp1 = 10'd464; b_exp2 = 10'd991; b_exp3 = 10'd89;
a_sign0 = 4'd1; a_sign1 = 4'd11; a_sign2 = 4'd3; a_sign3 = 4'd3;
b_sign0 = 4'd10; b_sign1 = 4'd11; b_sign2 = 4'd5; b_sign3 = 4'd14;
@(posedge clk_i);
a_mant0 = 8'd229; a_mant1 = 8'd187; a_mant2 = 8'd30; a_mant3 = 8'd100;
b_mant0 = 8'd30; b_mant1 = 8'd115; b_mant2 = 8'd155; b_mant3 = 8'd215;
a_exp0 = 10'd969; a_exp1 = 10'd877; a_exp2 = 10'd875; a_exp3 = 10'd58;
b_exp0 = 10'd687; b_exp1 = 10'd846; b_exp2 = 10'd623; b_exp3 = 10'd654;
a_sign0 = 4'd10; a_sign1 = 4'd16; a_sign2 = 4'd8; a_sign3 = 4'd1;
b_sign0 = 4'd12; b_sign1 = 4'd9; b_sign2 = 4'd14; b_sign3 = 4'd7;
@(posedge clk_i);
shared_exps0 = 8'd117;
shared_exps1 = 8'd153;
a_mant0 = 8'd205; a_mant1 = 8'd177; a_mant2 = 8'd12; a_mant3 = 8'd162;
b_mant0 = 8'd139; b_mant1 = 8'd138; b_mant2 = 8'd241; b_mant3 = 8'd198;
a_exp0 = 10'd600; a_exp1 = 10'd969; a_exp2 = 10'd818; a_exp3 = 10'd826;
b_exp0 = 10'd153; b_exp1 = 10'd672; b_exp2 = 10'd931; b_exp3 = 10'd159;
a_sign0 = 4'd15; a_sign1 = 4'd13; a_sign2 = 4'd10; a_sign3 = 4'd11;
b_sign0 = 4'd5; b_sign1 = 4'd0; b_sign2 = 4'd14; b_sign3 = 4'd0;
@(posedge clk_i);
a_mant0 = 8'd187; a_mant1 = 8'd51; a_mant2 = 8'd204; a_mant3 = 8'd148;
b_mant0 = 8'd160; b_mant1 = 8'd9; b_mant2 = 8'd62; b_mant3 = 8'd25;
a_exp0 = 10'd509; a_exp1 = 10'd255; a_exp2 = 10'd273; a_exp3 = 10'd917;
b_exp0 = 10'd307; b_exp1 = 10'd787; b_exp2 = 10'd453; b_exp3 = 10'd143;
a_sign0 = 4'd11; a_sign1 = 4'd8; a_sign2 = 4'd6; a_sign3 = 4'd9;
b_sign0 = 4'd14; b_sign1 = 4'd5; b_sign2 = 4'd2; b_sign3 = 4'd9;
@(posedge clk_i);
a_mant0 = 8'd220; a_mant1 = 8'd47; a_mant2 = 8'd246; a_mant3 = 8'd113;
b_mant0 = 8'd187; b_mant1 = 8'd230; b_mant2 = 8'd132; b_mant3 = 8'd48;
a_exp0 = 10'd853; a_exp1 = 10'd798; a_exp2 = 10'd108; a_exp3 = 10'd513;
b_exp0 = 10'd480; b_exp1 = 10'd634; b_exp2 = 10'd212; b_exp3 = 10'd940;
a_sign0 = 4'd4; a_sign1 = 4'd2; a_sign2 = 4'd2; a_sign3 = 4'd15;
b_sign0 = 4'd3; b_sign1 = 4'd5; b_sign2 = 4'd16; b_sign3 = 4'd9;
@(posedge clk_i);
a_mant0 = 8'd43; a_mant1 = 8'd93; a_mant2 = 8'd101; a_mant3 = 8'd214;
b_mant0 = 8'd143; b_mant1 = 8'd242; b_mant2 = 8'd156; b_mant3 = 8'd75;
a_exp0 = 10'd585; a_exp1 = 10'd807; a_exp2 = 10'd943; a_exp3 = 10'd716;
b_exp0 = 10'd361; b_exp1 = 10'd71; b_exp2 = 10'd564; b_exp3 = 10'd88;
a_sign0 = 4'd4; a_sign1 = 4'd15; a_sign2 = 4'd8; a_sign3 = 4'd12;
b_sign0 = 4'd2; b_sign1 = 4'd0; b_sign2 = 4'd8; b_sign3 = 4'd12;
@(posedge clk_i);
a_mant0 = 8'd66; a_mant1 = 8'd111; a_mant2 = 8'd162; a_mant3 = 8'd159;
b_mant0 = 8'd38; b_mant1 = 8'd68; b_mant2 = 8'd118; b_mant3 = 8'd37;
a_exp0 = 10'd654; a_exp1 = 10'd550; a_exp2 = 10'd314; a_exp3 = 10'd3;
b_exp0 = 10'd221; b_exp1 = 10'd769; b_exp2 = 10'd855; b_exp3 = 10'd229;
a_sign0 = 4'd5; a_sign1 = 4'd14; a_sign2 = 4'd4; a_sign3 = 4'd10;
b_sign0 = 4'd3; b_sign1 = 4'd12; b_sign2 = 4'd12; b_sign3 = 4'd15;
@(posedge clk_i);
a_mant0 = 8'd157; a_mant1 = 8'd175; a_mant2 = 8'd103; a_mant3 = 8'd8;
b_mant0 = 8'd169; b_mant1 = 8'd5; b_mant2 = 8'd103; b_mant3 = 8'd39;
a_exp0 = 10'd818; a_exp1 = 10'd122; a_exp2 = 10'd117; a_exp3 = 10'd19;
b_exp0 = 10'd698; b_exp1 = 10'd651; b_exp2 = 10'd431; b_exp3 = 10'd776;
a_sign0 = 4'd14; a_sign1 = 4'd9; a_sign2 = 4'd0; a_sign3 = 4'd15;
b_sign0 = 4'd11; b_sign1 = 4'd14; b_sign2 = 4'd10; b_sign3 = 4'd15;
@(posedge clk_i);
a_mant0 = 8'd50; a_mant1 = 8'd164; a_mant2 = 8'd182; a_mant3 = 8'd162;
b_mant0 = 8'd110; b_mant1 = 8'd191; b_mant2 = 8'd101; b_mant3 = 8'd161;
a_exp0 = 10'd666; a_exp1 = 10'd346; a_exp2 = 10'd489; a_exp3 = 10'd793;
b_exp0 = 10'd857; b_exp1 = 10'd668; b_exp2 = 10'd265; b_exp3 = 10'd96;
a_sign0 = 4'd9; a_sign1 = 4'd15; a_sign2 = 4'd13; a_sign3 = 4'd10;
b_sign0 = 4'd13; b_sign1 = 4'd6; b_sign2 = 4'd7; b_sign3 = 4'd9;
@(posedge clk_i);
a_mant0 = 8'd4; a_mant1 = 8'd75; a_mant2 = 8'd71; a_mant3 = 8'd42;
b_mant0 = 8'd161; b_mant1 = 8'd15; b_mant2 = 8'd107; b_mant3 = 8'd107;
a_exp0 = 10'd238; a_exp1 = 10'd664; a_exp2 = 10'd553; a_exp3 = 10'd981;
b_exp0 = 10'd212; b_exp1 = 10'd335; b_exp2 = 10'd766; b_exp3 = 10'd693;
a_sign0 = 4'd5; a_sign1 = 4'd14; a_sign2 = 4'd10; a_sign3 = 4'd13;
b_sign0 = 4'd11; b_sign1 = 4'd2; b_sign2 = 4'd7; b_sign3 = 4'd3;
@(posedge clk_i);
shared_exps0 = 8'd117;
shared_exps1 = 8'd130;
a_mant0 = 8'd220; a_mant1 = 8'd195; a_mant2 = 8'd70; a_mant3 = 8'd191;
b_mant0 = 8'd93; b_mant1 = 8'd133; b_mant2 = 8'd44; b_mant3 = 8'd142;
a_exp0 = 10'd507; a_exp1 = 10'd327; a_exp2 = 10'd589; a_exp3 = 10'd692;
b_exp0 = 10'd644; b_exp1 = 10'd104; b_exp2 = 10'd1017; b_exp3 = 10'd1009;
a_sign0 = 4'd1; a_sign1 = 4'd13; a_sign2 = 4'd16; a_sign3 = 4'd0;
b_sign0 = 4'd13; b_sign1 = 4'd14; b_sign2 = 4'd1; b_sign3 = 4'd1;
@(posedge clk_i);
a_mant0 = 8'd24; a_mant1 = 8'd192; a_mant2 = 8'd5; a_mant3 = 8'd62;
b_mant0 = 8'd4; b_mant1 = 8'd203; b_mant2 = 8'd50; b_mant3 = 8'd13;
a_exp0 = 10'd996; a_exp1 = 10'd161; a_exp2 = 10'd934; a_exp3 = 10'd590;
b_exp0 = 10'd773; b_exp1 = 10'd437; b_exp2 = 10'd410; b_exp3 = 10'd472;
a_sign0 = 4'd12; a_sign1 = 4'd16; a_sign2 = 4'd10; a_sign3 = 4'd9;
b_sign0 = 4'd12; b_sign1 = 4'd9; b_sign2 = 4'd1; b_sign3 = 4'd4;
@(posedge clk_i);
a_mant0 = 8'd133; a_mant1 = 8'd118; a_mant2 = 8'd154; a_mant3 = 8'd245;
b_mant0 = 8'd0; b_mant1 = 8'd24; b_mant2 = 8'd98; b_mant3 = 8'd32;
a_exp0 = 10'd678; a_exp1 = 10'd753; a_exp2 = 10'd419; a_exp3 = 10'd434;
b_exp0 = 10'd294; b_exp1 = 10'd690; b_exp2 = 10'd211; b_exp3 = 10'd925;
a_sign0 = 4'd15; a_sign1 = 4'd6; a_sign2 = 4'd6; a_sign3 = 4'd4;
b_sign0 = 4'd0; b_sign1 = 4'd2; b_sign2 = 4'd8; b_sign3 = 4'd14;
@(posedge clk_i);
a_mant0 = 8'd163; a_mant1 = 8'd19; a_mant2 = 8'd144; a_mant3 = 8'd178;
b_mant0 = 8'd168; b_mant1 = 8'd171; b_mant2 = 8'd162; b_mant3 = 8'd3;
a_exp0 = 10'd235; a_exp1 = 10'd961; a_exp2 = 10'd399; a_exp3 = 10'd287;
b_exp0 = 10'd296; b_exp1 = 10'd518; b_exp2 = 10'd450; b_exp3 = 10'd470;
a_sign0 = 4'd4; a_sign1 = 4'd4; a_sign2 = 4'd11; a_sign3 = 4'd3;
b_sign0 = 4'd11; b_sign1 = 4'd7; b_sign2 = 4'd8; b_sign3 = 4'd5;
@(posedge clk_i);
a_mant0 = 8'd146; a_mant1 = 8'd92; a_mant2 = 8'd121; a_mant3 = 8'd149;
b_mant0 = 8'd105; b_mant1 = 8'd191; b_mant2 = 8'd109; b_mant3 = 8'd205;
a_exp0 = 10'd81; a_exp1 = 10'd977; a_exp2 = 10'd469; a_exp3 = 10'd267;
b_exp0 = 10'd315; b_exp1 = 10'd653; b_exp2 = 10'd759; b_exp3 = 10'd796;
a_sign0 = 4'd0; a_sign1 = 4'd1; a_sign2 = 4'd1; a_sign3 = 4'd4;
b_sign0 = 4'd10; b_sign1 = 4'd7; b_sign2 = 4'd4; b_sign3 = 4'd4;
@(posedge clk_i);
a_mant0 = 8'd219; a_mant1 = 8'd216; a_mant2 = 8'd118; a_mant3 = 8'd150;
b_mant0 = 8'd170; b_mant1 = 8'd94; b_mant2 = 8'd122; b_mant3 = 8'd104;
a_exp0 = 10'd775; a_exp1 = 10'd354; a_exp2 = 10'd153; a_exp3 = 10'd302;
b_exp0 = 10'd665; b_exp1 = 10'd540; b_exp2 = 10'd813; b_exp3 = 10'd393;
a_sign0 = 4'd12; a_sign1 = 4'd0; a_sign2 = 4'd5; a_sign3 = 4'd0;
b_sign0 = 4'd15; b_sign1 = 4'd15; b_sign2 = 4'd7; b_sign3 = 4'd2;
@(posedge clk_i);
a_mant0 = 8'd107; a_mant1 = 8'd15; a_mant2 = 8'd236; a_mant3 = 8'd240;
b_mant0 = 8'd188; b_mant1 = 8'd202; b_mant2 = 8'd114; b_mant3 = 8'd252;
a_exp0 = 10'd309; a_exp1 = 10'd102; a_exp2 = 10'd413; a_exp3 = 10'd472;
b_exp0 = 10'd969; b_exp1 = 10'd147; b_exp2 = 10'd596; b_exp3 = 10'd1016;
a_sign0 = 4'd6; a_sign1 = 4'd14; a_sign2 = 4'd14; a_sign3 = 4'd13;
b_sign0 = 4'd1; b_sign1 = 4'd4; b_sign2 = 4'd11; b_sign3 = 4'd7;
@(posedge clk_i);
a_mant0 = 8'd95; a_mant1 = 8'd87; a_mant2 = 8'd133; a_mant3 = 8'd17;
b_mant0 = 8'd39; b_mant1 = 8'd74; b_mant2 = 8'd237; b_mant3 = 8'd112;
a_exp0 = 10'd777; a_exp1 = 10'd394; a_exp2 = 10'd442; a_exp3 = 10'd46;
b_exp0 = 10'd678; b_exp1 = 10'd266; b_exp2 = 10'd989; b_exp3 = 10'd776;
a_sign0 = 4'd11; a_sign1 = 4'd6; a_sign2 = 4'd15; a_sign3 = 4'd15;
b_sign0 = 4'd8; b_sign1 = 4'd10; b_sign2 = 4'd1; b_sign3 = 4'd6;
@(posedge clk_i);
shared_exps0 = 8'd119;
shared_exps1 = 8'd111;
rstn = 0;
@(posedge clk_i);
rstn = 1;
a_mant0 = 8'd59; a_mant1 = 8'd222; a_mant2 = 8'd22; a_mant3 = 8'd136;
b_mant0 = 8'd210; b_mant1 = 8'd73; b_mant2 = 8'd17; b_mant3 = 8'd218;
a_exp0 = 10'd802; a_exp1 = 10'd49; a_exp2 = 10'd873; a_exp3 = 10'd433;
b_exp0 = 10'd780; b_exp1 = 10'd751; b_exp2 = 10'd55; b_exp3 = 10'd589;
a_sign0 = 4'd11; a_sign1 = 4'd13; a_sign2 = 4'd12; a_sign3 = 4'd0;
b_sign0 = 4'd1; b_sign1 = 4'd9; b_sign2 = 4'd7; b_sign3 = 4'd12;
@(posedge clk_i);
a_mant0 = 8'd17; a_mant1 = 8'd70; a_mant2 = 8'd224; a_mant3 = 8'd92;
b_mant0 = 8'd115; b_mant1 = 8'd116; b_mant2 = 8'd128; b_mant3 = 8'd183;
a_exp0 = 10'd495; a_exp1 = 10'd949; a_exp2 = 10'd374; a_exp3 = 10'd173;
b_exp0 = 10'd174; b_exp1 = 10'd569; b_exp2 = 10'd955; b_exp3 = 10'd99;
a_sign0 = 4'd13; a_sign1 = 4'd1; a_sign2 = 4'd5; a_sign3 = 4'd6;
b_sign0 = 4'd0; b_sign1 = 4'd3; b_sign2 = 4'd6; b_sign3 = 4'd14;
@(posedge clk_i);
a_mant0 = 8'd237; a_mant1 = 8'd209; a_mant2 = 8'd147; a_mant3 = 8'd37;
b_mant0 = 8'd89; b_mant1 = 8'd197; b_mant2 = 8'd250; b_mant3 = 8'd245;
a_exp0 = 10'd103; a_exp1 = 10'd340; a_exp2 = 10'd354; a_exp3 = 10'd706;
b_exp0 = 10'd588; b_exp1 = 10'd999; b_exp2 = 10'd632; b_exp3 = 10'd167;
a_sign0 = 4'd15; a_sign1 = 4'd3; a_sign2 = 4'd13; a_sign3 = 4'd6;
b_sign0 = 4'd6; b_sign1 = 4'd9; b_sign2 = 4'd2; b_sign3 = 4'd6;
@(posedge clk_i);
a_mant0 = 8'd113; a_mant1 = 8'd214; a_mant2 = 8'd247; a_mant3 = 8'd166;
b_mant0 = 8'd16; b_mant1 = 8'd133; b_mant2 = 8'd77; b_mant3 = 8'd215;
a_exp0 = 10'd822; a_exp1 = 10'd719; a_exp2 = 10'd708; a_exp3 = 10'd41;
b_exp0 = 10'd615; b_exp1 = 10'd270; b_exp2 = 10'd888; b_exp3 = 10'd27;
a_sign0 = 4'd2; a_sign1 = 4'd16; a_sign2 = 4'd15; a_sign3 = 4'd9;
b_sign0 = 4'd15; b_sign1 = 4'd9; b_sign2 = 4'd3; b_sign3 = 4'd5;
@(posedge clk_i);
a_mant0 = 8'd137; a_mant1 = 8'd179; a_mant2 = 8'd175; a_mant3 = 8'd43;
b_mant0 = 8'd24; b_mant1 = 8'd13; b_mant2 = 8'd242; b_mant3 = 8'd165;
a_exp0 = 10'd143; a_exp1 = 10'd41; a_exp2 = 10'd562; a_exp3 = 10'd821;
b_exp0 = 10'd439; b_exp1 = 10'd683; b_exp2 = 10'd530; b_exp3 = 10'd412;
a_sign0 = 4'd10; a_sign1 = 4'd9; a_sign2 = 4'd11; a_sign3 = 4'd10;
b_sign0 = 4'd10; b_sign1 = 4'd9; b_sign2 = 4'd12; b_sign3 = 4'd3;
@(posedge clk_i);
a_mant0 = 8'd6; a_mant1 = 8'd1; a_mant2 = 8'd204; a_mant3 = 8'd242;
b_mant0 = 8'd157; b_mant1 = 8'd233; b_mant2 = 8'd151; b_mant3 = 8'd91;
a_exp0 = 10'd991; a_exp1 = 10'd334; a_exp2 = 10'd799; a_exp3 = 10'd532;
b_exp0 = 10'd337; b_exp1 = 10'd939; b_exp2 = 10'd713; b_exp3 = 10'd750;
a_sign0 = 4'd4; a_sign1 = 4'd1; a_sign2 = 4'd12; a_sign3 = 4'd6;
b_sign0 = 4'd8; b_sign1 = 4'd1; b_sign2 = 4'd9; b_sign3 = 4'd7;
@(posedge clk_i);
a_mant0 = 8'd145; a_mant1 = 8'd46; a_mant2 = 8'd225; a_mant3 = 8'd121;
b_mant0 = 8'd234; b_mant1 = 8'd73; b_mant2 = 8'd234; b_mant3 = 8'd95;
a_exp0 = 10'd291; a_exp1 = 10'd663; a_exp2 = 10'd778; a_exp3 = 10'd464;
b_exp0 = 10'd956; b_exp1 = 10'd945; b_exp2 = 10'd966; b_exp3 = 10'd799;
a_sign0 = 4'd11; a_sign1 = 4'd4; a_sign2 = 4'd11; a_sign3 = 4'd3;
b_sign0 = 4'd8; b_sign1 = 4'd3; b_sign2 = 4'd5; b_sign3 = 4'd5;
@(posedge clk_i);
shared_exps0 = 8'd122;
shared_exps1 = 8'd119;
a_mant0 = 8'd224; a_mant1 = 8'd22; a_mant2 = 8'd112; a_mant3 = 8'd55;
b_mant0 = 8'd155; b_mant1 = 8'd239; b_mant2 = 8'd238; b_mant3 = 8'd116;
a_exp0 = 10'd775; a_exp1 = 10'd585; a_exp2 = 10'd973; a_exp3 = 10'd475;
b_exp0 = 10'd363; b_exp1 = 10'd638; b_exp2 = 10'd356; b_exp3 = 10'd987;
a_sign0 = 4'd4; a_sign1 = 4'd12; a_sign2 = 4'd13; a_sign3 = 4'd9;
b_sign0 = 4'd6; b_sign1 = 4'd6; b_sign2 = 4'd15; b_sign3 = 4'd1;
@(posedge clk_i);
a_mant0 = 8'd195; a_mant1 = 8'd209; a_mant2 = 8'd44; a_mant3 = 8'd57;
b_mant0 = 8'd83; b_mant1 = 8'd50; b_mant2 = 8'd170; b_mant3 = 8'd207;
a_exp0 = 10'd30; a_exp1 = 10'd637; a_exp2 = 10'd305; a_exp3 = 10'd614;
b_exp0 = 10'd428; b_exp1 = 10'd986; b_exp2 = 10'd542; b_exp3 = 10'd525;
a_sign0 = 4'd0; a_sign1 = 4'd2; a_sign2 = 4'd8; a_sign3 = 4'd6;
b_sign0 = 4'd5; b_sign1 = 4'd11; b_sign2 = 4'd14; b_sign3 = 4'd3;
@(posedge clk_i);
a_mant0 = 8'd127; a_mant1 = 8'd82; a_mant2 = 8'd46; a_mant3 = 8'd152;
b_mant0 = 8'd54; b_mant1 = 8'd118; b_mant2 = 8'd45; b_mant3 = 8'd131;
a_exp0 = 10'd541; a_exp1 = 10'd66; a_exp2 = 10'd977; a_exp3 = 10'd897;
b_exp0 = 10'd529; b_exp1 = 10'd458; b_exp2 = 10'd18; b_exp3 = 10'd596;
a_sign0 = 4'd3; a_sign1 = 4'd1; a_sign2 = 4'd7; a_sign3 = 4'd6;
b_sign0 = 4'd9; b_sign1 = 4'd8; b_sign2 = 4'd13; b_sign3 = 4'd3;
@(posedge clk_i);
a_mant0 = 8'd210; a_mant1 = 8'd243; a_mant2 = 8'd245; a_mant3 = 8'd98;
b_mant0 = 8'd15; b_mant1 = 8'd185; b_mant2 = 8'd252; b_mant3 = 8'd138;
a_exp0 = 10'd341; a_exp1 = 10'd69; a_exp2 = 10'd141; a_exp3 = 10'd810;
b_exp0 = 10'd412; b_exp1 = 10'd128; b_exp2 = 10'd622; b_exp3 = 10'd622;
a_sign0 = 4'd12; a_sign1 = 4'd7; a_sign2 = 4'd3; a_sign3 = 4'd1;
b_sign0 = 4'd0; b_sign1 = 4'd8; b_sign2 = 4'd12; b_sign3 = 4'd2;
@(posedge clk_i);
a_mant0 = 8'd173; a_mant1 = 8'd140; a_mant2 = 8'd192; a_mant3 = 8'd252;
b_mant0 = 8'd68; b_mant1 = 8'd93; b_mant2 = 8'd155; b_mant3 = 8'd192;
a_exp0 = 10'd0; a_exp1 = 10'd971; a_exp2 = 10'd848; a_exp3 = 10'd569;
b_exp0 = 10'd958; b_exp1 = 10'd988; b_exp2 = 10'd698; b_exp3 = 10'd194;
a_sign0 = 4'd7; a_sign1 = 4'd8; a_sign2 = 4'd1; a_sign3 = 4'd15;
b_sign0 = 4'd3; b_sign1 = 4'd6; b_sign2 = 4'd5; b_sign3 = 4'd2;
@(posedge clk_i);
a_mant0 = 8'd184; a_mant1 = 8'd142; a_mant2 = 8'd153; a_mant3 = 8'd44;
b_mant0 = 8'd126; b_mant1 = 8'd85; b_mant2 = 8'd67; b_mant3 = 8'd156;
a_exp0 = 10'd892; a_exp1 = 10'd187; a_exp2 = 10'd1005; a_exp3 = 10'd206;
b_exp0 = 10'd137; b_exp1 = 10'd786; b_exp2 = 10'd504; b_exp3 = 10'd711;
a_sign0 = 4'd4; a_sign1 = 4'd12; a_sign2 = 4'd6; a_sign3 = 4'd0;
b_sign0 = 4'd6; b_sign1 = 4'd12; b_sign2 = 4'd15; b_sign3 = 4'd4;
@(posedge clk_i);
a_mant0 = 8'd132; a_mant1 = 8'd226; a_mant2 = 8'd204; a_mant3 = 8'd99;
b_mant0 = 8'd29; b_mant1 = 8'd170; b_mant2 = 8'd85; b_mant3 = 8'd102;
a_exp0 = 10'd301; a_exp1 = 10'd582; a_exp2 = 10'd185; a_exp3 = 10'd902;
b_exp0 = 10'd950; b_exp1 = 10'd321; b_exp2 = 10'd288; b_exp3 = 10'd264;
a_sign0 = 4'd15; a_sign1 = 4'd9; a_sign2 = 4'd14; a_sign3 = 4'd9;
b_sign0 = 4'd0; b_sign1 = 4'd0; b_sign2 = 4'd3; b_sign3 = 4'd2;
@(posedge clk_i);
a_mant0 = 8'd29; a_mant1 = 8'd115; a_mant2 = 8'd183; a_mant3 = 8'd122;
b_mant0 = 8'd149; b_mant1 = 8'd20; b_mant2 = 8'd247; b_mant3 = 8'd160;
a_exp0 = 10'd699; a_exp1 = 10'd413; a_exp2 = 10'd261; a_exp3 = 10'd173;
b_exp0 = 10'd108; b_exp1 = 10'd287; b_exp2 = 10'd935; b_exp3 = 10'd456;
a_sign0 = 4'd8; a_sign1 = 4'd4; a_sign2 = 4'd13; a_sign3 = 4'd12;
b_sign0 = 4'd14; b_sign1 = 4'd2; b_sign2 = 4'd7; b_sign3 = 4'd2;
@(posedge clk_i);
shared_exps0 = 8'd153;
shared_exps1 = 8'd128;
a_mant0 = 8'd222; a_mant1 = 8'd71; a_mant2 = 8'd4; a_mant3 = 8'd230;
b_mant0 = 8'd195; b_mant1 = 8'd77; b_mant2 = 8'd49; b_mant3 = 8'd253;
a_exp0 = 10'd124; a_exp1 = 10'd729; a_exp2 = 10'd231; a_exp3 = 10'd925;
b_exp0 = 10'd641; b_exp1 = 10'd42; b_exp2 = 10'd927; b_exp3 = 10'd576;
a_sign0 = 4'd0; a_sign1 = 4'd3; a_sign2 = 4'd0; a_sign3 = 4'd14;
b_sign0 = 4'd2; b_sign1 = 4'd6; b_sign2 = 4'd0; b_sign3 = 4'd8;
@(posedge clk_i);
a_mant0 = 8'd5; a_mant1 = 8'd45; a_mant2 = 8'd188; a_mant3 = 8'd31;
b_mant0 = 8'd198; b_mant1 = 8'd252; b_mant2 = 8'd165; b_mant3 = 8'd145;
a_exp0 = 10'd239; a_exp1 = 10'd783; a_exp2 = 10'd302; a_exp3 = 10'd1003;
b_exp0 = 10'd361; b_exp1 = 10'd557; b_exp2 = 10'd38; b_exp3 = 10'd121;
a_sign0 = 4'd16; a_sign1 = 4'd9; a_sign2 = 4'd14; a_sign3 = 4'd6;
b_sign0 = 4'd8; b_sign1 = 4'd13; b_sign2 = 4'd9; b_sign3 = 4'd0;
@(posedge clk_i);
a_mant0 = 8'd105; a_mant1 = 8'd4; a_mant2 = 8'd177; a_mant3 = 8'd166;
b_mant0 = 8'd221; b_mant1 = 8'd177; b_mant2 = 8'd182; b_mant3 = 8'd210;
a_exp0 = 10'd632; a_exp1 = 10'd508; a_exp2 = 10'd366; a_exp3 = 10'd256;
b_exp0 = 10'd397; b_exp1 = 10'd248; b_exp2 = 10'd651; b_exp3 = 10'd376;
a_sign0 = 4'd9; a_sign1 = 4'd16; a_sign2 = 4'd16; a_sign3 = 4'd13;
b_sign0 = 4'd16; b_sign1 = 4'd14; b_sign2 = 4'd11; b_sign3 = 4'd4;
@(posedge clk_i);
a_mant0 = 8'd32; a_mant1 = 8'd213; a_mant2 = 8'd1; a_mant3 = 8'd170;
b_mant0 = 8'd210; b_mant1 = 8'd121; b_mant2 = 8'd166; b_mant3 = 8'd137;
a_exp0 = 10'd974; a_exp1 = 10'd21; a_exp2 = 10'd941; a_exp3 = 10'd752;
b_exp0 = 10'd676; b_exp1 = 10'd307; b_exp2 = 10'd802; b_exp3 = 10'd235;
a_sign0 = 4'd2; a_sign1 = 4'd9; a_sign2 = 4'd14; a_sign3 = 4'd11;
b_sign0 = 4'd7; b_sign1 = 4'd5; b_sign2 = 4'd1; b_sign3 = 4'd8;
@(posedge clk_i);
a_mant0 = 8'd66; a_mant1 = 8'd68; a_mant2 = 8'd215; a_mant3 = 8'd93;
b_mant0 = 8'd33; b_mant1 = 8'd28; b_mant2 = 8'd102; b_mant3 = 8'd7;
a_exp0 = 10'd242; a_exp1 = 10'd60; a_exp2 = 10'd458; a_exp3 = 10'd282;
b_exp0 = 10'd904; b_exp1 = 10'd738; b_exp2 = 10'd746; b_exp3 = 10'd963;
a_sign0 = 4'd15; a_sign1 = 4'd14; a_sign2 = 4'd10; a_sign3 = 4'd4;
b_sign0 = 4'd16; b_sign1 = 4'd12; b_sign2 = 4'd0; b_sign3 = 4'd11;
@(posedge clk_i);
a_mant0 = 8'd203; a_mant1 = 8'd160; a_mant2 = 8'd164; a_mant3 = 8'd144;
b_mant0 = 8'd112; b_mant1 = 8'd42; b_mant2 = 8'd63; b_mant3 = 8'd160;
a_exp0 = 10'd595; a_exp1 = 10'd156; a_exp2 = 10'd416; a_exp3 = 10'd215;
b_exp0 = 10'd199; b_exp1 = 10'd402; b_exp2 = 10'd887; b_exp3 = 10'd350;
a_sign0 = 4'd11; a_sign1 = 4'd14; a_sign2 = 4'd3; a_sign3 = 4'd1;
b_sign0 = 4'd16; b_sign1 = 4'd3; b_sign2 = 4'd13; b_sign3 = 4'd5;
@(posedge clk_i);
a_mant0 = 8'd121; a_mant1 = 8'd79; a_mant2 = 8'd203; a_mant3 = 8'd4;
b_mant0 = 8'd101; b_mant1 = 8'd36; b_mant2 = 8'd254; b_mant3 = 8'd254;
a_exp0 = 10'd861; a_exp1 = 10'd777; a_exp2 = 10'd299; a_exp3 = 10'd279;
b_exp0 = 10'd994; b_exp1 = 10'd290; b_exp2 = 10'd646; b_exp3 = 10'd388;
a_sign0 = 4'd5; a_sign1 = 4'd1; a_sign2 = 4'd16; a_sign3 = 4'd14;
b_sign0 = 4'd1; b_sign1 = 4'd1; b_sign2 = 4'd9; b_sign3 = 4'd5;
@(posedge clk_i);
a_mant0 = 8'd7; a_mant1 = 8'd115; a_mant2 = 8'd103; a_mant3 = 8'd253;
b_mant0 = 8'd73; b_mant1 = 8'd36; b_mant2 = 8'd89; b_mant3 = 8'd70;
a_exp0 = 10'd933; a_exp1 = 10'd818; a_exp2 = 10'd219; a_exp3 = 10'd267;
b_exp0 = 10'd740; b_exp1 = 10'd939; b_exp2 = 10'd708; b_exp3 = 10'd574;
a_sign0 = 4'd4; a_sign1 = 4'd9; a_sign2 = 4'd3; a_sign3 = 4'd13;
b_sign0 = 4'd6; b_sign1 = 4'd2; b_sign2 = 4'd8; b_sign3 = 4'd16;
@(posedge clk_i);
shared_exps0 = 8'd133;
shared_exps1 = 8'd146;
a_mant0 = 8'd145; a_mant1 = 8'd123; a_mant2 = 8'd174; a_mant3 = 8'd10;
b_mant0 = 8'd4; b_mant1 = 8'd198; b_mant2 = 8'd129; b_mant3 = 8'd90;
a_exp0 = 10'd345; a_exp1 = 10'd456; a_exp2 = 10'd575; a_exp3 = 10'd65;
b_exp0 = 10'd146; b_exp1 = 10'd319; b_exp2 = 10'd580; b_exp3 = 10'd354;
a_sign0 = 4'd10; a_sign1 = 4'd5; a_sign2 = 4'd7; a_sign3 = 4'd8;
b_sign0 = 4'd8; b_sign1 = 4'd3; b_sign2 = 4'd8; b_sign3 = 4'd11;
@(posedge clk_i);
a_mant0 = 8'd132; a_mant1 = 8'd45; a_mant2 = 8'd35; a_mant3 = 8'd224;
b_mant0 = 8'd83; b_mant1 = 8'd194; b_mant2 = 8'd118; b_mant3 = 8'd88;
a_exp0 = 10'd658; a_exp1 = 10'd214; a_exp2 = 10'd91; a_exp3 = 10'd672;
b_exp0 = 10'd482; b_exp1 = 10'd444; b_exp2 = 10'd619; b_exp3 = 10'd641;
a_sign0 = 4'd2; a_sign1 = 4'd10; a_sign2 = 4'd4; a_sign3 = 4'd6;
b_sign0 = 4'd12; b_sign1 = 4'd14; b_sign2 = 4'd5; b_sign3 = 4'd16;
@(posedge clk_i);
a_mant0 = 8'd140; a_mant1 = 8'd217; a_mant2 = 8'd225; a_mant3 = 8'd35;
b_mant0 = 8'd149; b_mant1 = 8'd98; b_mant2 = 8'd204; b_mant3 = 8'd68;
a_exp0 = 10'd419; a_exp1 = 10'd893; a_exp2 = 10'd825; a_exp3 = 10'd723;
b_exp0 = 10'd433; b_exp1 = 10'd711; b_exp2 = 10'd208; b_exp3 = 10'd622;
a_sign0 = 4'd15; a_sign1 = 4'd3; a_sign2 = 4'd7; a_sign3 = 4'd15;
b_sign0 = 4'd8; b_sign1 = 4'd2; b_sign2 = 4'd8; b_sign3 = 4'd7;
@(posedge clk_i);
a_mant0 = 8'd104; a_mant1 = 8'd253; a_mant2 = 8'd45; a_mant3 = 8'd242;
b_mant0 = 8'd19; b_mant1 = 8'd180; b_mant2 = 8'd132; b_mant3 = 8'd234;
a_exp0 = 10'd481; a_exp1 = 10'd809; a_exp2 = 10'd283; a_exp3 = 10'd404;
b_exp0 = 10'd389; b_exp1 = 10'd52; b_exp2 = 10'd439; b_exp3 = 10'd419;
a_sign0 = 4'd2; a_sign1 = 4'd11; a_sign2 = 4'd6; a_sign3 = 4'd4;
b_sign0 = 4'd2; b_sign1 = 4'd11; b_sign2 = 4'd6; b_sign3 = 4'd5;
@(posedge clk_i);
a_mant0 = 8'd195; a_mant1 = 8'd75; a_mant2 = 8'd156; a_mant3 = 8'd119;
b_mant0 = 8'd83; b_mant1 = 8'd84; b_mant2 = 8'd50; b_mant3 = 8'd87;
a_exp0 = 10'd733; a_exp1 = 10'd430; a_exp2 = 10'd536; a_exp3 = 10'd841;
b_exp0 = 10'd220; b_exp1 = 10'd210; b_exp2 = 10'd717; b_exp3 = 10'd973;
a_sign0 = 4'd2; a_sign1 = 4'd0; a_sign2 = 4'd9; a_sign3 = 4'd2;
b_sign0 = 4'd1; b_sign1 = 4'd14; b_sign2 = 4'd0; b_sign3 = 4'd10;
@(posedge clk_i);
a_mant0 = 8'd164; a_mant1 = 8'd196; a_mant2 = 8'd105; a_mant3 = 8'd42;
b_mant0 = 8'd143; b_mant1 = 8'd248; b_mant2 = 8'd81; b_mant3 = 8'd197;
a_exp0 = 10'd800; a_exp1 = 10'd117; a_exp2 = 10'd67; a_exp3 = 10'd387;
b_exp0 = 10'd38; b_exp1 = 10'd77; b_exp2 = 10'd859; b_exp3 = 10'd667;
a_sign0 = 4'd2; a_sign1 = 4'd8; a_sign2 = 4'd0; a_sign3 = 4'd10;
b_sign0 = 4'd11; b_sign1 = 4'd5; b_sign2 = 4'd8; b_sign3 = 4'd11;
@(posedge clk_i);
a_mant0 = 8'd15; a_mant1 = 8'd12; a_mant2 = 8'd195; a_mant3 = 8'd0;
b_mant0 = 8'd190; b_mant1 = 8'd248; b_mant2 = 8'd160; b_mant3 = 8'd68;
a_exp0 = 10'd480; a_exp1 = 10'd595; a_exp2 = 10'd492; a_exp3 = 10'd753;
b_exp0 = 10'd287; b_exp1 = 10'd102; b_exp2 = 10'd852; b_exp3 = 10'd651;
a_sign0 = 4'd16; a_sign1 = 4'd6; a_sign2 = 4'd12; a_sign3 = 4'd3;
b_sign0 = 4'd16; b_sign1 = 4'd9; b_sign2 = 4'd7; b_sign3 = 4'd16;
@(posedge clk_i);
a_mant0 = 8'd237; a_mant1 = 8'd252; a_mant2 = 8'd222; a_mant3 = 8'd0;
b_mant0 = 8'd202; b_mant1 = 8'd185; b_mant2 = 8'd121; b_mant3 = 8'd156;
a_exp0 = 10'd208; a_exp1 = 10'd714; a_exp2 = 10'd400; a_exp3 = 10'd941;
b_exp0 = 10'd195; b_exp1 = 10'd901; b_exp2 = 10'd583; b_exp3 = 10'd553;
a_sign0 = 4'd1; a_sign1 = 4'd0; a_sign2 = 4'd7; a_sign3 = 4'd0;
b_sign0 = 4'd14; b_sign1 = 4'd12; b_sign2 = 4'd16; b_sign3 = 4'd13;
@(posedge clk_i);
shared_exps0 = 8'd131;
shared_exps1 = 8'd127;
rstn = 0;
@(posedge clk_i);
rstn = 1;
a_mant0 = 8'd173; a_mant1 = 8'd210; a_mant2 = 8'd183; a_mant3 = 8'd15;
b_mant0 = 8'd112; b_mant1 = 8'd35; b_mant2 = 8'd227; b_mant3 = 8'd145;
a_exp0 = 10'd209; a_exp1 = 10'd822; a_exp2 = 10'd416; a_exp3 = 10'd279;
b_exp0 = 10'd28; b_exp1 = 10'd132; b_exp2 = 10'd657; b_exp3 = 10'd383;
a_sign0 = 4'd11; a_sign1 = 4'd14; a_sign2 = 4'd15; a_sign3 = 4'd9;
b_sign0 = 4'd14; b_sign1 = 4'd16; b_sign2 = 4'd8; b_sign3 = 4'd5;
@(posedge clk_i);
a_mant0 = 8'd134; a_mant1 = 8'd70; a_mant2 = 8'd45; a_mant3 = 8'd200;
b_mant0 = 8'd118; b_mant1 = 8'd240; b_mant2 = 8'd244; b_mant3 = 8'd223;
a_exp0 = 10'd653; a_exp1 = 10'd972; a_exp2 = 10'd746; a_exp3 = 10'd995;
b_exp0 = 10'd119; b_exp1 = 10'd837; b_exp2 = 10'd744; b_exp3 = 10'd578;
a_sign0 = 4'd12; a_sign1 = 4'd6; a_sign2 = 4'd2; a_sign3 = 4'd16;
b_sign0 = 4'd6; b_sign1 = 4'd12; b_sign2 = 4'd6; b_sign3 = 4'd10;
@(posedge clk_i);
a_mant0 = 8'd103; a_mant1 = 8'd243; a_mant2 = 8'd158; a_mant3 = 8'd100;
b_mant0 = 8'd127; b_mant1 = 8'd28; b_mant2 = 8'd14; b_mant3 = 8'd62;
a_exp0 = 10'd198; a_exp1 = 10'd51; a_exp2 = 10'd449; a_exp3 = 10'd1004;
b_exp0 = 10'd468; b_exp1 = 10'd246; b_exp2 = 10'd665; b_exp3 = 10'd665;
a_sign0 = 4'd6; a_sign1 = 4'd10; a_sign2 = 4'd9; a_sign3 = 4'd8;
b_sign0 = 4'd0; b_sign1 = 4'd3; b_sign2 = 4'd14; b_sign3 = 4'd3;
@(posedge clk_i);
a_mant0 = 8'd48; a_mant1 = 8'd59; a_mant2 = 8'd165; a_mant3 = 8'd10;
b_mant0 = 8'd146; b_mant1 = 8'd219; b_mant2 = 8'd159; b_mant3 = 8'd101;
a_exp0 = 10'd1006; a_exp1 = 10'd86; a_exp2 = 10'd172; a_exp3 = 10'd249;
b_exp0 = 10'd564; b_exp1 = 10'd563; b_exp2 = 10'd320; b_exp3 = 10'd488;
a_sign0 = 4'd14; a_sign1 = 4'd9; a_sign2 = 4'd16; a_sign3 = 4'd1;
b_sign0 = 4'd9; b_sign1 = 4'd16; b_sign2 = 4'd2; b_sign3 = 4'd15;
@(posedge clk_i);
a_mant0 = 8'd82; a_mant1 = 8'd71; a_mant2 = 8'd84; a_mant3 = 8'd64;
b_mant0 = 8'd219; b_mant1 = 8'd152; b_mant2 = 8'd224; b_mant3 = 8'd190;
a_exp0 = 10'd110; a_exp1 = 10'd714; a_exp2 = 10'd201; a_exp3 = 10'd618;
b_exp0 = 10'd234; b_exp1 = 10'd491; b_exp2 = 10'd394; b_exp3 = 10'd441;
a_sign0 = 4'd2; a_sign1 = 4'd0; a_sign2 = 4'd11; a_sign3 = 4'd6;
b_sign0 = 4'd13; b_sign1 = 4'd10; b_sign2 = 4'd8; b_sign3 = 4'd15;
@(posedge clk_i);
a_mant0 = 8'd143; a_mant1 = 8'd183; a_mant2 = 8'd209; a_mant3 = 8'd81;
b_mant0 = 8'd103; b_mant1 = 8'd31; b_mant2 = 8'd55; b_mant3 = 8'd87;
a_exp0 = 10'd947; a_exp1 = 10'd893; a_exp2 = 10'd166; a_exp3 = 10'd406;
b_exp0 = 10'd55; b_exp1 = 10'd105; b_exp2 = 10'd329; b_exp3 = 10'd707;
a_sign0 = 4'd8; a_sign1 = 4'd2; a_sign2 = 4'd0; a_sign3 = 4'd13;
b_sign0 = 4'd16; b_sign1 = 4'd13; b_sign2 = 4'd2; b_sign3 = 4'd4;
@(posedge clk_i);
a_mant0 = 8'd73; a_mant1 = 8'd218; a_mant2 = 8'd10; a_mant3 = 8'd242;
b_mant0 = 8'd255; b_mant1 = 8'd58; b_mant2 = 8'd137; b_mant3 = 8'd0;
a_exp0 = 10'd843; a_exp1 = 10'd80; a_exp2 = 10'd161; a_exp3 = 10'd844;
b_exp0 = 10'd807; b_exp1 = 10'd821; b_exp2 = 10'd251; b_exp3 = 10'd505;
a_sign0 = 4'd4; a_sign1 = 4'd5; a_sign2 = 4'd7; a_sign3 = 4'd6;
b_sign0 = 4'd7; b_sign1 = 4'd7; b_sign2 = 4'd5; b_sign3 = 4'd4;
@(posedge clk_i);
shared_exps0 = 8'd128;
shared_exps1 = 8'd127;
a_mant0 = 8'd142; a_mant1 = 8'd8; a_mant2 = 8'd142; a_mant3 = 8'd105;
b_mant0 = 8'd254; b_mant1 = 8'd46; b_mant2 = 8'd106; b_mant3 = 8'd104;
a_exp0 = 10'd295; a_exp1 = 10'd169; a_exp2 = 10'd683; a_exp3 = 10'd60;
b_exp0 = 10'd201; b_exp1 = 10'd780; b_exp2 = 10'd117; b_exp3 = 10'd770;
a_sign0 = 4'd1; a_sign1 = 4'd5; a_sign2 = 4'd13; a_sign3 = 4'd0;
b_sign0 = 4'd4; b_sign1 = 4'd13; b_sign2 = 4'd3; b_sign3 = 4'd4;
@(posedge clk_i);
a_mant0 = 8'd226; a_mant1 = 8'd103; a_mant2 = 8'd155; a_mant3 = 8'd135;
b_mant0 = 8'd115; b_mant1 = 8'd98; b_mant2 = 8'd4; b_mant3 = 8'd19;
a_exp0 = 10'd357; a_exp1 = 10'd603; a_exp2 = 10'd997; a_exp3 = 10'd451;
b_exp0 = 10'd543; b_exp1 = 10'd338; b_exp2 = 10'd601; b_exp3 = 10'd597;
a_sign0 = 4'd9; a_sign1 = 4'd10; a_sign2 = 4'd2; a_sign3 = 4'd0;
b_sign0 = 4'd13; b_sign1 = 4'd8; b_sign2 = 4'd15; b_sign3 = 4'd1;
@(posedge clk_i);
a_mant0 = 8'd186; a_mant1 = 8'd55; a_mant2 = 8'd108; a_mant3 = 8'd69;
b_mant0 = 8'd165; b_mant1 = 8'd166; b_mant2 = 8'd234; b_mant3 = 8'd97;
a_exp0 = 10'd560; a_exp1 = 10'd863; a_exp2 = 10'd457; a_exp3 = 10'd908;
b_exp0 = 10'd57; b_exp1 = 10'd120; b_exp2 = 10'd219; b_exp3 = 10'd191;
a_sign0 = 4'd5; a_sign1 = 4'd0; a_sign2 = 4'd2; a_sign3 = 4'd7;
b_sign0 = 4'd0; b_sign1 = 4'd3; b_sign2 = 4'd12; b_sign3 = 4'd2;
@(posedge clk_i);
a_mant0 = 8'd88; a_mant1 = 8'd105; a_mant2 = 8'd177; a_mant3 = 8'd237;
b_mant0 = 8'd90; b_mant1 = 8'd177; b_mant2 = 8'd225; b_mant3 = 8'd45;
a_exp0 = 10'd947; a_exp1 = 10'd349; a_exp2 = 10'd686; a_exp3 = 10'd895;
b_exp0 = 10'd430; b_exp1 = 10'd257; b_exp2 = 10'd352; b_exp3 = 10'd121;
a_sign0 = 4'd2; a_sign1 = 4'd9; a_sign2 = 4'd2; a_sign3 = 4'd2;
b_sign0 = 4'd10; b_sign1 = 4'd6; b_sign2 = 4'd4; b_sign3 = 4'd1;
@(posedge clk_i);
a_mant0 = 8'd239; a_mant1 = 8'd35; a_mant2 = 8'd224; a_mant3 = 8'd155;
b_mant0 = 8'd154; b_mant1 = 8'd110; b_mant2 = 8'd152; b_mant3 = 8'd219;
a_exp0 = 10'd799; a_exp1 = 10'd13; a_exp2 = 10'd216; a_exp3 = 10'd628;
b_exp0 = 10'd549; b_exp1 = 10'd207; b_exp2 = 10'd278; b_exp3 = 10'd863;
a_sign0 = 4'd16; a_sign1 = 4'd1; a_sign2 = 4'd2; a_sign3 = 4'd13;
b_sign0 = 4'd11; b_sign1 = 4'd9; b_sign2 = 4'd14; b_sign3 = 4'd2;
@(posedge clk_i);
a_mant0 = 8'd76; a_mant1 = 8'd228; a_mant2 = 8'd127; a_mant3 = 8'd213;
b_mant0 = 8'd1; b_mant1 = 8'd226; b_mant2 = 8'd20; b_mant3 = 8'd150;
a_exp0 = 10'd275; a_exp1 = 10'd675; a_exp2 = 10'd200; a_exp3 = 10'd160;
b_exp0 = 10'd809; b_exp1 = 10'd482; b_exp2 = 10'd256; b_exp3 = 10'd709;
a_sign0 = 4'd3; a_sign1 = 4'd4; a_sign2 = 4'd9; a_sign3 = 4'd9;
b_sign0 = 4'd13; b_sign1 = 4'd14; b_sign2 = 4'd15; b_sign3 = 4'd11;
@(posedge clk_i);
a_mant0 = 8'd131; a_mant1 = 8'd18; a_mant2 = 8'd31; a_mant3 = 8'd154;
b_mant0 = 8'd32; b_mant1 = 8'd207; b_mant2 = 8'd177; b_mant3 = 8'd229;
a_exp0 = 10'd824; a_exp1 = 10'd599; a_exp2 = 10'd914; a_exp3 = 10'd726;
b_exp0 = 10'd107; b_exp1 = 10'd564; b_exp2 = 10'd470; b_exp3 = 10'd54;
a_sign0 = 4'd12; a_sign1 = 4'd16; a_sign2 = 4'd1; a_sign3 = 4'd2;
b_sign0 = 4'd2; b_sign1 = 4'd4; b_sign2 = 4'd9; b_sign3 = 4'd2;
@(posedge clk_i);
a_mant0 = 8'd158; a_mant1 = 8'd1; a_mant2 = 8'd22; a_mant3 = 8'd162;
b_mant0 = 8'd58; b_mant1 = 8'd124; b_mant2 = 8'd183; b_mant3 = 8'd101;
a_exp0 = 10'd329; a_exp1 = 10'd883; a_exp2 = 10'd997; a_exp3 = 10'd130;
b_exp0 = 10'd723; b_exp1 = 10'd345; b_exp2 = 10'd668; b_exp3 = 10'd508;
a_sign0 = 4'd0; a_sign1 = 4'd2; a_sign2 = 4'd16; a_sign3 = 4'd14;
b_sign0 = 4'd15; b_sign1 = 4'd11; b_sign2 = 4'd6; b_sign3 = 4'd6;
@(posedge clk_i);
shared_exps0 = 8'd113;
shared_exps1 = 8'd131;
a_mant0 = 8'd69; a_mant1 = 8'd163; a_mant2 = 8'd155; a_mant3 = 8'd50;
b_mant0 = 8'd162; b_mant1 = 8'd201; b_mant2 = 8'd66; b_mant3 = 8'd34;
a_exp0 = 10'd5; a_exp1 = 10'd524; a_exp2 = 10'd459; a_exp3 = 10'd716;
b_exp0 = 10'd982; b_exp1 = 10'd135; b_exp2 = 10'd627; b_exp3 = 10'd560;
a_sign0 = 4'd4; a_sign1 = 4'd4; a_sign2 = 4'd7; a_sign3 = 4'd10;
b_sign0 = 4'd9; b_sign1 = 4'd13; b_sign2 = 4'd0; b_sign3 = 4'd16;
@(posedge clk_i);
a_mant0 = 8'd17; a_mant1 = 8'd223; a_mant2 = 8'd219; a_mant3 = 8'd96;
b_mant0 = 8'd190; b_mant1 = 8'd19; b_mant2 = 8'd17; b_mant3 = 8'd237;
a_exp0 = 10'd928; a_exp1 = 10'd360; a_exp2 = 10'd611; a_exp3 = 10'd127;
b_exp0 = 10'd233; b_exp1 = 10'd547; b_exp2 = 10'd580; b_exp3 = 10'd363;
a_sign0 = 4'd10; a_sign1 = 4'd11; a_sign2 = 4'd1; a_sign3 = 4'd9;
b_sign0 = 4'd15; b_sign1 = 4'd2; b_sign2 = 4'd12; b_sign3 = 4'd15;
@(posedge clk_i);
a_mant0 = 8'd115; a_mant1 = 8'd173; a_mant2 = 8'd115; a_mant3 = 8'd71;
b_mant0 = 8'd236; b_mant1 = 8'd63; b_mant2 = 8'd241; b_mant3 = 8'd170;
a_exp0 = 10'd296; a_exp1 = 10'd249; a_exp2 = 10'd572; a_exp3 = 10'd318;
b_exp0 = 10'd125; b_exp1 = 10'd830; b_exp2 = 10'd557; b_exp3 = 10'd597;
a_sign0 = 4'd3; a_sign1 = 4'd9; a_sign2 = 4'd0; a_sign3 = 4'd14;
b_sign0 = 4'd2; b_sign1 = 4'd3; b_sign2 = 4'd0; b_sign3 = 4'd5;
@(posedge clk_i);
a_mant0 = 8'd109; a_mant1 = 8'd74; a_mant2 = 8'd3; a_mant3 = 8'd44;
b_mant0 = 8'd28; b_mant1 = 8'd214; b_mant2 = 8'd212; b_mant3 = 8'd166;
a_exp0 = 10'd728; a_exp1 = 10'd724; a_exp2 = 10'd215; a_exp3 = 10'd40;
b_exp0 = 10'd349; b_exp1 = 10'd275; b_exp2 = 10'd570; b_exp3 = 10'd531;
a_sign0 = 4'd7; a_sign1 = 4'd11; a_sign2 = 4'd3; a_sign3 = 4'd9;
b_sign0 = 4'd12; b_sign1 = 4'd1; b_sign2 = 4'd2; b_sign3 = 4'd7;
@(posedge clk_i);
a_mant0 = 8'd119; a_mant1 = 8'd235; a_mant2 = 8'd170; a_mant3 = 8'd50;
b_mant0 = 8'd89; b_mant1 = 8'd143; b_mant2 = 8'd225; b_mant3 = 8'd45;
a_exp0 = 10'd913; a_exp1 = 10'd287; a_exp2 = 10'd546; a_exp3 = 10'd7;
b_exp0 = 10'd997; b_exp1 = 10'd81; b_exp2 = 10'd329; b_exp3 = 10'd900;
a_sign0 = 4'd2; a_sign1 = 4'd8; a_sign2 = 4'd13; a_sign3 = 4'd0;
b_sign0 = 4'd10; b_sign1 = 4'd9; b_sign2 = 4'd13; b_sign3 = 4'd1;
@(posedge clk_i);
a_mant0 = 8'd41; a_mant1 = 8'd178; a_mant2 = 8'd111; a_mant3 = 8'd18;
b_mant0 = 8'd23; b_mant1 = 8'd37; b_mant2 = 8'd132; b_mant3 = 8'd125;
a_exp0 = 10'd707; a_exp1 = 10'd605; a_exp2 = 10'd474; a_exp3 = 10'd998;
b_exp0 = 10'd405; b_exp1 = 10'd210; b_exp2 = 10'd283; b_exp3 = 10'd385;
a_sign0 = 4'd3; a_sign1 = 4'd1; a_sign2 = 4'd0; a_sign3 = 4'd16;
b_sign0 = 4'd3; b_sign1 = 4'd1; b_sign2 = 4'd11; b_sign3 = 4'd12;
@(posedge clk_i);
a_mant0 = 8'd98; a_mant1 = 8'd249; a_mant2 = 8'd250; a_mant3 = 8'd99;
b_mant0 = 8'd189; b_mant1 = 8'd105; b_mant2 = 8'd160; b_mant3 = 8'd223;
a_exp0 = 10'd18; a_exp1 = 10'd558; a_exp2 = 10'd922; a_exp3 = 10'd934;
b_exp0 = 10'd600; b_exp1 = 10'd485; b_exp2 = 10'd876; b_exp3 = 10'd839;
a_sign0 = 4'd13; a_sign1 = 4'd16; a_sign2 = 4'd14; a_sign3 = 4'd6;
b_sign0 = 4'd16; b_sign1 = 4'd9; b_sign2 = 4'd1; b_sign3 = 4'd14;
@(posedge clk_i);
a_mant0 = 8'd150; a_mant1 = 8'd234; a_mant2 = 8'd122; a_mant3 = 8'd200;
b_mant0 = 8'd41; b_mant1 = 8'd79; b_mant2 = 8'd63; b_mant3 = 8'd33;
a_exp0 = 10'd348; a_exp1 = 10'd721; a_exp2 = 10'd108; a_exp3 = 10'd883;
b_exp0 = 10'd50; b_exp1 = 10'd233; b_exp2 = 10'd442; b_exp3 = 10'd868;
a_sign0 = 4'd5; a_sign1 = 4'd16; a_sign2 = 4'd10; a_sign3 = 4'd5;
b_sign0 = 4'd16; b_sign1 = 4'd3; b_sign2 = 4'd15; b_sign3 = 4'd8;
@(posedge clk_i);
shared_exps0 = 8'd103;
shared_exps1 = 8'd131;
a_mant0 = 8'd61; a_mant1 = 8'd236; a_mant2 = 8'd60; a_mant3 = 8'd119;
b_mant0 = 8'd24; b_mant1 = 8'd152; b_mant2 = 8'd32; b_mant3 = 8'd38;
a_exp0 = 10'd230; a_exp1 = 10'd782; a_exp2 = 10'd382; a_exp3 = 10'd132;
b_exp0 = 10'd409; b_exp1 = 10'd626; b_exp2 = 10'd544; b_exp3 = 10'd459;
a_sign0 = 4'd1; a_sign1 = 4'd3; a_sign2 = 4'd14; a_sign3 = 4'd7;
b_sign0 = 4'd0; b_sign1 = 4'd15; b_sign2 = 4'd9; b_sign3 = 4'd3;
@(posedge clk_i);
a_mant0 = 8'd38; a_mant1 = 8'd174; a_mant2 = 8'd251; a_mant3 = 8'd150;
b_mant0 = 8'd216; b_mant1 = 8'd53; b_mant2 = 8'd83; b_mant3 = 8'd118;
a_exp0 = 10'd683; a_exp1 = 10'd250; a_exp2 = 10'd571; a_exp3 = 10'd64;
b_exp0 = 10'd271; b_exp1 = 10'd394; b_exp2 = 10'd793; b_exp3 = 10'd722;
a_sign0 = 4'd0; a_sign1 = 4'd8; a_sign2 = 4'd16; a_sign3 = 4'd9;
b_sign0 = 4'd3; b_sign1 = 4'd9; b_sign2 = 4'd15; b_sign3 = 4'd3;
@(posedge clk_i);
a_mant0 = 8'd6; a_mant1 = 8'd154; a_mant2 = 8'd108; a_mant3 = 8'd94;
b_mant0 = 8'd60; b_mant1 = 8'd104; b_mant2 = 8'd79; b_mant3 = 8'd232;
a_exp0 = 10'd312; a_exp1 = 10'd748; a_exp2 = 10'd207; a_exp3 = 10'd936;
b_exp0 = 10'd248; b_exp1 = 10'd665; b_exp2 = 10'd735; b_exp3 = 10'd153;
a_sign0 = 4'd5; a_sign1 = 4'd5; a_sign2 = 4'd5; a_sign3 = 4'd16;
b_sign0 = 4'd4; b_sign1 = 4'd12; b_sign2 = 4'd11; b_sign3 = 4'd1;
@(posedge clk_i);
a_mant0 = 8'd96; a_mant1 = 8'd35; a_mant2 = 8'd149; a_mant3 = 8'd248;
b_mant0 = 8'd15; b_mant1 = 8'd240; b_mant2 = 8'd55; b_mant3 = 8'd72;
a_exp0 = 10'd223; a_exp1 = 10'd788; a_exp2 = 10'd658; a_exp3 = 10'd748;
b_exp0 = 10'd609; b_exp1 = 10'd216; b_exp2 = 10'd255; b_exp3 = 10'd609;
a_sign0 = 4'd6; a_sign1 = 4'd16; a_sign2 = 4'd8; a_sign3 = 4'd12;
b_sign0 = 4'd5; b_sign1 = 4'd3; b_sign2 = 4'd15; b_sign3 = 4'd0;
@(posedge clk_i);
a_mant0 = 8'd197; a_mant1 = 8'd94; a_mant2 = 8'd27; a_mant3 = 8'd49;
b_mant0 = 8'd52; b_mant1 = 8'd40; b_mant2 = 8'd94; b_mant3 = 8'd86;
a_exp0 = 10'd942; a_exp1 = 10'd607; a_exp2 = 10'd127; a_exp3 = 10'd385;
b_exp0 = 10'd373; b_exp1 = 10'd915; b_exp2 = 10'd406; b_exp3 = 10'd396;
a_sign0 = 4'd2; a_sign1 = 4'd11; a_sign2 = 4'd8; a_sign3 = 4'd12;
b_sign0 = 4'd14; b_sign1 = 4'd16; b_sign2 = 4'd10; b_sign3 = 4'd3;
@(posedge clk_i);
a_mant0 = 8'd63; a_mant1 = 8'd133; a_mant2 = 8'd221; a_mant3 = 8'd127;
b_mant0 = 8'd78; b_mant1 = 8'd108; b_mant2 = 8'd216; b_mant3 = 8'd162;
a_exp0 = 10'd110; a_exp1 = 10'd207; a_exp2 = 10'd55; a_exp3 = 10'd187;
b_exp0 = 10'd654; b_exp1 = 10'd733; b_exp2 = 10'd329; b_exp3 = 10'd243;
a_sign0 = 4'd12; a_sign1 = 4'd10; a_sign2 = 4'd4; a_sign3 = 4'd13;
b_sign0 = 4'd14; b_sign1 = 4'd9; b_sign2 = 4'd5; b_sign3 = 4'd7;
@(posedge clk_i);
a_mant0 = 8'd255; a_mant1 = 8'd232; a_mant2 = 8'd139; a_mant3 = 8'd56;
b_mant0 = 8'd89; b_mant1 = 8'd213; b_mant2 = 8'd157; b_mant3 = 8'd202;
a_exp0 = 10'd156; a_exp1 = 10'd335; a_exp2 = 10'd897; a_exp3 = 10'd928;
b_exp0 = 10'd1000; b_exp1 = 10'd914; b_exp2 = 10'd812; b_exp3 = 10'd863;
a_sign0 = 4'd10; a_sign1 = 4'd15; a_sign2 = 4'd15; a_sign3 = 4'd8;
b_sign0 = 4'd12; b_sign1 = 4'd16; b_sign2 = 4'd16; b_sign3 = 4'd1;
@(posedge clk_i);
a_mant0 = 8'd197; a_mant1 = 8'd39; a_mant2 = 8'd202; a_mant3 = 8'd186;
b_mant0 = 8'd15; b_mant1 = 8'd190; b_mant2 = 8'd21; b_mant3 = 8'd230;
a_exp0 = 10'd811; a_exp1 = 10'd133; a_exp2 = 10'd69; a_exp3 = 10'd398;
b_exp0 = 10'd966; b_exp1 = 10'd822; b_exp2 = 10'd293; b_exp3 = 10'd252;
a_sign0 = 4'd15; a_sign1 = 4'd16; a_sign2 = 4'd1; a_sign3 = 4'd4;
b_sign0 = 4'd9; b_sign1 = 4'd12; b_sign2 = 4'd5; b_sign3 = 4'd3;
@(posedge clk_i);
shared_exps0 = 8'd149;
shared_exps1 = 8'd152;
rstn = 0;
@(posedge clk_i);
rstn = 1;
a_mant0 = 8'd209; a_mant1 = 8'd9; a_mant2 = 8'd21; a_mant3 = 8'd224;
b_mant0 = 8'd108; b_mant1 = 8'd102; b_mant2 = 8'd203; b_mant3 = 8'd207;
a_exp0 = 10'd1011; a_exp1 = 10'd354; a_exp2 = 10'd922; a_exp3 = 10'd828;
b_exp0 = 10'd588; b_exp1 = 10'd651; b_exp2 = 10'd273; b_exp3 = 10'd750;
a_sign0 = 4'd0; a_sign1 = 4'd3; a_sign2 = 4'd5; a_sign3 = 4'd2;
b_sign0 = 4'd4; b_sign1 = 4'd3; b_sign2 = 4'd1; b_sign3 = 4'd11;
@(posedge clk_i);
a_mant0 = 8'd194; a_mant1 = 8'd212; a_mant2 = 8'd154; a_mant3 = 8'd64;
b_mant0 = 8'd119; b_mant1 = 8'd247; b_mant2 = 8'd49; b_mant3 = 8'd169;
a_exp0 = 10'd579; a_exp1 = 10'd587; a_exp2 = 10'd525; a_exp3 = 10'd34;
b_exp0 = 10'd747; b_exp1 = 10'd706; b_exp2 = 10'd645; b_exp3 = 10'd590;
a_sign0 = 4'd9; a_sign1 = 4'd15; a_sign2 = 4'd2; a_sign3 = 4'd4;
b_sign0 = 4'd7; b_sign1 = 4'd3; b_sign2 = 4'd15; b_sign3 = 4'd7;
@(posedge clk_i);
a_mant0 = 8'd9; a_mant1 = 8'd245; a_mant2 = 8'd155; a_mant3 = 8'd45;
b_mant0 = 8'd190; b_mant1 = 8'd132; b_mant2 = 8'd189; b_mant3 = 8'd53;
a_exp0 = 10'd786; a_exp1 = 10'd470; a_exp2 = 10'd282; a_exp3 = 10'd399;
b_exp0 = 10'd870; b_exp1 = 10'd273; b_exp2 = 10'd583; b_exp3 = 10'd1022;
a_sign0 = 4'd16; a_sign1 = 4'd13; a_sign2 = 4'd0; a_sign3 = 4'd15;
b_sign0 = 4'd1; b_sign1 = 4'd15; b_sign2 = 4'd10; b_sign3 = 4'd14;
@(posedge clk_i);
a_mant0 = 8'd204; a_mant1 = 8'd151; a_mant2 = 8'd255; a_mant3 = 8'd98;
b_mant0 = 8'd79; b_mant1 = 8'd82; b_mant2 = 8'd54; b_mant3 = 8'd245;
a_exp0 = 10'd553; a_exp1 = 10'd397; a_exp2 = 10'd719; a_exp3 = 10'd394;
b_exp0 = 10'd187; b_exp1 = 10'd813; b_exp2 = 10'd448; b_exp3 = 10'd565;
a_sign0 = 4'd6; a_sign1 = 4'd0; a_sign2 = 4'd7; a_sign3 = 4'd15;
b_sign0 = 4'd11; b_sign1 = 4'd12; b_sign2 = 4'd15; b_sign3 = 4'd1;
@(posedge clk_i);
a_mant0 = 8'd146; a_mant1 = 8'd145; a_mant2 = 8'd227; a_mant3 = 8'd6;
b_mant0 = 8'd106; b_mant1 = 8'd52; b_mant2 = 8'd114; b_mant3 = 8'd78;
a_exp0 = 10'd426; a_exp1 = 10'd1009; a_exp2 = 10'd116; a_exp3 = 10'd967;
b_exp0 = 10'd715; b_exp1 = 10'd615; b_exp2 = 10'd27; b_exp3 = 10'd258;
a_sign0 = 4'd7; a_sign1 = 4'd8; a_sign2 = 4'd10; a_sign3 = 4'd3;
b_sign0 = 4'd11; b_sign1 = 4'd8; b_sign2 = 4'd13; b_sign3 = 4'd12;
@(posedge clk_i);
a_mant0 = 8'd140; a_mant1 = 8'd142; a_mant2 = 8'd184; a_mant3 = 8'd60;
b_mant0 = 8'd135; b_mant1 = 8'd208; b_mant2 = 8'd119; b_mant3 = 8'd197;
a_exp0 = 10'd347; a_exp1 = 10'd760; a_exp2 = 10'd650; a_exp3 = 10'd870;
b_exp0 = 10'd857; b_exp1 = 10'd530; b_exp2 = 10'd879; b_exp3 = 10'd562;
a_sign0 = 4'd1; a_sign1 = 4'd0; a_sign2 = 4'd5; a_sign3 = 4'd12;
b_sign0 = 4'd0; b_sign1 = 4'd5; b_sign2 = 4'd1; b_sign3 = 4'd1;
@(posedge clk_i);
a_mant0 = 8'd87; a_mant1 = 8'd152; a_mant2 = 8'd63; a_mant3 = 8'd200;
b_mant0 = 8'd119; b_mant1 = 8'd115; b_mant2 = 8'd229; b_mant3 = 8'd60;
a_exp0 = 10'd111; a_exp1 = 10'd650; a_exp2 = 10'd233; a_exp3 = 10'd54;
b_exp0 = 10'd922; b_exp1 = 10'd371; b_exp2 = 10'd332; b_exp3 = 10'd347;
a_sign0 = 4'd2; a_sign1 = 4'd10; a_sign2 = 4'd11; a_sign3 = 4'd0;
b_sign0 = 4'd6; b_sign1 = 4'd8; b_sign2 = 4'd2; b_sign3 = 4'd8;
@(posedge clk_i);
shared_exps0 = 8'd125;
shared_exps1 = 8'd118;
a_mant0 = 8'd82; a_mant1 = 8'd14; a_mant2 = 8'd84; a_mant3 = 8'd205;
b_mant0 = 8'd170; b_mant1 = 8'd238; b_mant2 = 8'd124; b_mant3 = 8'd93;
a_exp0 = 10'd794; a_exp1 = 10'd281; a_exp2 = 10'd369; a_exp3 = 10'd50;
b_exp0 = 10'd425; b_exp1 = 10'd210; b_exp2 = 10'd802; b_exp3 = 10'd863;
a_sign0 = 4'd13; a_sign1 = 4'd4; a_sign2 = 4'd4; a_sign3 = 4'd7;
b_sign0 = 4'd5; b_sign1 = 4'd5; b_sign2 = 4'd9; b_sign3 = 4'd2;
@(posedge clk_i);
a_mant0 = 8'd188; a_mant1 = 8'd102; a_mant2 = 8'd235; a_mant3 = 8'd237;
b_mant0 = 8'd108; b_mant1 = 8'd2; b_mant2 = 8'd147; b_mant3 = 8'd14;
a_exp0 = 10'd484; a_exp1 = 10'd849; a_exp2 = 10'd281; a_exp3 = 10'd988;
b_exp0 = 10'd45; b_exp1 = 10'd615; b_exp2 = 10'd569; b_exp3 = 10'd642;
a_sign0 = 4'd10; a_sign1 = 4'd2; a_sign2 = 4'd13; a_sign3 = 4'd1;
b_sign0 = 4'd0; b_sign1 = 4'd3; b_sign2 = 4'd1; b_sign3 = 4'd15;
@(posedge clk_i);
a_mant0 = 8'd227; a_mant1 = 8'd227; a_mant2 = 8'd92; a_mant3 = 8'd172;
b_mant0 = 8'd200; b_mant1 = 8'd135; b_mant2 = 8'd234; b_mant3 = 8'd219;
a_exp0 = 10'd954; a_exp1 = 10'd955; a_exp2 = 10'd35; a_exp3 = 10'd836;
b_exp0 = 10'd33; b_exp1 = 10'd711; b_exp2 = 10'd969; b_exp3 = 10'd896;
a_sign0 = 4'd11; a_sign1 = 4'd7; a_sign2 = 4'd14; a_sign3 = 4'd12;
b_sign0 = 4'd15; b_sign1 = 4'd2; b_sign2 = 4'd2; b_sign3 = 4'd2;
@(posedge clk_i);
a_mant0 = 8'd167; a_mant1 = 8'd48; a_mant2 = 8'd149; a_mant3 = 8'd104;
b_mant0 = 8'd28; b_mant1 = 8'd183; b_mant2 = 8'd60; b_mant3 = 8'd147;
a_exp0 = 10'd30; a_exp1 = 10'd357; a_exp2 = 10'd438; a_exp3 = 10'd857;
b_exp0 = 10'd987; b_exp1 = 10'd184; b_exp2 = 10'd9; b_exp3 = 10'd586;
a_sign0 = 4'd8; a_sign1 = 4'd6; a_sign2 = 4'd10; a_sign3 = 4'd13;
b_sign0 = 4'd12; b_sign1 = 4'd6; b_sign2 = 4'd9; b_sign3 = 4'd0;
@(posedge clk_i);
a_mant0 = 8'd172; a_mant1 = 8'd142; a_mant2 = 8'd145; a_mant3 = 8'd119;
b_mant0 = 8'd52; b_mant1 = 8'd153; b_mant2 = 8'd50; b_mant3 = 8'd70;
a_exp0 = 10'd790; a_exp1 = 10'd772; a_exp2 = 10'd583; a_exp3 = 10'd421;
b_exp0 = 10'd263; b_exp1 = 10'd266; b_exp2 = 10'd214; b_exp3 = 10'd118;
a_sign0 = 4'd1; a_sign1 = 4'd0; a_sign2 = 4'd1; a_sign3 = 4'd13;
b_sign0 = 4'd7; b_sign1 = 4'd11; b_sign2 = 4'd8; b_sign3 = 4'd4;
@(posedge clk_i);
a_mant0 = 8'd103; a_mant1 = 8'd8; a_mant2 = 8'd193; a_mant3 = 8'd199;
b_mant0 = 8'd241; b_mant1 = 8'd137; b_mant2 = 8'd190; b_mant3 = 8'd85;
a_exp0 = 10'd692; a_exp1 = 10'd117; a_exp2 = 10'd521; a_exp3 = 10'd744;
b_exp0 = 10'd607; b_exp1 = 10'd942; b_exp2 = 10'd636; b_exp3 = 10'd172;
a_sign0 = 4'd12; a_sign1 = 4'd0; a_sign2 = 4'd14; a_sign3 = 4'd9;
b_sign0 = 4'd14; b_sign1 = 4'd5; b_sign2 = 4'd13; b_sign3 = 4'd0;
@(posedge clk_i);
a_mant0 = 8'd247; a_mant1 = 8'd95; a_mant2 = 8'd155; a_mant3 = 8'd110;
b_mant0 = 8'd168; b_mant1 = 8'd37; b_mant2 = 8'd33; b_mant3 = 8'd153;
a_exp0 = 10'd843; a_exp1 = 10'd54; a_exp2 = 10'd727; a_exp3 = 10'd733;
b_exp0 = 10'd905; b_exp1 = 10'd159; b_exp2 = 10'd940; b_exp3 = 10'd64;
a_sign0 = 4'd10; a_sign1 = 4'd3; a_sign2 = 4'd9; a_sign3 = 4'd10;
b_sign0 = 4'd13; b_sign1 = 4'd4; b_sign2 = 4'd7; b_sign3 = 4'd14;
@(posedge clk_i);
a_mant0 = 8'd185; a_mant1 = 8'd158; a_mant2 = 8'd10; a_mant3 = 8'd6;
b_mant0 = 8'd175; b_mant1 = 8'd255; b_mant2 = 8'd174; b_mant3 = 8'd45;
a_exp0 = 10'd846; a_exp1 = 10'd298; a_exp2 = 10'd610; a_exp3 = 10'd942;
b_exp0 = 10'd695; b_exp1 = 10'd718; b_exp2 = 10'd777; b_exp3 = 10'd245;
a_sign0 = 4'd2; a_sign1 = 4'd5; a_sign2 = 4'd2; a_sign3 = 4'd5;
b_sign0 = 4'd14; b_sign1 = 4'd13; b_sign2 = 4'd3; b_sign3 = 4'd3;
@(posedge clk_i);
shared_exps0 = 8'd138;
shared_exps1 = 8'd147;
a_mant0 = 8'd87; a_mant1 = 8'd176; a_mant2 = 8'd57; a_mant3 = 8'd46;
b_mant0 = 8'd121; b_mant1 = 8'd16; b_mant2 = 8'd66; b_mant3 = 8'd175;
a_exp0 = 10'd43; a_exp1 = 10'd244; a_exp2 = 10'd652; a_exp3 = 10'd1001;
b_exp0 = 10'd149; b_exp1 = 10'd944; b_exp2 = 10'd117; b_exp3 = 10'd765;
a_sign0 = 4'd7; a_sign1 = 4'd8; a_sign2 = 4'd7; a_sign3 = 4'd12;
b_sign0 = 4'd11; b_sign1 = 4'd2; b_sign2 = 4'd14; b_sign3 = 4'd10;
@(posedge clk_i);
a_mant0 = 8'd214; a_mant1 = 8'd203; a_mant2 = 8'd130; a_mant3 = 8'd113;
b_mant0 = 8'd132; b_mant1 = 8'd225; b_mant2 = 8'd215; b_mant3 = 8'd18;
a_exp0 = 10'd104; a_exp1 = 10'd233; a_exp2 = 10'd924; a_exp3 = 10'd222;
b_exp0 = 10'd1011; b_exp1 = 10'd526; b_exp2 = 10'd620; b_exp3 = 10'd304;
a_sign0 = 4'd5; a_sign1 = 4'd14; a_sign2 = 4'd0; a_sign3 = 4'd7;
b_sign0 = 4'd3; b_sign1 = 4'd1; b_sign2 = 4'd4; b_sign3 = 4'd1;
@(posedge clk_i);
a_mant0 = 8'd110; a_mant1 = 8'd54; a_mant2 = 8'd112; a_mant3 = 8'd128;
b_mant0 = 8'd183; b_mant1 = 8'd27; b_mant2 = 8'd110; b_mant3 = 8'd106;
a_exp0 = 10'd150; a_exp1 = 10'd915; a_exp2 = 10'd465; a_exp3 = 10'd940;
b_exp0 = 10'd911; b_exp1 = 10'd446; b_exp2 = 10'd729; b_exp3 = 10'd653;
a_sign0 = 4'd12; a_sign1 = 4'd13; a_sign2 = 4'd10; a_sign3 = 4'd4;
b_sign0 = 4'd7; b_sign1 = 4'd7; b_sign2 = 4'd16; b_sign3 = 4'd5;
@(posedge clk_i);
a_mant0 = 8'd99; a_mant1 = 8'd94; a_mant2 = 8'd106; a_mant3 = 8'd225;
b_mant0 = 8'd251; b_mant1 = 8'd44; b_mant2 = 8'd162; b_mant3 = 8'd15;
a_exp0 = 10'd394; a_exp1 = 10'd882; a_exp2 = 10'd1006; a_exp3 = 10'd320;
b_exp0 = 10'd805; b_exp1 = 10'd1017; b_exp2 = 10'd982; b_exp3 = 10'd495;
a_sign0 = 4'd13; a_sign1 = 4'd0; a_sign2 = 4'd6; a_sign3 = 4'd16;
b_sign0 = 4'd11; b_sign1 = 4'd12; b_sign2 = 4'd6; b_sign3 = 4'd10;
@(posedge clk_i);
a_mant0 = 8'd12; a_mant1 = 8'd214; a_mant2 = 8'd49; a_mant3 = 8'd162;
b_mant0 = 8'd88; b_mant1 = 8'd245; b_mant2 = 8'd144; b_mant3 = 8'd88;
a_exp0 = 10'd234; a_exp1 = 10'd874; a_exp2 = 10'd551; a_exp3 = 10'd851;
b_exp0 = 10'd453; b_exp1 = 10'd264; b_exp2 = 10'd378; b_exp3 = 10'd127;
a_sign0 = 4'd16; a_sign1 = 4'd14; a_sign2 = 4'd6; a_sign3 = 4'd14;
b_sign0 = 4'd1; b_sign1 = 4'd9; b_sign2 = 4'd7; b_sign3 = 4'd11;
@(posedge clk_i);
a_mant0 = 8'd215; a_mant1 = 8'd109; a_mant2 = 8'd136; a_mant3 = 8'd156;
b_mant0 = 8'd211; b_mant1 = 8'd152; b_mant2 = 8'd252; b_mant3 = 8'd78;
a_exp0 = 10'd584; a_exp1 = 10'd137; a_exp2 = 10'd287; a_exp3 = 10'd886;
b_exp0 = 10'd320; b_exp1 = 10'd746; b_exp2 = 10'd561; b_exp3 = 10'd674;
a_sign0 = 4'd6; a_sign1 = 4'd14; a_sign2 = 4'd8; a_sign3 = 4'd9;
b_sign0 = 4'd5; b_sign1 = 4'd11; b_sign2 = 4'd6; b_sign3 = 4'd5;
@(posedge clk_i);
a_mant0 = 8'd15; a_mant1 = 8'd158; a_mant2 = 8'd20; a_mant3 = 8'd176;
b_mant0 = 8'd215; b_mant1 = 8'd27; b_mant2 = 8'd163; b_mant3 = 8'd160;
a_exp0 = 10'd82; a_exp1 = 10'd56; a_exp2 = 10'd555; a_exp3 = 10'd10;
b_exp0 = 10'd201; b_exp1 = 10'd20; b_exp2 = 10'd918; b_exp3 = 10'd587;
a_sign0 = 4'd0; a_sign1 = 4'd5; a_sign2 = 4'd6; a_sign3 = 4'd10;
b_sign0 = 4'd3; b_sign1 = 4'd16; b_sign2 = 4'd1; b_sign3 = 4'd13;
@(posedge clk_i);
a_mant0 = 8'd93; a_mant1 = 8'd68; a_mant2 = 8'd163; a_mant3 = 8'd170;
b_mant0 = 8'd227; b_mant1 = 8'd113; b_mant2 = 8'd17; b_mant3 = 8'd118;
a_exp0 = 10'd563; a_exp1 = 10'd308; a_exp2 = 10'd483; a_exp3 = 10'd389;
b_exp0 = 10'd866; b_exp1 = 10'd48; b_exp2 = 10'd112; b_exp3 = 10'd916;
a_sign0 = 4'd1; a_sign1 = 4'd14; a_sign2 = 4'd4; a_sign3 = 4'd10;
b_sign0 = 4'd0; b_sign1 = 4'd2; b_sign2 = 4'd13; b_sign3 = 4'd1;
@(posedge clk_i);
shared_exps0 = 8'd136;
shared_exps1 = 8'd123;
a_mant0 = 8'd245; a_mant1 = 8'd142; a_mant2 = 8'd130; a_mant3 = 8'd88;
b_mant0 = 8'd53; b_mant1 = 8'd14; b_mant2 = 8'd3; b_mant3 = 8'd25;
a_exp0 = 10'd463; a_exp1 = 10'd727; a_exp2 = 10'd410; a_exp3 = 10'd532;
b_exp0 = 10'd979; b_exp1 = 10'd111; b_exp2 = 10'd664; b_exp3 = 10'd82;
a_sign0 = 4'd3; a_sign1 = 4'd16; a_sign2 = 4'd9; a_sign3 = 4'd13;
b_sign0 = 4'd4; b_sign1 = 4'd2; b_sign2 = 4'd13; b_sign3 = 4'd12;
@(posedge clk_i);
a_mant0 = 8'd61; a_mant1 = 8'd104; a_mant2 = 8'd114; a_mant3 = 8'd156;
b_mant0 = 8'd200; b_mant1 = 8'd208; b_mant2 = 8'd178; b_mant3 = 8'd111;
a_exp0 = 10'd534; a_exp1 = 10'd130; a_exp2 = 10'd942; a_exp3 = 10'd615;
b_exp0 = 10'd413; b_exp1 = 10'd469; b_exp2 = 10'd470; b_exp3 = 10'd772;
a_sign0 = 4'd2; a_sign1 = 4'd5; a_sign2 = 4'd11; a_sign3 = 4'd7;
b_sign0 = 4'd10; b_sign1 = 4'd9; b_sign2 = 4'd13; b_sign3 = 4'd11;
@(posedge clk_i);
a_mant0 = 8'd240; a_mant1 = 8'd95; a_mant2 = 8'd196; a_mant3 = 8'd157;
b_mant0 = 8'd124; b_mant1 = 8'd26; b_mant2 = 8'd63; b_mant3 = 8'd5;
a_exp0 = 10'd320; a_exp1 = 10'd840; a_exp2 = 10'd794; a_exp3 = 10'd855;
b_exp0 = 10'd35; b_exp1 = 10'd97; b_exp2 = 10'd590; b_exp3 = 10'd763;
a_sign0 = 4'd1; a_sign1 = 4'd4; a_sign2 = 4'd10; a_sign3 = 4'd7;
b_sign0 = 4'd4; b_sign1 = 4'd10; b_sign2 = 4'd8; b_sign3 = 4'd1;
@(posedge clk_i);
a_mant0 = 8'd189; a_mant1 = 8'd246; a_mant2 = 8'd214; a_mant3 = 8'd58;
b_mant0 = 8'd196; b_mant1 = 8'd147; b_mant2 = 8'd175; b_mant3 = 8'd149;
a_exp0 = 10'd803; a_exp1 = 10'd996; a_exp2 = 10'd376; a_exp3 = 10'd433;
b_exp0 = 10'd626; b_exp1 = 10'd663; b_exp2 = 10'd329; b_exp3 = 10'd299;
a_sign0 = 4'd2; a_sign1 = 4'd8; a_sign2 = 4'd10; a_sign3 = 4'd12;
b_sign0 = 4'd0; b_sign1 = 4'd3; b_sign2 = 4'd10; b_sign3 = 4'd14;
@(posedge clk_i);
a_mant0 = 8'd123; a_mant1 = 8'd189; a_mant2 = 8'd239; a_mant3 = 8'd249;
b_mant0 = 8'd109; b_mant1 = 8'd32; b_mant2 = 8'd199; b_mant3 = 8'd251;
a_exp0 = 10'd913; a_exp1 = 10'd480; a_exp2 = 10'd156; a_exp3 = 10'd190;
b_exp0 = 10'd809; b_exp1 = 10'd61; b_exp2 = 10'd754; b_exp3 = 10'd845;
a_sign0 = 4'd15; a_sign1 = 4'd12; a_sign2 = 4'd11; a_sign3 = 4'd15;
b_sign0 = 4'd7; b_sign1 = 4'd10; b_sign2 = 4'd0; b_sign3 = 4'd11;
@(posedge clk_i);
a_mant0 = 8'd255; a_mant1 = 8'd109; a_mant2 = 8'd200; a_mant3 = 8'd40;
b_mant0 = 8'd166; b_mant1 = 8'd149; b_mant2 = 8'd174; b_mant3 = 8'd117;
a_exp0 = 10'd183; a_exp1 = 10'd1010; a_exp2 = 10'd584; a_exp3 = 10'd621;
b_exp0 = 10'd310; b_exp1 = 10'd649; b_exp2 = 10'd396; b_exp3 = 10'd539;
a_sign0 = 4'd5; a_sign1 = 4'd7; a_sign2 = 4'd11; a_sign3 = 4'd11;
b_sign0 = 4'd12; b_sign1 = 4'd12; b_sign2 = 4'd9; b_sign3 = 4'd3;
@(posedge clk_i);
a_mant0 = 8'd16; a_mant1 = 8'd205; a_mant2 = 8'd229; a_mant3 = 8'd1;
b_mant0 = 8'd16; b_mant1 = 8'd10; b_mant2 = 8'd6; b_mant3 = 8'd80;
a_exp0 = 10'd20; a_exp1 = 10'd709; a_exp2 = 10'd368; a_exp3 = 10'd841;
b_exp0 = 10'd241; b_exp1 = 10'd919; b_exp2 = 10'd429; b_exp3 = 10'd568;
a_sign0 = 4'd15; a_sign1 = 4'd5; a_sign2 = 4'd2; a_sign3 = 4'd5;
b_sign0 = 4'd16; b_sign1 = 4'd9; b_sign2 = 4'd6; b_sign3 = 4'd5;
@(posedge clk_i);
a_mant0 = 8'd144; a_mant1 = 8'd193; a_mant2 = 8'd121; a_mant3 = 8'd107;
b_mant0 = 8'd9; b_mant1 = 8'd210; b_mant2 = 8'd60; b_mant3 = 8'd209;
a_exp0 = 10'd338; a_exp1 = 10'd607; a_exp2 = 10'd86; a_exp3 = 10'd324;
b_exp0 = 10'd973; b_exp1 = 10'd75; b_exp2 = 10'd291; b_exp3 = 10'd357;
a_sign0 = 4'd11; a_sign1 = 4'd16; a_sign2 = 4'd6; a_sign3 = 4'd5;
b_sign0 = 4'd7; b_sign1 = 4'd10; b_sign2 = 4'd5; b_sign3 = 4'd16;
@(posedge clk_i);
shared_exps0 = 8'd152;
shared_exps1 = 8'd126;
rstn = 0;
@(posedge clk_i);
rstn = 1;
a_mant0 = 8'd81; a_mant1 = 8'd170; a_mant2 = 8'd63; a_mant3 = 8'd97;
b_mant0 = 8'd235; b_mant1 = 8'd55; b_mant2 = 8'd216; b_mant3 = 8'd173;
a_exp0 = 10'd849; a_exp1 = 10'd199; a_exp2 = 10'd387; a_exp3 = 10'd235;
b_exp0 = 10'd149; b_exp1 = 10'd62; b_exp2 = 10'd160; b_exp3 = 10'd787;
a_sign0 = 4'd4; a_sign1 = 4'd11; a_sign2 = 4'd6; a_sign3 = 4'd4;
b_sign0 = 4'd6; b_sign1 = 4'd1; b_sign2 = 4'd4; b_sign3 = 4'd9;
@(posedge clk_i);
a_mant0 = 8'd40; a_mant1 = 8'd27; a_mant2 = 8'd198; a_mant3 = 8'd35;
b_mant0 = 8'd128; b_mant1 = 8'd229; b_mant2 = 8'd31; b_mant3 = 8'd60;
a_exp0 = 10'd866; a_exp1 = 10'd529; a_exp2 = 10'd487; a_exp3 = 10'd902;
b_exp0 = 10'd206; b_exp1 = 10'd494; b_exp2 = 10'd914; b_exp3 = 10'd145;
a_sign0 = 4'd3; a_sign1 = 4'd15; a_sign2 = 4'd9; a_sign3 = 4'd4;
b_sign0 = 4'd16; b_sign1 = 4'd3; b_sign2 = 4'd16; b_sign3 = 4'd0;
@(posedge clk_i);
a_mant0 = 8'd216; a_mant1 = 8'd199; a_mant2 = 8'd149; a_mant3 = 8'd141;
b_mant0 = 8'd109; b_mant1 = 8'd103; b_mant2 = 8'd246; b_mant3 = 8'd91;
a_exp0 = 10'd640; a_exp1 = 10'd359; a_exp2 = 10'd433; a_exp3 = 10'd188;
b_exp0 = 10'd635; b_exp1 = 10'd769; b_exp2 = 10'd358; b_exp3 = 10'd316;
a_sign0 = 4'd16; a_sign1 = 4'd15; a_sign2 = 4'd0; a_sign3 = 4'd13;
b_sign0 = 4'd3; b_sign1 = 4'd14; b_sign2 = 4'd5; b_sign3 = 4'd13;
@(posedge clk_i);
a_mant0 = 8'd35; a_mant1 = 8'd28; a_mant2 = 8'd40; a_mant3 = 8'd71;
b_mant0 = 8'd202; b_mant1 = 8'd81; b_mant2 = 8'd229; b_mant3 = 8'd223;
a_exp0 = 10'd478; a_exp1 = 10'd181; a_exp2 = 10'd851; a_exp3 = 10'd214;
b_exp0 = 10'd794; b_exp1 = 10'd433; b_exp2 = 10'd302; b_exp3 = 10'd119;
a_sign0 = 4'd1; a_sign1 = 4'd10; a_sign2 = 4'd6; a_sign3 = 4'd13;
b_sign0 = 4'd4; b_sign1 = 4'd8; b_sign2 = 4'd4; b_sign3 = 4'd12;
@(posedge clk_i);
a_mant0 = 8'd214; a_mant1 = 8'd134; a_mant2 = 8'd99; a_mant3 = 8'd131;
b_mant0 = 8'd151; b_mant1 = 8'd22; b_mant2 = 8'd151; b_mant3 = 8'd163;
a_exp0 = 10'd14; a_exp1 = 10'd721; a_exp2 = 10'd902; a_exp3 = 10'd838;
b_exp0 = 10'd210; b_exp1 = 10'd373; b_exp2 = 10'd959; b_exp3 = 10'd144;
a_sign0 = 4'd16; a_sign1 = 4'd9; a_sign2 = 4'd1; a_sign3 = 4'd9;
b_sign0 = 4'd16; b_sign1 = 4'd1; b_sign2 = 4'd9; b_sign3 = 4'd12;
@(posedge clk_i);
a_mant0 = 8'd117; a_mant1 = 8'd194; a_mant2 = 8'd186; a_mant3 = 8'd226;
b_mant0 = 8'd76; b_mant1 = 8'd186; b_mant2 = 8'd145; b_mant3 = 8'd99;
a_exp0 = 10'd233; a_exp1 = 10'd716; a_exp2 = 10'd21; a_exp3 = 10'd261;
b_exp0 = 10'd655; b_exp1 = 10'd164; b_exp2 = 10'd602; b_exp3 = 10'd254;
a_sign0 = 4'd15; a_sign1 = 4'd5; a_sign2 = 4'd14; a_sign3 = 4'd7;
b_sign0 = 4'd8; b_sign1 = 4'd14; b_sign2 = 4'd12; b_sign3 = 4'd6;
@(posedge clk_i);
a_mant0 = 8'd245; a_mant1 = 8'd110; a_mant2 = 8'd181; a_mant3 = 8'd32;
b_mant0 = 8'd157; b_mant1 = 8'd162; b_mant2 = 8'd153; b_mant3 = 8'd212;
a_exp0 = 10'd205; a_exp1 = 10'd915; a_exp2 = 10'd89; a_exp3 = 10'd357;
b_exp0 = 10'd461; b_exp1 = 10'd794; b_exp2 = 10'd657; b_exp3 = 10'd477;
a_sign0 = 4'd11; a_sign1 = 4'd5; a_sign2 = 4'd7; a_sign3 = 4'd12;
b_sign0 = 4'd8; b_sign1 = 4'd7; b_sign2 = 4'd1; b_sign3 = 4'd2;
@(posedge clk_i);
shared_exps0 = 8'd132;
shared_exps1 = 8'd143;
a_mant0 = 8'd113; a_mant1 = 8'd63; a_mant2 = 8'd78; a_mant3 = 8'd106;
b_mant0 = 8'd71; b_mant1 = 8'd108; b_mant2 = 8'd199; b_mant3 = 8'd147;
a_exp0 = 10'd864; a_exp1 = 10'd664; a_exp2 = 10'd787; a_exp3 = 10'd432;
b_exp0 = 10'd961; b_exp1 = 10'd662; b_exp2 = 10'd423; b_exp3 = 10'd571;
a_sign0 = 4'd14; a_sign1 = 4'd14; a_sign2 = 4'd16; a_sign3 = 4'd5;
b_sign0 = 4'd10; b_sign1 = 4'd13; b_sign2 = 4'd12; b_sign3 = 4'd14;
@(posedge clk_i);
a_mant0 = 8'd115; a_mant1 = 8'd48; a_mant2 = 8'd140; a_mant3 = 8'd9;
b_mant0 = 8'd177; b_mant1 = 8'd170; b_mant2 = 8'd174; b_mant3 = 8'd77;
a_exp0 = 10'd735; a_exp1 = 10'd971; a_exp2 = 10'd640; a_exp3 = 10'd610;
b_exp0 = 10'd686; b_exp1 = 10'd610; b_exp2 = 10'd281; b_exp3 = 10'd29;
a_sign0 = 4'd6; a_sign1 = 4'd2; a_sign2 = 4'd7; a_sign3 = 4'd6;
b_sign0 = 4'd8; b_sign1 = 4'd14; b_sign2 = 4'd12; b_sign3 = 4'd16;
@(posedge clk_i);
a_mant0 = 8'd248; a_mant1 = 8'd79; a_mant2 = 8'd110; a_mant3 = 8'd114;
b_mant0 = 8'd115; b_mant1 = 8'd111; b_mant2 = 8'd109; b_mant3 = 8'd61;
a_exp0 = 10'd116; a_exp1 = 10'd63; a_exp2 = 10'd155; a_exp3 = 10'd444;
b_exp0 = 10'd1015; b_exp1 = 10'd182; b_exp2 = 10'd780; b_exp3 = 10'd301;
a_sign0 = 4'd9; a_sign1 = 4'd0; a_sign2 = 4'd11; a_sign3 = 4'd14;
b_sign0 = 4'd10; b_sign1 = 4'd8; b_sign2 = 4'd11; b_sign3 = 4'd11;
@(posedge clk_i);
a_mant0 = 8'd85; a_mant1 = 8'd4; a_mant2 = 8'd127; a_mant3 = 8'd49;
b_mant0 = 8'd105; b_mant1 = 8'd83; b_mant2 = 8'd165; b_mant3 = 8'd43;
a_exp0 = 10'd634; a_exp1 = 10'd243; a_exp2 = 10'd343; a_exp3 = 10'd12;
b_exp0 = 10'd297; b_exp1 = 10'd218; b_exp2 = 10'd551; b_exp3 = 10'd15;
a_sign0 = 4'd5; a_sign1 = 4'd13; a_sign2 = 4'd10; a_sign3 = 4'd2;
b_sign0 = 4'd7; b_sign1 = 4'd10; b_sign2 = 4'd2; b_sign3 = 4'd7;
@(posedge clk_i);
a_mant0 = 8'd91; a_mant1 = 8'd225; a_mant2 = 8'd177; a_mant3 = 8'd72;
b_mant0 = 8'd121; b_mant1 = 8'd221; b_mant2 = 8'd209; b_mant3 = 8'd237;
a_exp0 = 10'd204; a_exp1 = 10'd18; a_exp2 = 10'd250; a_exp3 = 10'd916;
b_exp0 = 10'd473; b_exp1 = 10'd251; b_exp2 = 10'd803; b_exp3 = 10'd103;
a_sign0 = 4'd12; a_sign1 = 4'd6; a_sign2 = 4'd7; a_sign3 = 4'd14;
b_sign0 = 4'd2; b_sign1 = 4'd13; b_sign2 = 4'd9; b_sign3 = 4'd15;
@(posedge clk_i);
a_mant0 = 8'd201; a_mant1 = 8'd40; a_mant2 = 8'd252; a_mant3 = 8'd211;
b_mant0 = 8'd244; b_mant1 = 8'd120; b_mant2 = 8'd126; b_mant3 = 8'd149;
a_exp0 = 10'd825; a_exp1 = 10'd462; a_exp2 = 10'd298; a_exp3 = 10'd405;
b_exp0 = 10'd700; b_exp1 = 10'd555; b_exp2 = 10'd554; b_exp3 = 10'd232;
a_sign0 = 4'd15; a_sign1 = 4'd6; a_sign2 = 4'd9; a_sign3 = 4'd6;
b_sign0 = 4'd1; b_sign1 = 4'd12; b_sign2 = 4'd4; b_sign3 = 4'd13;
@(posedge clk_i);
a_mant0 = 8'd8; a_mant1 = 8'd112; a_mant2 = 8'd130; a_mant3 = 8'd159;
b_mant0 = 8'd128; b_mant1 = 8'd53; b_mant2 = 8'd156; b_mant3 = 8'd196;
a_exp0 = 10'd660; a_exp1 = 10'd317; a_exp2 = 10'd584; a_exp3 = 10'd459;
b_exp0 = 10'd87; b_exp1 = 10'd744; b_exp2 = 10'd631; b_exp3 = 10'd992;
a_sign0 = 4'd1; a_sign1 = 4'd16; a_sign2 = 4'd4; a_sign3 = 4'd15;
b_sign0 = 4'd8; b_sign1 = 4'd1; b_sign2 = 4'd7; b_sign3 = 4'd5;
@(posedge clk_i);
a_mant0 = 8'd23; a_mant1 = 8'd46; a_mant2 = 8'd41; a_mant3 = 8'd121;
b_mant0 = 8'd90; b_mant1 = 8'd111; b_mant2 = 8'd75; b_mant3 = 8'd75;
a_exp0 = 10'd811; a_exp1 = 10'd290; a_exp2 = 10'd890; a_exp3 = 10'd266;
b_exp0 = 10'd437; b_exp1 = 10'd196; b_exp2 = 10'd909; b_exp3 = 10'd345;
a_sign0 = 4'd15; a_sign1 = 4'd4; a_sign2 = 4'd8; a_sign3 = 4'd4;
b_sign0 = 4'd14; b_sign1 = 4'd14; b_sign2 = 4'd3; b_sign3 = 4'd9;
@(posedge clk_i);
shared_exps0 = 8'd129;
shared_exps1 = 8'd113;
a_mant0 = 8'd5; a_mant1 = 8'd234; a_mant2 = 8'd122; a_mant3 = 8'd53;
b_mant0 = 8'd142; b_mant1 = 8'd116; b_mant2 = 8'd86; b_mant3 = 8'd68;
a_exp0 = 10'd340; a_exp1 = 10'd882; a_exp2 = 10'd624; a_exp3 = 10'd163;
b_exp0 = 10'd260; b_exp1 = 10'd600; b_exp2 = 10'd340; b_exp3 = 10'd876;
a_sign0 = 4'd10; a_sign1 = 4'd8; a_sign2 = 4'd14; a_sign3 = 4'd13;
b_sign0 = 4'd10; b_sign1 = 4'd10; b_sign2 = 4'd16; b_sign3 = 4'd1;
@(posedge clk_i);
a_mant0 = 8'd9; a_mant1 = 8'd222; a_mant2 = 8'd53; a_mant3 = 8'd51;
b_mant0 = 8'd216; b_mant1 = 8'd233; b_mant2 = 8'd5; b_mant3 = 8'd101;
a_exp0 = 10'd118; a_exp1 = 10'd759; a_exp2 = 10'd952; a_exp3 = 10'd295;
b_exp0 = 10'd805; b_exp1 = 10'd683; b_exp2 = 10'd206; b_exp3 = 10'd55;
a_sign0 = 4'd11; a_sign1 = 4'd4; a_sign2 = 4'd10; a_sign3 = 4'd2;
b_sign0 = 4'd7; b_sign1 = 4'd9; b_sign2 = 4'd10; b_sign3 = 4'd7;
@(posedge clk_i);
a_mant0 = 8'd99; a_mant1 = 8'd227; a_mant2 = 8'd222; a_mant3 = 8'd4;
b_mant0 = 8'd249; b_mant1 = 8'd217; b_mant2 = 8'd64; b_mant3 = 8'd173;
a_exp0 = 10'd32; a_exp1 = 10'd736; a_exp2 = 10'd191; a_exp3 = 10'd884;
b_exp0 = 10'd957; b_exp1 = 10'd920; b_exp2 = 10'd724; b_exp3 = 10'd986;
a_sign0 = 4'd10; a_sign1 = 4'd0; a_sign2 = 4'd1; a_sign3 = 4'd6;
b_sign0 = 4'd1; b_sign1 = 4'd10; b_sign2 = 4'd6; b_sign3 = 4'd14;
@(posedge clk_i);
a_mant0 = 8'd107; a_mant1 = 8'd86; a_mant2 = 8'd33; a_mant3 = 8'd42;
b_mant0 = 8'd248; b_mant1 = 8'd247; b_mant2 = 8'd20; b_mant3 = 8'd249;
a_exp0 = 10'd582; a_exp1 = 10'd752; a_exp2 = 10'd887; a_exp3 = 10'd8;
b_exp0 = 10'd630; b_exp1 = 10'd913; b_exp2 = 10'd987; b_exp3 = 10'd696;
a_sign0 = 4'd8; a_sign1 = 4'd11; a_sign2 = 4'd6; a_sign3 = 4'd12;
b_sign0 = 4'd7; b_sign1 = 4'd5; b_sign2 = 4'd8; b_sign3 = 4'd16;
@(posedge clk_i);
a_mant0 = 8'd198; a_mant1 = 8'd71; a_mant2 = 8'd32; a_mant3 = 8'd24;
b_mant0 = 8'd224; b_mant1 = 8'd204; b_mant2 = 8'd140; b_mant3 = 8'd70;
a_exp0 = 10'd343; a_exp1 = 10'd743; a_exp2 = 10'd57; a_exp3 = 10'd950;
b_exp0 = 10'd889; b_exp1 = 10'd280; b_exp2 = 10'd873; b_exp3 = 10'd751;
a_sign0 = 4'd14; a_sign1 = 4'd8; a_sign2 = 4'd7; a_sign3 = 4'd7;
b_sign0 = 4'd10; b_sign1 = 4'd12; b_sign2 = 4'd15; b_sign3 = 4'd2;
@(posedge clk_i);
a_mant0 = 8'd228; a_mant1 = 8'd174; a_mant2 = 8'd209; a_mant3 = 8'd190;
b_mant0 = 8'd15; b_mant1 = 8'd96; b_mant2 = 8'd83; b_mant3 = 8'd209;
a_exp0 = 10'd18; a_exp1 = 10'd992; a_exp2 = 10'd580; a_exp3 = 10'd989;
b_exp0 = 10'd661; b_exp1 = 10'd639; b_exp2 = 10'd48; b_exp3 = 10'd418;
a_sign0 = 4'd10; a_sign1 = 4'd10; a_sign2 = 4'd15; a_sign3 = 4'd3;
b_sign0 = 4'd7; b_sign1 = 4'd13; b_sign2 = 4'd2; b_sign3 = 4'd4;
@(posedge clk_i);
a_mant0 = 8'd25; a_mant1 = 8'd121; a_mant2 = 8'd94; a_mant3 = 8'd33;
b_mant0 = 8'd166; b_mant1 = 8'd96; b_mant2 = 8'd136; b_mant3 = 8'd214;
a_exp0 = 10'd858; a_exp1 = 10'd770; a_exp2 = 10'd654; a_exp3 = 10'd984;
b_exp0 = 10'd548; b_exp1 = 10'd101; b_exp2 = 10'd894; b_exp3 = 10'd783;
a_sign0 = 4'd8; a_sign1 = 4'd5; a_sign2 = 4'd7; a_sign3 = 4'd12;
b_sign0 = 4'd13; b_sign1 = 4'd3; b_sign2 = 4'd10; b_sign3 = 4'd7;
@(posedge clk_i);
a_mant0 = 8'd1; a_mant1 = 8'd114; a_mant2 = 8'd121; a_mant3 = 8'd196;
b_mant0 = 8'd43; b_mant1 = 8'd178; b_mant2 = 8'd33; b_mant3 = 8'd12;
a_exp0 = 10'd645; a_exp1 = 10'd346; a_exp2 = 10'd362; a_exp3 = 10'd659;
b_exp0 = 10'd356; b_exp1 = 10'd355; b_exp2 = 10'd0; b_exp3 = 10'd878;
a_sign0 = 4'd11; a_sign1 = 4'd2; a_sign2 = 4'd9; a_sign3 = 4'd2;
b_sign0 = 4'd10; b_sign1 = 4'd13; b_sign2 = 4'd13; b_sign3 = 4'd4;
@(posedge clk_i);
shared_exps0 = 8'd111;
shared_exps1 = 8'd115;
a_mant0 = 8'd196; a_mant1 = 8'd197; a_mant2 = 8'd75; a_mant3 = 8'd181;
b_mant0 = 8'd164; b_mant1 = 8'd109; b_mant2 = 8'd129; b_mant3 = 8'd96;
a_exp0 = 10'd914; a_exp1 = 10'd288; a_exp2 = 10'd279; a_exp3 = 10'd734;
b_exp0 = 10'd850; b_exp1 = 10'd389; b_exp2 = 10'd332; b_exp3 = 10'd297;
a_sign0 = 4'd4; a_sign1 = 4'd7; a_sign2 = 4'd14; a_sign3 = 4'd9;
b_sign0 = 4'd6; b_sign1 = 4'd5; b_sign2 = 4'd2; b_sign3 = 4'd10;
@(posedge clk_i);
a_mant0 = 8'd14; a_mant1 = 8'd83; a_mant2 = 8'd80; a_mant3 = 8'd188;
b_mant0 = 8'd75; b_mant1 = 8'd88; b_mant2 = 8'd18; b_mant3 = 8'd134;
a_exp0 = 10'd163; a_exp1 = 10'd283; a_exp2 = 10'd861; a_exp3 = 10'd888;
b_exp0 = 10'd769; b_exp1 = 10'd335; b_exp2 = 10'd24; b_exp3 = 10'd1000;
a_sign0 = 4'd13; a_sign1 = 4'd2; a_sign2 = 4'd1; a_sign3 = 4'd13;
b_sign0 = 4'd4; b_sign1 = 4'd6; b_sign2 = 4'd5; b_sign3 = 4'd7;
@(posedge clk_i);
a_mant0 = 8'd247; a_mant1 = 8'd218; a_mant2 = 8'd122; a_mant3 = 8'd43;
b_mant0 = 8'd139; b_mant1 = 8'd139; b_mant2 = 8'd112; b_mant3 = 8'd63;
a_exp0 = 10'd403; a_exp1 = 10'd83; a_exp2 = 10'd495; a_exp3 = 10'd968;
b_exp0 = 10'd77; b_exp1 = 10'd839; b_exp2 = 10'd336; b_exp3 = 10'd323;
a_sign0 = 4'd4; a_sign1 = 4'd11; a_sign2 = 4'd13; a_sign3 = 4'd9;
b_sign0 = 4'd12; b_sign1 = 4'd11; b_sign2 = 4'd3; b_sign3 = 4'd16;
@(posedge clk_i);
a_mant0 = 8'd35; a_mant1 = 8'd202; a_mant2 = 8'd159; a_mant3 = 8'd196;
b_mant0 = 8'd242; b_mant1 = 8'd244; b_mant2 = 8'd218; b_mant3 = 8'd111;
a_exp0 = 10'd972; a_exp1 = 10'd576; a_exp2 = 10'd727; a_exp3 = 10'd706;
b_exp0 = 10'd2; b_exp1 = 10'd675; b_exp2 = 10'd372; b_exp3 = 10'd535;
a_sign0 = 4'd14; a_sign1 = 4'd5; a_sign2 = 4'd6; a_sign3 = 4'd1;
b_sign0 = 4'd15; b_sign1 = 4'd8; b_sign2 = 4'd16; b_sign3 = 4'd8;
@(posedge clk_i);
a_mant0 = 8'd69; a_mant1 = 8'd129; a_mant2 = 8'd149; a_mant3 = 8'd241;
b_mant0 = 8'd19; b_mant1 = 8'd54; b_mant2 = 8'd244; b_mant3 = 8'd119;
a_exp0 = 10'd702; a_exp1 = 10'd27; a_exp2 = 10'd648; a_exp3 = 10'd54;
b_exp0 = 10'd507; b_exp1 = 10'd638; b_exp2 = 10'd830; b_exp3 = 10'd767;
a_sign0 = 4'd11; a_sign1 = 4'd9; a_sign2 = 4'd2; a_sign3 = 4'd8;
b_sign0 = 4'd16; b_sign1 = 4'd0; b_sign2 = 4'd2; b_sign3 = 4'd7;
@(posedge clk_i);
a_mant0 = 8'd89; a_mant1 = 8'd3; a_mant2 = 8'd228; a_mant3 = 8'd135;
b_mant0 = 8'd179; b_mant1 = 8'd14; b_mant2 = 8'd213; b_mant3 = 8'd182;
a_exp0 = 10'd928; a_exp1 = 10'd328; a_exp2 = 10'd592; a_exp3 = 10'd378;
b_exp0 = 10'd526; b_exp1 = 10'd619; b_exp2 = 10'd59; b_exp3 = 10'd777;
a_sign0 = 4'd6; a_sign1 = 4'd14; a_sign2 = 4'd0; a_sign3 = 4'd8;
b_sign0 = 4'd1; b_sign1 = 4'd5; b_sign2 = 4'd10; b_sign3 = 4'd8;
@(posedge clk_i);
a_mant0 = 8'd26; a_mant1 = 8'd101; a_mant2 = 8'd220; a_mant3 = 8'd109;
b_mant0 = 8'd20; b_mant1 = 8'd201; b_mant2 = 8'd250; b_mant3 = 8'd188;
a_exp0 = 10'd1003; a_exp1 = 10'd95; a_exp2 = 10'd93; a_exp3 = 10'd746;
b_exp0 = 10'd409; b_exp1 = 10'd253; b_exp2 = 10'd50; b_exp3 = 10'd29;
a_sign0 = 4'd14; a_sign1 = 4'd5; a_sign2 = 4'd15; a_sign3 = 4'd16;
b_sign0 = 4'd16; b_sign1 = 4'd2; b_sign2 = 4'd1; b_sign3 = 4'd8;
@(posedge clk_i);
a_mant0 = 8'd42; a_mant1 = 8'd160; a_mant2 = 8'd133; a_mant3 = 8'd47;
b_mant0 = 8'd84; b_mant1 = 8'd228; b_mant2 = 8'd181; b_mant3 = 8'd15;
a_exp0 = 10'd128; a_exp1 = 10'd542; a_exp2 = 10'd98; a_exp3 = 10'd475;
b_exp0 = 10'd807; b_exp1 = 10'd665; b_exp2 = 10'd733; b_exp3 = 10'd276;
a_sign0 = 4'd14; a_sign1 = 4'd16; a_sign2 = 4'd7; a_sign3 = 4'd5;
b_sign0 = 4'd11; b_sign1 = 4'd9; b_sign2 = 4'd2; b_sign3 = 4'd14;
@(posedge clk_i);
shared_exps0 = 8'd141;
shared_exps1 = 8'd133;
rstn = 0;
@(posedge clk_i);
rstn = 1;
a_mant0 = 8'd251; a_mant1 = 8'd203; a_mant2 = 8'd248; a_mant3 = 8'd169;
b_mant0 = 8'd143; b_mant1 = 8'd234; b_mant2 = 8'd84; b_mant3 = 8'd126;
a_exp0 = 10'd107; a_exp1 = 10'd890; a_exp2 = 10'd645; a_exp3 = 10'd908;
b_exp0 = 10'd859; b_exp1 = 10'd697; b_exp2 = 10'd630; b_exp3 = 10'd484;
a_sign0 = 4'd16; a_sign1 = 4'd5; a_sign2 = 4'd8; a_sign3 = 4'd15;
b_sign0 = 4'd3; b_sign1 = 4'd5; b_sign2 = 4'd7; b_sign3 = 4'd8;
@(posedge clk_i);
a_mant0 = 8'd250; a_mant1 = 8'd106; a_mant2 = 8'd146; a_mant3 = 8'd111;
b_mant0 = 8'd45; b_mant1 = 8'd62; b_mant2 = 8'd183; b_mant3 = 8'd94;
a_exp0 = 10'd197; a_exp1 = 10'd418; a_exp2 = 10'd358; a_exp3 = 10'd668;
b_exp0 = 10'd155; b_exp1 = 10'd345; b_exp2 = 10'd533; b_exp3 = 10'd314;
a_sign0 = 4'd0; a_sign1 = 4'd16; a_sign2 = 4'd14; a_sign3 = 4'd10;
b_sign0 = 4'd15; b_sign1 = 4'd0; b_sign2 = 4'd0; b_sign3 = 4'd16;
@(posedge clk_i);
a_mant0 = 8'd69; a_mant1 = 8'd103; a_mant2 = 8'd94; a_mant3 = 8'd62;
b_mant0 = 8'd179; b_mant1 = 8'd198; b_mant2 = 8'd175; b_mant3 = 8'd15;
a_exp0 = 10'd728; a_exp1 = 10'd296; a_exp2 = 10'd155; a_exp3 = 10'd841;
b_exp0 = 10'd261; b_exp1 = 10'd710; b_exp2 = 10'd613; b_exp3 = 10'd295;
a_sign0 = 4'd2; a_sign1 = 4'd13; a_sign2 = 4'd5; a_sign3 = 4'd12;
b_sign0 = 4'd4; b_sign1 = 4'd6; b_sign2 = 4'd9; b_sign3 = 4'd11;
@(posedge clk_i);
a_mant0 = 8'd126; a_mant1 = 8'd205; a_mant2 = 8'd195; a_mant3 = 8'd37;
b_mant0 = 8'd96; b_mant1 = 8'd136; b_mant2 = 8'd55; b_mant3 = 8'd132;
a_exp0 = 10'd8; a_exp1 = 10'd998; a_exp2 = 10'd65; a_exp3 = 10'd779;
b_exp0 = 10'd231; b_exp1 = 10'd3; b_exp2 = 10'd885; b_exp3 = 10'd63;
a_sign0 = 4'd12; a_sign1 = 4'd9; a_sign2 = 4'd8; a_sign3 = 4'd10;
b_sign0 = 4'd4; b_sign1 = 4'd1; b_sign2 = 4'd4; b_sign3 = 4'd10;
@(posedge clk_i);
a_mant0 = 8'd106; a_mant1 = 8'd131; a_mant2 = 8'd85; a_mant3 = 8'd225;
b_mant0 = 8'd133; b_mant1 = 8'd18; b_mant2 = 8'd216; b_mant3 = 8'd213;
a_exp0 = 10'd913; a_exp1 = 10'd314; a_exp2 = 10'd725; a_exp3 = 10'd495;
b_exp0 = 10'd762; b_exp1 = 10'd645; b_exp2 = 10'd956; b_exp3 = 10'd740;
a_sign0 = 4'd5; a_sign1 = 4'd8; a_sign2 = 4'd13; a_sign3 = 4'd11;
b_sign0 = 4'd8; b_sign1 = 4'd16; b_sign2 = 4'd10; b_sign3 = 4'd0;
@(posedge clk_i);
a_mant0 = 8'd109; a_mant1 = 8'd222; a_mant2 = 8'd116; a_mant3 = 8'd196;
b_mant0 = 8'd12; b_mant1 = 8'd104; b_mant2 = 8'd143; b_mant3 = 8'd148;
a_exp0 = 10'd452; a_exp1 = 10'd773; a_exp2 = 10'd394; a_exp3 = 10'd471;
b_exp0 = 10'd475; b_exp1 = 10'd873; b_exp2 = 10'd912; b_exp3 = 10'd433;
a_sign0 = 4'd5; a_sign1 = 4'd0; a_sign2 = 4'd1; a_sign3 = 4'd6;
b_sign0 = 4'd15; b_sign1 = 4'd2; b_sign2 = 4'd4; b_sign3 = 4'd10;
@(posedge clk_i);
a_mant0 = 8'd181; a_mant1 = 8'd239; a_mant2 = 8'd175; a_mant3 = 8'd30;
b_mant0 = 8'd245; b_mant1 = 8'd81; b_mant2 = 8'd246; b_mant3 = 8'd139;
a_exp0 = 10'd799; a_exp1 = 10'd269; a_exp2 = 10'd668; a_exp3 = 10'd825;
b_exp0 = 10'd935; b_exp1 = 10'd673; b_exp2 = 10'd1015; b_exp3 = 10'd554;
a_sign0 = 4'd11; a_sign1 = 4'd6; a_sign2 = 4'd7; a_sign3 = 4'd11;
b_sign0 = 4'd11; b_sign1 = 4'd11; b_sign2 = 4'd2; b_sign3 = 4'd16;
@(posedge clk_i);
shared_exps0 = 8'd122;
shared_exps1 = 8'd144;
a_mant0 = 8'd165; a_mant1 = 8'd199; a_mant2 = 8'd29; a_mant3 = 8'd89;
b_mant0 = 8'd74; b_mant1 = 8'd207; b_mant2 = 8'd235; b_mant3 = 8'd186;
a_exp0 = 10'd459; a_exp1 = 10'd351; a_exp2 = 10'd453; a_exp3 = 10'd274;
b_exp0 = 10'd156; b_exp1 = 10'd191; b_exp2 = 10'd1023; b_exp3 = 10'd654;
a_sign0 = 4'd5; a_sign1 = 4'd16; a_sign2 = 4'd11; a_sign3 = 4'd16;
b_sign0 = 4'd5; b_sign1 = 4'd8; b_sign2 = 4'd8; b_sign3 = 4'd14;
@(posedge clk_i);
a_mant0 = 8'd153; a_mant1 = 8'd197; a_mant2 = 8'd168; a_mant3 = 8'd157;
b_mant0 = 8'd200; b_mant1 = 8'd29; b_mant2 = 8'd219; b_mant3 = 8'd162;
a_exp0 = 10'd983; a_exp1 = 10'd17; a_exp2 = 10'd942; a_exp3 = 10'd143;
b_exp0 = 10'd938; b_exp1 = 10'd175; b_exp2 = 10'd888; b_exp3 = 10'd43;
a_sign0 = 4'd8; a_sign1 = 4'd10; a_sign2 = 4'd5; a_sign3 = 4'd0;
b_sign0 = 4'd8; b_sign1 = 4'd5; b_sign2 = 4'd16; b_sign3 = 4'd2;
@(posedge clk_i);
a_mant0 = 8'd137; a_mant1 = 8'd13; a_mant2 = 8'd212; a_mant3 = 8'd103;
b_mant0 = 8'd52; b_mant1 = 8'd16; b_mant2 = 8'd60; b_mant3 = 8'd183;
a_exp0 = 10'd1010; a_exp1 = 10'd117; a_exp2 = 10'd981; a_exp3 = 10'd82;
b_exp0 = 10'd894; b_exp1 = 10'd860; b_exp2 = 10'd708; b_exp3 = 10'd181;
a_sign0 = 4'd11; a_sign1 = 4'd7; a_sign2 = 4'd7; a_sign3 = 4'd9;
b_sign0 = 4'd4; b_sign1 = 4'd3; b_sign2 = 4'd1; b_sign3 = 4'd4;
@(posedge clk_i);
a_mant0 = 8'd16; a_mant1 = 8'd9; a_mant2 = 8'd223; a_mant3 = 8'd112;
b_mant0 = 8'd62; b_mant1 = 8'd242; b_mant2 = 8'd219; b_mant3 = 8'd161;
a_exp0 = 10'd558; a_exp1 = 10'd215; a_exp2 = 10'd226; a_exp3 = 10'd33;
b_exp0 = 10'd563; b_exp1 = 10'd779; b_exp2 = 10'd659; b_exp3 = 10'd682;
a_sign0 = 4'd1; a_sign1 = 4'd4; a_sign2 = 4'd11; a_sign3 = 4'd9;
b_sign0 = 4'd9; b_sign1 = 4'd16; b_sign2 = 4'd2; b_sign3 = 4'd7;
@(posedge clk_i);
a_mant0 = 8'd242; a_mant1 = 8'd107; a_mant2 = 8'd171; a_mant3 = 8'd99;
b_mant0 = 8'd144; b_mant1 = 8'd229; b_mant2 = 8'd188; b_mant3 = 8'd215;
a_exp0 = 10'd318; a_exp1 = 10'd676; a_exp2 = 10'd760; a_exp3 = 10'd207;
b_exp0 = 10'd459; b_exp1 = 10'd221; b_exp2 = 10'd865; b_exp3 = 10'd357;
a_sign0 = 4'd9; a_sign1 = 4'd4; a_sign2 = 4'd2; a_sign3 = 4'd1;
b_sign0 = 4'd12; b_sign1 = 4'd9; b_sign2 = 4'd7; b_sign3 = 4'd11;
@(posedge clk_i);
a_mant0 = 8'd38; a_mant1 = 8'd20; a_mant2 = 8'd222; a_mant3 = 8'd127;
b_mant0 = 8'd58; b_mant1 = 8'd187; b_mant2 = 8'd48; b_mant3 = 8'd85;
a_exp0 = 10'd20; a_exp1 = 10'd841; a_exp2 = 10'd545; a_exp3 = 10'd208;
b_exp0 = 10'd924; b_exp1 = 10'd626; b_exp2 = 10'd864; b_exp3 = 10'd257;
a_sign0 = 4'd5; a_sign1 = 4'd1; a_sign2 = 4'd4; a_sign3 = 4'd16;
b_sign0 = 4'd6; b_sign1 = 4'd2; b_sign2 = 4'd16; b_sign3 = 4'd1;
@(posedge clk_i);
a_mant0 = 8'd209; a_mant1 = 8'd244; a_mant2 = 8'd97; a_mant3 = 8'd9;
b_mant0 = 8'd54; b_mant1 = 8'd4; b_mant2 = 8'd132; b_mant3 = 8'd115;
a_exp0 = 10'd236; a_exp1 = 10'd473; a_exp2 = 10'd594; a_exp3 = 10'd869;
b_exp0 = 10'd320; b_exp1 = 10'd235; b_exp2 = 10'd645; b_exp3 = 10'd780;
a_sign0 = 4'd12; a_sign1 = 4'd7; a_sign2 = 4'd6; a_sign3 = 4'd15;
b_sign0 = 4'd9; b_sign1 = 4'd6; b_sign2 = 4'd4; b_sign3 = 4'd10;
@(posedge clk_i);
a_mant0 = 8'd32; a_mant1 = 8'd115; a_mant2 = 8'd140; a_mant3 = 8'd254;
b_mant0 = 8'd135; b_mant1 = 8'd56; b_mant2 = 8'd8; b_mant3 = 8'd111;
a_exp0 = 10'd84; a_exp1 = 10'd447; a_exp2 = 10'd402; a_exp3 = 10'd308;
b_exp0 = 10'd877; b_exp1 = 10'd1023; b_exp2 = 10'd684; b_exp3 = 10'd872;
a_sign0 = 4'd12; a_sign1 = 4'd9; a_sign2 = 4'd4; a_sign3 = 4'd5;
b_sign0 = 4'd7; b_sign1 = 4'd1; b_sign2 = 4'd8; b_sign3 = 4'd15;
@(posedge clk_i);
shared_exps0 = 8'd135;
shared_exps1 = 8'd141;
a_mant0 = 8'd179; a_mant1 = 8'd4; a_mant2 = 8'd145; a_mant3 = 8'd177;
b_mant0 = 8'd185; b_mant1 = 8'd86; b_mant2 = 8'd168; b_mant3 = 8'd215;
a_exp0 = 10'd4; a_exp1 = 10'd899; a_exp2 = 10'd755; a_exp3 = 10'd623;
b_exp0 = 10'd434; b_exp1 = 10'd457; b_exp2 = 10'd890; b_exp3 = 10'd921;
a_sign0 = 4'd12; a_sign1 = 4'd11; a_sign2 = 4'd14; a_sign3 = 4'd5;
b_sign0 = 4'd14; b_sign1 = 4'd3; b_sign2 = 4'd2; b_sign3 = 4'd5;
@(posedge clk_i);
a_mant0 = 8'd105; a_mant1 = 8'd60; a_mant2 = 8'd235; a_mant3 = 8'd13;
b_mant0 = 8'd118; b_mant1 = 8'd10; b_mant2 = 8'd158; b_mant3 = 8'd29;
a_exp0 = 10'd929; a_exp1 = 10'd195; a_exp2 = 10'd8; a_exp3 = 10'd488;
b_exp0 = 10'd932; b_exp1 = 10'd643; b_exp2 = 10'd1010; b_exp3 = 10'd245;
a_sign0 = 4'd9; a_sign1 = 4'd14; a_sign2 = 4'd2; a_sign3 = 4'd16;
b_sign0 = 4'd1; b_sign1 = 4'd0; b_sign2 = 4'd8; b_sign3 = 4'd3;
@(posedge clk_i);
a_mant0 = 8'd37; a_mant1 = 8'd67; a_mant2 = 8'd201; a_mant3 = 8'd184;
b_mant0 = 8'd147; b_mant1 = 8'd87; b_mant2 = 8'd229; b_mant3 = 8'd213;
a_exp0 = 10'd765; a_exp1 = 10'd337; a_exp2 = 10'd356; a_exp3 = 10'd935;
b_exp0 = 10'd871; b_exp1 = 10'd1019; b_exp2 = 10'd336; b_exp3 = 10'd131;
a_sign0 = 4'd0; a_sign1 = 4'd12; a_sign2 = 4'd5; a_sign3 = 4'd11;
b_sign0 = 4'd8; b_sign1 = 4'd13; b_sign2 = 4'd9; b_sign3 = 4'd6;
@(posedge clk_i);
a_mant0 = 8'd194; a_mant1 = 8'd47; a_mant2 = 8'd61; a_mant3 = 8'd34;
b_mant0 = 8'd47; b_mant1 = 8'd165; b_mant2 = 8'd44; b_mant3 = 8'd240;
a_exp0 = 10'd268; a_exp1 = 10'd678; a_exp2 = 10'd235; a_exp3 = 10'd385;
b_exp0 = 10'd26; b_exp1 = 10'd16; b_exp2 = 10'd926; b_exp3 = 10'd558;
a_sign0 = 4'd10; a_sign1 = 4'd2; a_sign2 = 4'd7; a_sign3 = 4'd7;
b_sign0 = 4'd10; b_sign1 = 4'd6; b_sign2 = 4'd8; b_sign3 = 4'd16;
@(posedge clk_i);
a_mant0 = 8'd107; a_mant1 = 8'd0; a_mant2 = 8'd72; a_mant3 = 8'd47;
b_mant0 = 8'd224; b_mant1 = 8'd71; b_mant2 = 8'd154; b_mant3 = 8'd24;
a_exp0 = 10'd233; a_exp1 = 10'd241; a_exp2 = 10'd598; a_exp3 = 10'd358;
b_exp0 = 10'd661; b_exp1 = 10'd990; b_exp2 = 10'd52; b_exp3 = 10'd1009;
a_sign0 = 4'd8; a_sign1 = 4'd14; a_sign2 = 4'd4; a_sign3 = 4'd10;
b_sign0 = 4'd13; b_sign1 = 4'd1; b_sign2 = 4'd8; b_sign3 = 4'd8;
@(posedge clk_i);
a_mant0 = 8'd222; a_mant1 = 8'd18; a_mant2 = 8'd61; a_mant3 = 8'd111;
b_mant0 = 8'd107; b_mant1 = 8'd231; b_mant2 = 8'd131; b_mant3 = 8'd134;
a_exp0 = 10'd142; a_exp1 = 10'd878; a_exp2 = 10'd52; a_exp3 = 10'd553;
b_exp0 = 10'd412; b_exp1 = 10'd540; b_exp2 = 10'd898; b_exp3 = 10'd76;
a_sign0 = 4'd3; a_sign1 = 4'd12; a_sign2 = 4'd13; a_sign3 = 4'd14;
b_sign0 = 4'd15; b_sign1 = 4'd1; b_sign2 = 4'd10; b_sign3 = 4'd4;
@(posedge clk_i);
a_mant0 = 8'd86; a_mant1 = 8'd215; a_mant2 = 8'd55; a_mant3 = 8'd245;
b_mant0 = 8'd148; b_mant1 = 8'd191; b_mant2 = 8'd19; b_mant3 = 8'd7;
a_exp0 = 10'd116; a_exp1 = 10'd137; a_exp2 = 10'd813; a_exp3 = 10'd1004;
b_exp0 = 10'd877; b_exp1 = 10'd392; b_exp2 = 10'd763; b_exp3 = 10'd444;
a_sign0 = 4'd3; a_sign1 = 4'd8; a_sign2 = 4'd11; a_sign3 = 4'd9;
b_sign0 = 4'd8; b_sign1 = 4'd15; b_sign2 = 4'd8; b_sign3 = 4'd8;
@(posedge clk_i);
a_mant0 = 8'd124; a_mant1 = 8'd67; a_mant2 = 8'd206; a_mant3 = 8'd76;
b_mant0 = 8'd130; b_mant1 = 8'd104; b_mant2 = 8'd140; b_mant3 = 8'd64;
a_exp0 = 10'd990; a_exp1 = 10'd261; a_exp2 = 10'd684; a_exp3 = 10'd102;
b_exp0 = 10'd136; b_exp1 = 10'd35; b_exp2 = 10'd228; b_exp3 = 10'd678;
a_sign0 = 4'd8; a_sign1 = 4'd16; a_sign2 = 4'd6; a_sign3 = 4'd14;
b_sign0 = 4'd13; b_sign1 = 4'd10; b_sign2 = 4'd13; b_sign3 = 4'd12;
@(posedge clk_i);
shared_exps0 = 8'd151;
shared_exps1 = 8'd156;
a_mant0 = 8'd12; a_mant1 = 8'd11; a_mant2 = 8'd84; a_mant3 = 8'd172;
b_mant0 = 8'd60; b_mant1 = 8'd172; b_mant2 = 8'd1; b_mant3 = 8'd157;
a_exp0 = 10'd154; a_exp1 = 10'd636; a_exp2 = 10'd517; a_exp3 = 10'd50;
b_exp0 = 10'd962; b_exp1 = 10'd486; b_exp2 = 10'd281; b_exp3 = 10'd954;
a_sign0 = 4'd7; a_sign1 = 4'd2; a_sign2 = 4'd8; a_sign3 = 4'd10;
b_sign0 = 4'd6; b_sign1 = 4'd5; b_sign2 = 4'd4; b_sign3 = 4'd16;
@(posedge clk_i);
a_mant0 = 8'd138; a_mant1 = 8'd98; a_mant2 = 8'd59; a_mant3 = 8'd67;
b_mant0 = 8'd230; b_mant1 = 8'd81; b_mant2 = 8'd92; b_mant3 = 8'd47;
a_exp0 = 10'd913; a_exp1 = 10'd384; a_exp2 = 10'd893; a_exp3 = 10'd714;
b_exp0 = 10'd178; b_exp1 = 10'd102; b_exp2 = 10'd732; b_exp3 = 10'd311;
a_sign0 = 4'd2; a_sign1 = 4'd2; a_sign2 = 4'd2; a_sign3 = 4'd1;
b_sign0 = 4'd11; b_sign1 = 4'd9; b_sign2 = 4'd14; b_sign3 = 4'd15;
@(posedge clk_i);
a_mant0 = 8'd209; a_mant1 = 8'd199; a_mant2 = 8'd19; a_mant3 = 8'd16;
b_mant0 = 8'd118; b_mant1 = 8'd10; b_mant2 = 8'd222; b_mant3 = 8'd30;
a_exp0 = 10'd296; a_exp1 = 10'd109; a_exp2 = 10'd647; a_exp3 = 10'd1018;
b_exp0 = 10'd144; b_exp1 = 10'd323; b_exp2 = 10'd466; b_exp3 = 10'd819;
a_sign0 = 4'd4; a_sign1 = 4'd9; a_sign2 = 4'd9; a_sign3 = 4'd7;
b_sign0 = 4'd4; b_sign1 = 4'd0; b_sign2 = 4'd2; b_sign3 = 4'd6;
@(posedge clk_i);
a_mant0 = 8'd44; a_mant1 = 8'd221; a_mant2 = 8'd170; a_mant3 = 8'd72;
b_mant0 = 8'd82; b_mant1 = 8'd239; b_mant2 = 8'd123; b_mant3 = 8'd55;
a_exp0 = 10'd798; a_exp1 = 10'd176; a_exp2 = 10'd877; a_exp3 = 10'd845;
b_exp0 = 10'd376; b_exp1 = 10'd923; b_exp2 = 10'd815; b_exp3 = 10'd655;
a_sign0 = 4'd11; a_sign1 = 4'd11; a_sign2 = 4'd0; a_sign3 = 4'd0;
b_sign0 = 4'd10; b_sign1 = 4'd4; b_sign2 = 4'd14; b_sign3 = 4'd12;
@(posedge clk_i);
a_mant0 = 8'd108; a_mant1 = 8'd72; a_mant2 = 8'd205; a_mant3 = 8'd141;
b_mant0 = 8'd215; b_mant1 = 8'd7; b_mant2 = 8'd136; b_mant3 = 8'd135;
a_exp0 = 10'd971; a_exp1 = 10'd1017; a_exp2 = 10'd150; a_exp3 = 10'd258;
b_exp0 = 10'd12; b_exp1 = 10'd928; b_exp2 = 10'd138; b_exp3 = 10'd580;
a_sign0 = 4'd10; a_sign1 = 4'd16; a_sign2 = 4'd6; a_sign3 = 4'd9;
b_sign0 = 4'd10; b_sign1 = 4'd7; b_sign2 = 4'd11; b_sign3 = 4'd7;
@(posedge clk_i);
a_mant0 = 8'd8; a_mant1 = 8'd180; a_mant2 = 8'd13; a_mant3 = 8'd82;
b_mant0 = 8'd6; b_mant1 = 8'd198; b_mant2 = 8'd161; b_mant3 = 8'd150;
a_exp0 = 10'd391; a_exp1 = 10'd406; a_exp2 = 10'd740; a_exp3 = 10'd704;
b_exp0 = 10'd63; b_exp1 = 10'd587; b_exp2 = 10'd590; b_exp3 = 10'd762;
a_sign0 = 4'd1; a_sign1 = 4'd8; a_sign2 = 4'd8; a_sign3 = 4'd10;
b_sign0 = 4'd2; b_sign1 = 4'd1; b_sign2 = 4'd3; b_sign3 = 4'd11;
@(posedge clk_i);
a_mant0 = 8'd126; a_mant1 = 8'd17; a_mant2 = 8'd57; a_mant3 = 8'd87;
b_mant0 = 8'd125; b_mant1 = 8'd198; b_mant2 = 8'd122; b_mant3 = 8'd21;
a_exp0 = 10'd914; a_exp1 = 10'd607; a_exp2 = 10'd221; a_exp3 = 10'd747;
b_exp0 = 10'd499; b_exp1 = 10'd572; b_exp2 = 10'd201; b_exp3 = 10'd908;
a_sign0 = 4'd16; a_sign1 = 4'd14; a_sign2 = 4'd10; a_sign3 = 4'd16;
b_sign0 = 4'd4; b_sign1 = 4'd6; b_sign2 = 4'd10; b_sign3 = 4'd15;
@(posedge clk_i);
a_mant0 = 8'd119; a_mant1 = 8'd53; a_mant2 = 8'd74; a_mant3 = 8'd10;
b_mant0 = 8'd84; b_mant1 = 8'd132; b_mant2 = 8'd116; b_mant3 = 8'd156;
a_exp0 = 10'd984; a_exp1 = 10'd15; a_exp2 = 10'd725; a_exp3 = 10'd369;
b_exp0 = 10'd225; b_exp1 = 10'd771; b_exp2 = 10'd985; b_exp3 = 10'd201;
a_sign0 = 4'd11; a_sign1 = 4'd12; a_sign2 = 4'd10; a_sign3 = 4'd16;
b_sign0 = 4'd14; b_sign1 = 4'd12; b_sign2 = 4'd11; b_sign3 = 4'd0;
@(posedge clk_i);
shared_exps0 = 8'd84;
shared_exps1 = 8'd143;
rstn = 0;
@(posedge clk_i);
rstn = 1;
a_mant0 = 8'd142; a_mant1 = 8'd151; a_mant2 = 8'd11; a_mant3 = 8'd162;
b_mant0 = 8'd134; b_mant1 = 8'd100; b_mant2 = 8'd92; b_mant3 = 8'd221;
a_exp0 = 10'd541; a_exp1 = 10'd143; a_exp2 = 10'd746; a_exp3 = 10'd806;
b_exp0 = 10'd434; b_exp1 = 10'd109; b_exp2 = 10'd175; b_exp3 = 10'd108;
a_sign0 = 4'd9; a_sign1 = 4'd6; a_sign2 = 4'd9; a_sign3 = 4'd12;
b_sign0 = 4'd13; b_sign1 = 4'd1; b_sign2 = 4'd9; b_sign3 = 4'd4;
@(posedge clk_i);
a_mant0 = 8'd111; a_mant1 = 8'd87; a_mant2 = 8'd92; a_mant3 = 8'd112;
b_mant0 = 8'd98; b_mant1 = 8'd77; b_mant2 = 8'd205; b_mant3 = 8'd97;
a_exp0 = 10'd511; a_exp1 = 10'd20; a_exp2 = 10'd804; a_exp3 = 10'd114;
b_exp0 = 10'd623; b_exp1 = 10'd798; b_exp2 = 10'd171; b_exp3 = 10'd996;
a_sign0 = 4'd0; a_sign1 = 4'd13; a_sign2 = 4'd9; a_sign3 = 4'd11;
b_sign0 = 4'd9; b_sign1 = 4'd7; b_sign2 = 4'd0; b_sign3 = 4'd3;
@(posedge clk_i);
a_mant0 = 8'd215; a_mant1 = 8'd148; a_mant2 = 8'd189; a_mant3 = 8'd64;
b_mant0 = 8'd67; b_mant1 = 8'd4; b_mant2 = 8'd39; b_mant3 = 8'd250;
a_exp0 = 10'd535; a_exp1 = 10'd509; a_exp2 = 10'd743; a_exp3 = 10'd873;
b_exp0 = 10'd162; b_exp1 = 10'd50; b_exp2 = 10'd366; b_exp3 = 10'd116;
a_sign0 = 4'd9; a_sign1 = 4'd12; a_sign2 = 4'd5; a_sign3 = 4'd15;
b_sign0 = 4'd16; b_sign1 = 4'd16; b_sign2 = 4'd2; b_sign3 = 4'd8;
@(posedge clk_i);
a_mant0 = 8'd129; a_mant1 = 8'd116; a_mant2 = 8'd103; a_mant3 = 8'd124;
b_mant0 = 8'd16; b_mant1 = 8'd112; b_mant2 = 8'd104; b_mant3 = 8'd248;
a_exp0 = 10'd761; a_exp1 = 10'd356; a_exp2 = 10'd298; a_exp3 = 10'd375;
b_exp0 = 10'd883; b_exp1 = 10'd925; b_exp2 = 10'd450; b_exp3 = 10'd367;
a_sign0 = 4'd14; a_sign1 = 4'd0; a_sign2 = 4'd1; a_sign3 = 4'd14;
b_sign0 = 4'd0; b_sign1 = 4'd9; b_sign2 = 4'd8; b_sign3 = 4'd12;
@(posedge clk_i);
a_mant0 = 8'd118; a_mant1 = 8'd50; a_mant2 = 8'd27; a_mant3 = 8'd251;
b_mant0 = 8'd77; b_mant1 = 8'd120; b_mant2 = 8'd20; b_mant3 = 8'd105;
a_exp0 = 10'd322; a_exp1 = 10'd416; a_exp2 = 10'd713; a_exp3 = 10'd820;
b_exp0 = 10'd482; b_exp1 = 10'd830; b_exp2 = 10'd161; b_exp3 = 10'd846;
a_sign0 = 4'd5; a_sign1 = 4'd14; a_sign2 = 4'd8; a_sign3 = 4'd15;
b_sign0 = 4'd16; b_sign1 = 4'd14; b_sign2 = 4'd2; b_sign3 = 4'd0;
@(posedge clk_i);
a_mant0 = 8'd194; a_mant1 = 8'd76; a_mant2 = 8'd69; a_mant3 = 8'd239;
b_mant0 = 8'd215; b_mant1 = 8'd208; b_mant2 = 8'd97; b_mant3 = 8'd180;
a_exp0 = 10'd413; a_exp1 = 10'd996; a_exp2 = 10'd592; a_exp3 = 10'd610;
b_exp0 = 10'd952; b_exp1 = 10'd708; b_exp2 = 10'd892; b_exp3 = 10'd282;
a_sign0 = 4'd0; a_sign1 = 4'd7; a_sign2 = 4'd3; a_sign3 = 4'd6;
b_sign0 = 4'd11; b_sign1 = 4'd13; b_sign2 = 4'd9; b_sign3 = 4'd16;
@(posedge clk_i);
a_mant0 = 8'd167; a_mant1 = 8'd82; a_mant2 = 8'd1; a_mant3 = 8'd89;
b_mant0 = 8'd251; b_mant1 = 8'd90; b_mant2 = 8'd51; b_mant3 = 8'd18;
a_exp0 = 10'd235; a_exp1 = 10'd130; a_exp2 = 10'd322; a_exp3 = 10'd260;
b_exp0 = 10'd244; b_exp1 = 10'd187; b_exp2 = 10'd336; b_exp3 = 10'd955;
a_sign0 = 4'd9; a_sign1 = 4'd12; a_sign2 = 4'd16; a_sign3 = 4'd15;
b_sign0 = 4'd7; b_sign1 = 4'd3; b_sign2 = 4'd11; b_sign3 = 4'd16;
@(posedge clk_i);
shared_exps0 = 8'd120;
shared_exps1 = 8'd155;
a_mant0 = 8'd124; a_mant1 = 8'd230; a_mant2 = 8'd228; a_mant3 = 8'd139;
b_mant0 = 8'd61; b_mant1 = 8'd132; b_mant2 = 8'd253; b_mant3 = 8'd179;
a_exp0 = 10'd484; a_exp1 = 10'd798; a_exp2 = 10'd672; a_exp3 = 10'd325;
b_exp0 = 10'd714; b_exp1 = 10'd508; b_exp2 = 10'd310; b_exp3 = 10'd1001;
a_sign0 = 4'd9; a_sign1 = 4'd6; a_sign2 = 4'd4; a_sign3 = 4'd2;
b_sign0 = 4'd6; b_sign1 = 4'd14; b_sign2 = 4'd9; b_sign3 = 4'd12;
@(posedge clk_i);
a_mant0 = 8'd230; a_mant1 = 8'd40; a_mant2 = 8'd16; a_mant3 = 8'd103;
b_mant0 = 8'd77; b_mant1 = 8'd133; b_mant2 = 8'd143; b_mant3 = 8'd54;
a_exp0 = 10'd243; a_exp1 = 10'd407; a_exp2 = 10'd875; a_exp3 = 10'd789;
b_exp0 = 10'd797; b_exp1 = 10'd996; b_exp2 = 10'd61; b_exp3 = 10'd378;
a_sign0 = 4'd10; a_sign1 = 4'd2; a_sign2 = 4'd6; a_sign3 = 4'd13;
b_sign0 = 4'd2; b_sign1 = 4'd10; b_sign2 = 4'd8; b_sign3 = 4'd9;
@(posedge clk_i);
a_mant0 = 8'd103; a_mant1 = 8'd139; a_mant2 = 8'd0; a_mant3 = 8'd60;
b_mant0 = 8'd219; b_mant1 = 8'd202; b_mant2 = 8'd60; b_mant3 = 8'd186;
a_exp0 = 10'd711; a_exp1 = 10'd199; a_exp2 = 10'd703; a_exp3 = 10'd935;
b_exp0 = 10'd662; b_exp1 = 10'd450; b_exp2 = 10'd603; b_exp3 = 10'd972;
a_sign0 = 4'd0; a_sign1 = 4'd14; a_sign2 = 4'd11; a_sign3 = 4'd13;
b_sign0 = 4'd11; b_sign1 = 4'd8; b_sign2 = 4'd9; b_sign3 = 4'd7;
@(posedge clk_i);
a_mant0 = 8'd215; a_mant1 = 8'd220; a_mant2 = 8'd77; a_mant3 = 8'd39;
b_mant0 = 8'd53; b_mant1 = 8'd27; b_mant2 = 8'd23; b_mant3 = 8'd228;
a_exp0 = 10'd744; a_exp1 = 10'd328; a_exp2 = 10'd1013; a_exp3 = 10'd146;
b_exp0 = 10'd1013; b_exp1 = 10'd736; b_exp2 = 10'd38; b_exp3 = 10'd525;
a_sign0 = 4'd1; a_sign1 = 4'd15; a_sign2 = 4'd5; a_sign3 = 4'd11;
b_sign0 = 4'd15; b_sign1 = 4'd8; b_sign2 = 4'd1; b_sign3 = 4'd15;
@(posedge clk_i);
a_mant0 = 8'd19; a_mant1 = 8'd182; a_mant2 = 8'd108; a_mant3 = 8'd179;
b_mant0 = 8'd203; b_mant1 = 8'd44; b_mant2 = 8'd228; b_mant3 = 8'd120;
a_exp0 = 10'd795; a_exp1 = 10'd348; a_exp2 = 10'd527; a_exp3 = 10'd907;
b_exp0 = 10'd411; b_exp1 = 10'd708; b_exp2 = 10'd190; b_exp3 = 10'd858;
a_sign0 = 4'd0; a_sign1 = 4'd5; a_sign2 = 4'd7; a_sign3 = 4'd10;
b_sign0 = 4'd7; b_sign1 = 4'd5; b_sign2 = 4'd10; b_sign3 = 4'd3;
@(posedge clk_i);
a_mant0 = 8'd229; a_mant1 = 8'd54; a_mant2 = 8'd29; a_mant3 = 8'd162;
b_mant0 = 8'd7; b_mant1 = 8'd35; b_mant2 = 8'd222; b_mant3 = 8'd225;
a_exp0 = 10'd473; a_exp1 = 10'd273; a_exp2 = 10'd7; a_exp3 = 10'd489;
b_exp0 = 10'd170; b_exp1 = 10'd153; b_exp2 = 10'd1009; b_exp3 = 10'd1020;
a_sign0 = 4'd2; a_sign1 = 4'd10; a_sign2 = 4'd1; a_sign3 = 4'd15;
b_sign0 = 4'd15; b_sign1 = 4'd4; b_sign2 = 4'd11; b_sign3 = 4'd5;
@(posedge clk_i);
a_mant0 = 8'd115; a_mant1 = 8'd104; a_mant2 = 8'd24; a_mant3 = 8'd167;
b_mant0 = 8'd140; b_mant1 = 8'd88; b_mant2 = 8'd178; b_mant3 = 8'd137;
a_exp0 = 10'd1003; a_exp1 = 10'd240; a_exp2 = 10'd48; a_exp3 = 10'd949;
b_exp0 = 10'd126; b_exp1 = 10'd631; b_exp2 = 10'd858; b_exp3 = 10'd351;
a_sign0 = 4'd10; a_sign1 = 4'd11; a_sign2 = 4'd6; a_sign3 = 4'd15;
b_sign0 = 4'd2; b_sign1 = 4'd5; b_sign2 = 4'd3; b_sign3 = 4'd15;
@(posedge clk_i);
a_mant0 = 8'd35; a_mant1 = 8'd20; a_mant2 = 8'd143; a_mant3 = 8'd113;
b_mant0 = 8'd23; b_mant1 = 8'd4; b_mant2 = 8'd155; b_mant3 = 8'd189;
a_exp0 = 10'd1014; a_exp1 = 10'd458; a_exp2 = 10'd1022; a_exp3 = 10'd993;
b_exp0 = 10'd627; b_exp1 = 10'd913; b_exp2 = 10'd944; b_exp3 = 10'd322;
a_sign0 = 4'd4; a_sign1 = 4'd10; a_sign2 = 4'd1; a_sign3 = 4'd3;
b_sign0 = 4'd3; b_sign1 = 4'd1; b_sign2 = 4'd16; b_sign3 = 4'd10;
@(posedge clk_i);
shared_exps0 = 8'd85;
shared_exps1 = 8'd154;
a_mant0 = 8'd217; a_mant1 = 8'd147; a_mant2 = 8'd250; a_mant3 = 8'd47;
b_mant0 = 8'd154; b_mant1 = 8'd90; b_mant2 = 8'd189; b_mant3 = 8'd28;
a_exp0 = 10'd471; a_exp1 = 10'd571; a_exp2 = 10'd942; a_exp3 = 10'd401;
b_exp0 = 10'd835; b_exp1 = 10'd856; b_exp2 = 10'd852; b_exp3 = 10'd102;
a_sign0 = 4'd8; a_sign1 = 4'd4; a_sign2 = 4'd16; a_sign3 = 4'd4;
b_sign0 = 4'd14; b_sign1 = 4'd9; b_sign2 = 4'd16; b_sign3 = 4'd3;
@(posedge clk_i);
a_mant0 = 8'd249; a_mant1 = 8'd118; a_mant2 = 8'd29; a_mant3 = 8'd236;
b_mant0 = 8'd142; b_mant1 = 8'd152; b_mant2 = 8'd4; b_mant3 = 8'd159;
a_exp0 = 10'd329; a_exp1 = 10'd560; a_exp2 = 10'd83; a_exp3 = 10'd607;
b_exp0 = 10'd141; b_exp1 = 10'd385; b_exp2 = 10'd756; b_exp3 = 10'd726;
a_sign0 = 4'd16; a_sign1 = 4'd12; a_sign2 = 4'd10; a_sign3 = 4'd1;
b_sign0 = 4'd14; b_sign1 = 4'd13; b_sign2 = 4'd3; b_sign3 = 4'd16;
@(posedge clk_i);
a_mant0 = 8'd253; a_mant1 = 8'd144; a_mant2 = 8'd241; a_mant3 = 8'd88;
b_mant0 = 8'd170; b_mant1 = 8'd1; b_mant2 = 8'd210; b_mant3 = 8'd111;
a_exp0 = 10'd794; a_exp1 = 10'd673; a_exp2 = 10'd230; a_exp3 = 10'd143;
b_exp0 = 10'd156; b_exp1 = 10'd40; b_exp2 = 10'd95; b_exp3 = 10'd438;
a_sign0 = 4'd6; a_sign1 = 4'd16; a_sign2 = 4'd2; a_sign3 = 4'd6;
b_sign0 = 4'd11; b_sign1 = 4'd11; b_sign2 = 4'd10; b_sign3 = 4'd2;
@(posedge clk_i);
a_mant0 = 8'd116; a_mant1 = 8'd229; a_mant2 = 8'd41; a_mant3 = 8'd153;
b_mant0 = 8'd240; b_mant1 = 8'd249; b_mant2 = 8'd230; b_mant3 = 8'd81;
a_exp0 = 10'd379; a_exp1 = 10'd359; a_exp2 = 10'd518; a_exp3 = 10'd178;
b_exp0 = 10'd913; b_exp1 = 10'd928; b_exp2 = 10'd360; b_exp3 = 10'd405;
a_sign0 = 4'd9; a_sign1 = 4'd11; a_sign2 = 4'd2; a_sign3 = 4'd1;
b_sign0 = 4'd8; b_sign1 = 4'd15; b_sign2 = 4'd12; b_sign3 = 4'd0;
@(posedge clk_i);
a_mant0 = 8'd0; a_mant1 = 8'd100; a_mant2 = 8'd52; a_mant3 = 8'd23;
b_mant0 = 8'd45; b_mant1 = 8'd131; b_mant2 = 8'd40; b_mant3 = 8'd248;
a_exp0 = 10'd865; a_exp1 = 10'd165; a_exp2 = 10'd217; a_exp3 = 10'd554;
b_exp0 = 10'd188; b_exp1 = 10'd132; b_exp2 = 10'd339; b_exp3 = 10'd18;
a_sign0 = 4'd9; a_sign1 = 4'd16; a_sign2 = 4'd9; a_sign3 = 4'd16;
b_sign0 = 4'd11; b_sign1 = 4'd11; b_sign2 = 4'd5; b_sign3 = 4'd14;
@(posedge clk_i);
a_mant0 = 8'd244; a_mant1 = 8'd78; a_mant2 = 8'd219; a_mant3 = 8'd4;
b_mant0 = 8'd7; b_mant1 = 8'd238; b_mant2 = 8'd79; b_mant3 = 8'd250;
a_exp0 = 10'd335; a_exp1 = 10'd439; a_exp2 = 10'd997; a_exp3 = 10'd142;
b_exp0 = 10'd789; b_exp1 = 10'd703; b_exp2 = 10'd356; b_exp3 = 10'd556;
a_sign0 = 4'd1; a_sign1 = 4'd12; a_sign2 = 4'd6; a_sign3 = 4'd6;
b_sign0 = 4'd7; b_sign1 = 4'd8; b_sign2 = 4'd9; b_sign3 = 4'd14;
@(posedge clk_i);
a_mant0 = 8'd157; a_mant1 = 8'd201; a_mant2 = 8'd155; a_mant3 = 8'd64;
b_mant0 = 8'd181; b_mant1 = 8'd236; b_mant2 = 8'd184; b_mant3 = 8'd223;
a_exp0 = 10'd612; a_exp1 = 10'd132; a_exp2 = 10'd94; a_exp3 = 10'd375;
b_exp0 = 10'd487; b_exp1 = 10'd287; b_exp2 = 10'd667; b_exp3 = 10'd1004;
a_sign0 = 4'd13; a_sign1 = 4'd0; a_sign2 = 4'd4; a_sign3 = 4'd10;
b_sign0 = 4'd4; b_sign1 = 4'd12; b_sign2 = 4'd14; b_sign3 = 4'd8;
@(posedge clk_i);
a_mant0 = 8'd51; a_mant1 = 8'd240; a_mant2 = 8'd64; a_mant3 = 8'd161;
b_mant0 = 8'd63; b_mant1 = 8'd132; b_mant2 = 8'd139; b_mant3 = 8'd29;
a_exp0 = 10'd676; a_exp1 = 10'd97; a_exp2 = 10'd661; a_exp3 = 10'd445;
b_exp0 = 10'd308; b_exp1 = 10'd838; b_exp2 = 10'd447; b_exp3 = 10'd203;
a_sign0 = 4'd16; a_sign1 = 4'd3; a_sign2 = 4'd1; a_sign3 = 4'd15;
b_sign0 = 4'd9; b_sign1 = 4'd15; b_sign2 = 4'd11; b_sign3 = 4'd4;
@(posedge clk_i);
shared_exps0 = 8'd115;
shared_exps1 = 8'd140;
a_mant0 = 8'd158; a_mant1 = 8'd202; a_mant2 = 8'd36; a_mant3 = 8'd90;
b_mant0 = 8'd85; b_mant1 = 8'd195; b_mant2 = 8'd170; b_mant3 = 8'd1;
a_exp0 = 10'd890; a_exp1 = 10'd24; a_exp2 = 10'd842; a_exp3 = 10'd890;
b_exp0 = 10'd515; b_exp1 = 10'd118; b_exp2 = 10'd449; b_exp3 = 10'd523;
a_sign0 = 4'd8; a_sign1 = 4'd10; a_sign2 = 4'd9; a_sign3 = 4'd10;
b_sign0 = 4'd2; b_sign1 = 4'd13; b_sign2 = 4'd3; b_sign3 = 4'd14;
@(posedge clk_i);
a_mant0 = 8'd194; a_mant1 = 8'd183; a_mant2 = 8'd54; a_mant3 = 8'd53;
b_mant0 = 8'd153; b_mant1 = 8'd65; b_mant2 = 8'd107; b_mant3 = 8'd6;
a_exp0 = 10'd281; a_exp1 = 10'd691; a_exp2 = 10'd259; a_exp3 = 10'd488;
b_exp0 = 10'd915; b_exp1 = 10'd260; b_exp2 = 10'd420; b_exp3 = 10'd229;
a_sign0 = 4'd13; a_sign1 = 4'd0; a_sign2 = 4'd14; a_sign3 = 4'd12;
b_sign0 = 4'd15; b_sign1 = 4'd6; b_sign2 = 4'd4; b_sign3 = 4'd15;
@(posedge clk_i);
a_mant0 = 8'd74; a_mant1 = 8'd168; a_mant2 = 8'd29; a_mant3 = 8'd104;
b_mant0 = 8'd65; b_mant1 = 8'd71; b_mant2 = 8'd1; b_mant3 = 8'd36;
a_exp0 = 10'd845; a_exp1 = 10'd234; a_exp2 = 10'd505; a_exp3 = 10'd716;
b_exp0 = 10'd165; b_exp1 = 10'd578; b_exp2 = 10'd4; b_exp3 = 10'd261;
a_sign0 = 4'd16; a_sign1 = 4'd7; a_sign2 = 4'd12; a_sign3 = 4'd3;
b_sign0 = 4'd9; b_sign1 = 4'd15; b_sign2 = 4'd5; b_sign3 = 4'd9;
@(posedge clk_i);
a_mant0 = 8'd161; a_mant1 = 8'd105; a_mant2 = 8'd241; a_mant3 = 8'd228;
b_mant0 = 8'd143; b_mant1 = 8'd224; b_mant2 = 8'd34; b_mant3 = 8'd148;
a_exp0 = 10'd898; a_exp1 = 10'd37; a_exp2 = 10'd438; a_exp3 = 10'd951;
b_exp0 = 10'd754; b_exp1 = 10'd445; b_exp2 = 10'd618; b_exp3 = 10'd326;
a_sign0 = 4'd4; a_sign1 = 4'd13; a_sign2 = 4'd2; a_sign3 = 4'd11;
b_sign0 = 4'd13; b_sign1 = 4'd14; b_sign2 = 4'd3; b_sign3 = 4'd14;
@(posedge clk_i);
a_mant0 = 8'd210; a_mant1 = 8'd255; a_mant2 = 8'd193; a_mant3 = 8'd50;
b_mant0 = 8'd241; b_mant1 = 8'd142; b_mant2 = 8'd175; b_mant3 = 8'd189;
a_exp0 = 10'd48; a_exp1 = 10'd480; a_exp2 = 10'd317; a_exp3 = 10'd596;
b_exp0 = 10'd688; b_exp1 = 10'd331; b_exp2 = 10'd34; b_exp3 = 10'd784;
a_sign0 = 4'd13; a_sign1 = 4'd0; a_sign2 = 4'd12; a_sign3 = 4'd14;
b_sign0 = 4'd6; b_sign1 = 4'd11; b_sign2 = 4'd11; b_sign3 = 4'd0;
@(posedge clk_i);
a_mant0 = 8'd5; a_mant1 = 8'd177; a_mant2 = 8'd103; a_mant3 = 8'd230;
b_mant0 = 8'd187; b_mant1 = 8'd218; b_mant2 = 8'd184; b_mant3 = 8'd86;
a_exp0 = 10'd933; a_exp1 = 10'd266; a_exp2 = 10'd779; a_exp3 = 10'd939;
b_exp0 = 10'd372; b_exp1 = 10'd916; b_exp2 = 10'd590; b_exp3 = 10'd880;
a_sign0 = 4'd3; a_sign1 = 4'd9; a_sign2 = 4'd15; a_sign3 = 4'd1;
b_sign0 = 4'd13; b_sign1 = 4'd10; b_sign2 = 4'd12; b_sign3 = 4'd6;
@(posedge clk_i);
a_mant0 = 8'd156; a_mant1 = 8'd231; a_mant2 = 8'd121; a_mant3 = 8'd27;
b_mant0 = 8'd90; b_mant1 = 8'd177; b_mant2 = 8'd118; b_mant3 = 8'd61;
a_exp0 = 10'd627; a_exp1 = 10'd69; a_exp2 = 10'd887; a_exp3 = 10'd397;
b_exp0 = 10'd457; b_exp1 = 10'd701; b_exp2 = 10'd412; b_exp3 = 10'd477;
a_sign0 = 4'd10; a_sign1 = 4'd3; a_sign2 = 4'd9; a_sign3 = 4'd0;
b_sign0 = 4'd5; b_sign1 = 4'd3; b_sign2 = 4'd4; b_sign3 = 4'd12;
@(posedge clk_i);
a_mant0 = 8'd108; a_mant1 = 8'd188; a_mant2 = 8'd148; a_mant3 = 8'd34;
b_mant0 = 8'd59; b_mant1 = 8'd207; b_mant2 = 8'd216; b_mant3 = 8'd109;
a_exp0 = 10'd888; a_exp1 = 10'd732; a_exp2 = 10'd943; a_exp3 = 10'd15;
b_exp0 = 10'd473; b_exp1 = 10'd872; b_exp2 = 10'd532; b_exp3 = 10'd203;
a_sign0 = 4'd3; a_sign1 = 4'd0; a_sign2 = 4'd10; a_sign3 = 4'd0;
b_sign0 = 4'd0; b_sign1 = 4'd3; b_sign2 = 4'd4; b_sign3 = 4'd8;
@(posedge clk_i);
shared_exps0 = 8'd117;
shared_exps1 = 8'd147;
rstn = 0;
@(posedge clk_i);
rstn = 1;
a_mant0 = 8'd34; a_mant1 = 8'd17; a_mant2 = 8'd18; a_mant3 = 8'd88;
b_mant0 = 8'd208; b_mant1 = 8'd249; b_mant2 = 8'd56; b_mant3 = 8'd136;
a_exp0 = 10'd651; a_exp1 = 10'd848; a_exp2 = 10'd7; a_exp3 = 10'd512;
b_exp0 = 10'd1003; b_exp1 = 10'd81; b_exp2 = 10'd509; b_exp3 = 10'd726;
a_sign0 = 4'd5; a_sign1 = 4'd9; a_sign2 = 4'd12; a_sign3 = 4'd15;
b_sign0 = 4'd16; b_sign1 = 4'd14; b_sign2 = 4'd8; b_sign3 = 4'd14;
@(posedge clk_i);
a_mant0 = 8'd209; a_mant1 = 8'd194; a_mant2 = 8'd226; a_mant3 = 8'd79;
b_mant0 = 8'd14; b_mant1 = 8'd219; b_mant2 = 8'd189; b_mant3 = 8'd134;
a_exp0 = 10'd485; a_exp1 = 10'd826; a_exp2 = 10'd995; a_exp3 = 10'd898;
b_exp0 = 10'd373; b_exp1 = 10'd223; b_exp2 = 10'd43; b_exp3 = 10'd349;
a_sign0 = 4'd14; a_sign1 = 4'd14; a_sign2 = 4'd10; a_sign3 = 4'd15;
b_sign0 = 4'd14; b_sign1 = 4'd8; b_sign2 = 4'd11; b_sign3 = 4'd16;
@(posedge clk_i);
a_mant0 = 8'd49; a_mant1 = 8'd3; a_mant2 = 8'd197; a_mant3 = 8'd32;
b_mant0 = 8'd22; b_mant1 = 8'd163; b_mant2 = 8'd121; b_mant3 = 8'd16;
a_exp0 = 10'd22; a_exp1 = 10'd199; a_exp2 = 10'd310; a_exp3 = 10'd992;
b_exp0 = 10'd934; b_exp1 = 10'd502; b_exp2 = 10'd387; b_exp3 = 10'd516;
a_sign0 = 4'd11; a_sign1 = 4'd7; a_sign2 = 4'd15; a_sign3 = 4'd14;
b_sign0 = 4'd7; b_sign1 = 4'd0; b_sign2 = 4'd2; b_sign3 = 4'd14;
@(posedge clk_i);
a_mant0 = 8'd205; a_mant1 = 8'd136; a_mant2 = 8'd188; a_mant3 = 8'd110;
b_mant0 = 8'd187; b_mant1 = 8'd182; b_mant2 = 8'd141; b_mant3 = 8'd194;
a_exp0 = 10'd943; a_exp1 = 10'd500; a_exp2 = 10'd808; a_exp3 = 10'd691;
b_exp0 = 10'd763; b_exp1 = 10'd386; b_exp2 = 10'd808; b_exp3 = 10'd53;
a_sign0 = 4'd4; a_sign1 = 4'd9; a_sign2 = 4'd0; a_sign3 = 4'd11;
b_sign0 = 4'd9; b_sign1 = 4'd9; b_sign2 = 4'd3; b_sign3 = 4'd7;
@(posedge clk_i);
a_mant0 = 8'd29; a_mant1 = 8'd112; a_mant2 = 8'd188; a_mant3 = 8'd86;
b_mant0 = 8'd20; b_mant1 = 8'd244; b_mant2 = 8'd188; b_mant3 = 8'd164;
a_exp0 = 10'd287; a_exp1 = 10'd350; a_exp2 = 10'd759; a_exp3 = 10'd327;
b_exp0 = 10'd200; b_exp1 = 10'd673; b_exp2 = 10'd300; b_exp3 = 10'd520;
a_sign0 = 4'd8; a_sign1 = 4'd6; a_sign2 = 4'd16; a_sign3 = 4'd10;
b_sign0 = 4'd15; b_sign1 = 4'd13; b_sign2 = 4'd3; b_sign3 = 4'd7;
@(posedge clk_i);
a_mant0 = 8'd152; a_mant1 = 8'd104; a_mant2 = 8'd42; a_mant3 = 8'd72;
b_mant0 = 8'd154; b_mant1 = 8'd82; b_mant2 = 8'd192; b_mant3 = 8'd116;
a_exp0 = 10'd754; a_exp1 = 10'd417; a_exp2 = 10'd88; a_exp3 = 10'd461;
b_exp0 = 10'd997; b_exp1 = 10'd966; b_exp2 = 10'd845; b_exp3 = 10'd507;
a_sign0 = 4'd3; a_sign1 = 4'd4; a_sign2 = 4'd16; a_sign3 = 4'd14;
b_sign0 = 4'd4; b_sign1 = 4'd8; b_sign2 = 4'd9; b_sign3 = 4'd11;
@(posedge clk_i);
a_mant0 = 8'd223; a_mant1 = 8'd5; a_mant2 = 8'd30; a_mant3 = 8'd231;
b_mant0 = 8'd43; b_mant1 = 8'd27; b_mant2 = 8'd66; b_mant3 = 8'd51;
a_exp0 = 10'd403; a_exp1 = 10'd135; a_exp2 = 10'd120; a_exp3 = 10'd573;
b_exp0 = 10'd641; b_exp1 = 10'd548; b_exp2 = 10'd348; b_exp3 = 10'd181;
a_sign0 = 4'd12; a_sign1 = 4'd13; a_sign2 = 4'd9; a_sign3 = 4'd4;
b_sign0 = 4'd7; b_sign1 = 4'd8; b_sign2 = 4'd13; b_sign3 = 4'd6;
@(posedge clk_i);
shared_exps0 = 8'd139;
shared_exps1 = 8'd127;
a_mant0 = 8'd194; a_mant1 = 8'd249; a_mant2 = 8'd112; a_mant3 = 8'd26;
b_mant0 = 8'd198; b_mant1 = 8'd8; b_mant2 = 8'd137; b_mant3 = 8'd193;
a_exp0 = 10'd191; a_exp1 = 10'd704; a_exp2 = 10'd426; a_exp3 = 10'd692;
b_exp0 = 10'd859; b_exp1 = 10'd53; b_exp2 = 10'd485; b_exp3 = 10'd250;
a_sign0 = 4'd14; a_sign1 = 4'd2; a_sign2 = 4'd16; a_sign3 = 4'd12;
b_sign0 = 4'd5; b_sign1 = 4'd10; b_sign2 = 4'd13; b_sign3 = 4'd14;
@(posedge clk_i);
a_mant0 = 8'd248; a_mant1 = 8'd128; a_mant2 = 8'd236; a_mant3 = 8'd6;
b_mant0 = 8'd212; b_mant1 = 8'd132; b_mant2 = 8'd95; b_mant3 = 8'd7;
a_exp0 = 10'd873; a_exp1 = 10'd449; a_exp2 = 10'd682; a_exp3 = 10'd923;
b_exp0 = 10'd739; b_exp1 = 10'd973; b_exp2 = 10'd924; b_exp3 = 10'd683;
a_sign0 = 4'd14; a_sign1 = 4'd9; a_sign2 = 4'd16; a_sign3 = 4'd10;
b_sign0 = 4'd2; b_sign1 = 4'd2; b_sign2 = 4'd6; b_sign3 = 4'd9;
@(posedge clk_i);
a_mant0 = 8'd166; a_mant1 = 8'd248; a_mant2 = 8'd78; a_mant3 = 8'd1;
b_mant0 = 8'd228; b_mant1 = 8'd253; b_mant2 = 8'd97; b_mant3 = 8'd17;
a_exp0 = 10'd154; a_exp1 = 10'd225; a_exp2 = 10'd353; a_exp3 = 10'd41;
b_exp0 = 10'd47; b_exp1 = 10'd740; b_exp2 = 10'd236; b_exp3 = 10'd821;
a_sign0 = 4'd12; a_sign1 = 4'd3; a_sign2 = 4'd2; a_sign3 = 4'd11;
b_sign0 = 4'd2; b_sign1 = 4'd12; b_sign2 = 4'd11; b_sign3 = 4'd5;
@(posedge clk_i);
a_mant0 = 8'd204; a_mant1 = 8'd53; a_mant2 = 8'd4; a_mant3 = 8'd100;
b_mant0 = 8'd216; b_mant1 = 8'd63; b_mant2 = 8'd5; b_mant3 = 8'd90;
a_exp0 = 10'd583; a_exp1 = 10'd278; a_exp2 = 10'd923; a_exp3 = 10'd296;
b_exp0 = 10'd869; b_exp1 = 10'd211; b_exp2 = 10'd89; b_exp3 = 10'd30;
a_sign0 = 4'd10; a_sign1 = 4'd8; a_sign2 = 4'd11; a_sign3 = 4'd9;
b_sign0 = 4'd14; b_sign1 = 4'd5; b_sign2 = 4'd2; b_sign3 = 4'd5;
@(posedge clk_i);
a_mant0 = 8'd219; a_mant1 = 8'd134; a_mant2 = 8'd73; a_mant3 = 8'd199;
b_mant0 = 8'd237; b_mant1 = 8'd116; b_mant2 = 8'd130; b_mant3 = 8'd233;
a_exp0 = 10'd799; a_exp1 = 10'd505; a_exp2 = 10'd112; a_exp3 = 10'd155;
b_exp0 = 10'd293; b_exp1 = 10'd122; b_exp2 = 10'd709; b_exp3 = 10'd18;
a_sign0 = 4'd3; a_sign1 = 4'd4; a_sign2 = 4'd0; a_sign3 = 4'd5;
b_sign0 = 4'd1; b_sign1 = 4'd16; b_sign2 = 4'd0; b_sign3 = 4'd3;
@(posedge clk_i);
a_mant0 = 8'd251; a_mant1 = 8'd162; a_mant2 = 8'd81; a_mant3 = 8'd112;
b_mant0 = 8'd30; b_mant1 = 8'd36; b_mant2 = 8'd252; b_mant3 = 8'd38;
a_exp0 = 10'd232; a_exp1 = 10'd245; a_exp2 = 10'd176; a_exp3 = 10'd103;
b_exp0 = 10'd467; b_exp1 = 10'd835; b_exp2 = 10'd208; b_exp3 = 10'd674;
a_sign0 = 4'd13; a_sign1 = 4'd6; a_sign2 = 4'd10; a_sign3 = 4'd12;
b_sign0 = 4'd8; b_sign1 = 4'd6; b_sign2 = 4'd13; b_sign3 = 4'd2;
@(posedge clk_i);
a_mant0 = 8'd11; a_mant1 = 8'd35; a_mant2 = 8'd175; a_mant3 = 8'd138;
b_mant0 = 8'd38; b_mant1 = 8'd58; b_mant2 = 8'd56; b_mant3 = 8'd234;
a_exp0 = 10'd993; a_exp1 = 10'd392; a_exp2 = 10'd56; a_exp3 = 10'd560;
b_exp0 = 10'd165; b_exp1 = 10'd276; b_exp2 = 10'd382; b_exp3 = 10'd111;
a_sign0 = 4'd11; a_sign1 = 4'd7; a_sign2 = 4'd15; a_sign3 = 4'd6;
b_sign0 = 4'd13; b_sign1 = 4'd8; b_sign2 = 4'd3; b_sign3 = 4'd2;
@(posedge clk_i);
a_mant0 = 8'd131; a_mant1 = 8'd64; a_mant2 = 8'd196; a_mant3 = 8'd227;
b_mant0 = 8'd101; b_mant1 = 8'd181; b_mant2 = 8'd208; b_mant3 = 8'd66;
a_exp0 = 10'd403; a_exp1 = 10'd515; a_exp2 = 10'd772; a_exp3 = 10'd650;
b_exp0 = 10'd35; b_exp1 = 10'd6; b_exp2 = 10'd284; b_exp3 = 10'd995;
a_sign0 = 4'd15; a_sign1 = 4'd0; a_sign2 = 4'd6; a_sign3 = 4'd3;
b_sign0 = 4'd14; b_sign1 = 4'd14; b_sign2 = 4'd0; b_sign3 = 4'd14;
@(posedge clk_i);
shared_exps0 = 8'd129;
shared_exps1 = 8'd113;
a_mant0 = 8'd160; a_mant1 = 8'd119; a_mant2 = 8'd66; a_mant3 = 8'd215;
b_mant0 = 8'd197; b_mant1 = 8'd156; b_mant2 = 8'd148; b_mant3 = 8'd167;
a_exp0 = 10'd414; a_exp1 = 10'd751; a_exp2 = 10'd815; a_exp3 = 10'd972;
b_exp0 = 10'd604; b_exp1 = 10'd429; b_exp2 = 10'd926; b_exp3 = 10'd290;
a_sign0 = 4'd13; a_sign1 = 4'd10; a_sign2 = 4'd4; a_sign3 = 4'd9;
b_sign0 = 4'd11; b_sign1 = 4'd5; b_sign2 = 4'd3; b_sign3 = 4'd11;
@(posedge clk_i);
a_mant0 = 8'd176; a_mant1 = 8'd69; a_mant2 = 8'd96; a_mant3 = 8'd217;
b_mant0 = 8'd235; b_mant1 = 8'd27; b_mant2 = 8'd62; b_mant3 = 8'd55;
a_exp0 = 10'd834; a_exp1 = 10'd714; a_exp2 = 10'd478; a_exp3 = 10'd162;
b_exp0 = 10'd503; b_exp1 = 10'd806; b_exp2 = 10'd916; b_exp3 = 10'd146;
a_sign0 = 4'd0; a_sign1 = 4'd3; a_sign2 = 4'd16; a_sign3 = 4'd16;
b_sign0 = 4'd6; b_sign1 = 4'd15; b_sign2 = 4'd3; b_sign3 = 4'd2;
@(posedge clk_i);
a_mant0 = 8'd43; a_mant1 = 8'd155; a_mant2 = 8'd187; a_mant3 = 8'd59;
b_mant0 = 8'd13; b_mant1 = 8'd192; b_mant2 = 8'd152; b_mant3 = 8'd145;
a_exp0 = 10'd744; a_exp1 = 10'd336; a_exp2 = 10'd956; a_exp3 = 10'd114;
b_exp0 = 10'd577; b_exp1 = 10'd583; b_exp2 = 10'd356; b_exp3 = 10'd557;
a_sign0 = 4'd15; a_sign1 = 4'd12; a_sign2 = 4'd15; a_sign3 = 4'd16;
b_sign0 = 4'd3; b_sign1 = 4'd5; b_sign2 = 4'd11; b_sign3 = 4'd12;
@(posedge clk_i);
a_mant0 = 8'd129; a_mant1 = 8'd248; a_mant2 = 8'd171; a_mant3 = 8'd78;
b_mant0 = 8'd25; b_mant1 = 8'd176; b_mant2 = 8'd31; b_mant3 = 8'd246;
a_exp0 = 10'd495; a_exp1 = 10'd884; a_exp2 = 10'd735; a_exp3 = 10'd698;
b_exp0 = 10'd17; b_exp1 = 10'd69; b_exp2 = 10'd440; b_exp3 = 10'd121;
a_sign0 = 4'd14; a_sign1 = 4'd6; a_sign2 = 4'd16; a_sign3 = 4'd12;
b_sign0 = 4'd16; b_sign1 = 4'd3; b_sign2 = 4'd13; b_sign3 = 4'd1;
@(posedge clk_i);
a_mant0 = 8'd222; a_mant1 = 8'd171; a_mant2 = 8'd246; a_mant3 = 8'd15;
b_mant0 = 8'd230; b_mant1 = 8'd140; b_mant2 = 8'd7; b_mant3 = 8'd254;
a_exp0 = 10'd891; a_exp1 = 10'd932; a_exp2 = 10'd257; a_exp3 = 10'd121;
b_exp0 = 10'd140; b_exp1 = 10'd562; b_exp2 = 10'd243; b_exp3 = 10'd809;
a_sign0 = 4'd7; a_sign1 = 4'd1; a_sign2 = 4'd3; a_sign3 = 4'd8;
b_sign0 = 4'd6; b_sign1 = 4'd16; b_sign2 = 4'd11; b_sign3 = 4'd9;
@(posedge clk_i);
a_mant0 = 8'd162; a_mant1 = 8'd115; a_mant2 = 8'd222; a_mant3 = 8'd42;
b_mant0 = 8'd13; b_mant1 = 8'd187; b_mant2 = 8'd16; b_mant3 = 8'd222;
a_exp0 = 10'd867; a_exp1 = 10'd437; a_exp2 = 10'd153; a_exp3 = 10'd674;
b_exp0 = 10'd551; b_exp1 = 10'd917; b_exp2 = 10'd276; b_exp3 = 10'd289;
a_sign0 = 4'd14; a_sign1 = 4'd16; a_sign2 = 4'd14; a_sign3 = 4'd9;
b_sign0 = 4'd8; b_sign1 = 4'd10; b_sign2 = 4'd15; b_sign3 = 4'd15;
@(posedge clk_i);
a_mant0 = 8'd152; a_mant1 = 8'd241; a_mant2 = 8'd35; a_mant3 = 8'd27;
b_mant0 = 8'd200; b_mant1 = 8'd235; b_mant2 = 8'd157; b_mant3 = 8'd157;
a_exp0 = 10'd249; a_exp1 = 10'd935; a_exp2 = 10'd666; a_exp3 = 10'd911;
b_exp0 = 10'd161; b_exp1 = 10'd233; b_exp2 = 10'd997; b_exp3 = 10'd170;
a_sign0 = 4'd7; a_sign1 = 4'd13; a_sign2 = 4'd2; a_sign3 = 4'd8;
b_sign0 = 4'd10; b_sign1 = 4'd1; b_sign2 = 4'd9; b_sign3 = 4'd6;
@(posedge clk_i);
a_mant0 = 8'd95; a_mant1 = 8'd147; a_mant2 = 8'd173; a_mant3 = 8'd28;
b_mant0 = 8'd33; b_mant1 = 8'd163; b_mant2 = 8'd69; b_mant3 = 8'd155;
a_exp0 = 10'd1005; a_exp1 = 10'd135; a_exp2 = 10'd479; a_exp3 = 10'd940;
b_exp0 = 10'd995; b_exp1 = 10'd152; b_exp2 = 10'd995; b_exp3 = 10'd1014;
a_sign0 = 4'd15; a_sign1 = 4'd0; a_sign2 = 4'd8; a_sign3 = 4'd12;
b_sign0 = 4'd5; b_sign1 = 4'd16; b_sign2 = 4'd4; b_sign3 = 4'd10;
@(posedge clk_i);
shared_exps0 = 8'd118;
shared_exps1 = 8'd137;
a_mant0 = 8'd60; a_mant1 = 8'd119; a_mant2 = 8'd36; a_mant3 = 8'd139;
b_mant0 = 8'd237; b_mant1 = 8'd181; b_mant2 = 8'd25; b_mant3 = 8'd0;
a_exp0 = 10'd973; a_exp1 = 10'd467; a_exp2 = 10'd857; a_exp3 = 10'd414;
b_exp0 = 10'd466; b_exp1 = 10'd627; b_exp2 = 10'd401; b_exp3 = 10'd19;
a_sign0 = 4'd2; a_sign1 = 4'd0; a_sign2 = 4'd15; a_sign3 = 4'd2;
b_sign0 = 4'd4; b_sign1 = 4'd7; b_sign2 = 4'd15; b_sign3 = 4'd12;
@(posedge clk_i);
a_mant0 = 8'd68; a_mant1 = 8'd229; a_mant2 = 8'd129; a_mant3 = 8'd206;
b_mant0 = 8'd99; b_mant1 = 8'd150; b_mant2 = 8'd40; b_mant3 = 8'd214;
a_exp0 = 10'd625; a_exp1 = 10'd945; a_exp2 = 10'd88; a_exp3 = 10'd846;
b_exp0 = 10'd100; b_exp1 = 10'd416; b_exp2 = 10'd770; b_exp3 = 10'd1;
a_sign0 = 4'd8; a_sign1 = 4'd10; a_sign2 = 4'd10; a_sign3 = 4'd14;
b_sign0 = 4'd11; b_sign1 = 4'd16; b_sign2 = 4'd12; b_sign3 = 4'd1;
@(posedge clk_i);
a_mant0 = 8'd8; a_mant1 = 8'd45; a_mant2 = 8'd46; a_mant3 = 8'd173;
b_mant0 = 8'd96; b_mant1 = 8'd77; b_mant2 = 8'd165; b_mant3 = 8'd172;
a_exp0 = 10'd157; a_exp1 = 10'd401; a_exp2 = 10'd6; a_exp3 = 10'd207;
b_exp0 = 10'd38; b_exp1 = 10'd487; b_exp2 = 10'd582; b_exp3 = 10'd379;
a_sign0 = 4'd10; a_sign1 = 4'd2; a_sign2 = 4'd7; a_sign3 = 4'd2;
b_sign0 = 4'd4; b_sign1 = 4'd1; b_sign2 = 4'd4; b_sign3 = 4'd3;
@(posedge clk_i);
a_mant0 = 8'd137; a_mant1 = 8'd10; a_mant2 = 8'd13; a_mant3 = 8'd171;
b_mant0 = 8'd121; b_mant1 = 8'd103; b_mant2 = 8'd107; b_mant3 = 8'd180;
a_exp0 = 10'd301; a_exp1 = 10'd846; a_exp2 = 10'd40; a_exp3 = 10'd425;
b_exp0 = 10'd54; b_exp1 = 10'd91; b_exp2 = 10'd682; b_exp3 = 10'd970;
a_sign0 = 4'd4; a_sign1 = 4'd2; a_sign2 = 4'd4; a_sign3 = 4'd3;
b_sign0 = 4'd12; b_sign1 = 4'd2; b_sign2 = 4'd7; b_sign3 = 4'd9;
@(posedge clk_i);
a_mant0 = 8'd247; a_mant1 = 8'd195; a_mant2 = 8'd19; a_mant3 = 8'd197;
b_mant0 = 8'd90; b_mant1 = 8'd139; b_mant2 = 8'd6; b_mant3 = 8'd8;
a_exp0 = 10'd517; a_exp1 = 10'd158; a_exp2 = 10'd67; a_exp3 = 10'd985;
b_exp0 = 10'd393; b_exp1 = 10'd503; b_exp2 = 10'd753; b_exp3 = 10'd711;
a_sign0 = 4'd12; a_sign1 = 4'd16; a_sign2 = 4'd6; a_sign3 = 4'd11;
b_sign0 = 4'd8; b_sign1 = 4'd2; b_sign2 = 4'd10; b_sign3 = 4'd15;
@(posedge clk_i);
a_mant0 = 8'd24; a_mant1 = 8'd217; a_mant2 = 8'd136; a_mant3 = 8'd170;
b_mant0 = 8'd84; b_mant1 = 8'd129; b_mant2 = 8'd120; b_mant3 = 8'd224;
a_exp0 = 10'd237; a_exp1 = 10'd693; a_exp2 = 10'd453; a_exp3 = 10'd660;
b_exp0 = 10'd735; b_exp1 = 10'd687; b_exp2 = 10'd764; b_exp3 = 10'd768;
a_sign0 = 4'd15; a_sign1 = 4'd8; a_sign2 = 4'd7; a_sign3 = 4'd2;
b_sign0 = 4'd10; b_sign1 = 4'd0; b_sign2 = 4'd3; b_sign3 = 4'd0;
@(posedge clk_i);
a_mant0 = 8'd239; a_mant1 = 8'd75; a_mant2 = 8'd19; a_mant3 = 8'd47;
b_mant0 = 8'd183; b_mant1 = 8'd67; b_mant2 = 8'd22; b_mant3 = 8'd186;
a_exp0 = 10'd450; a_exp1 = 10'd762; a_exp2 = 10'd199; a_exp3 = 10'd273;
b_exp0 = 10'd858; b_exp1 = 10'd790; b_exp2 = 10'd277; b_exp3 = 10'd14;
a_sign0 = 4'd1; a_sign1 = 4'd10; a_sign2 = 4'd4; a_sign3 = 4'd4;
b_sign0 = 4'd0; b_sign1 = 4'd7; b_sign2 = 4'd12; b_sign3 = 4'd14;
@(posedge clk_i);
a_mant0 = 8'd32; a_mant1 = 8'd166; a_mant2 = 8'd130; a_mant3 = 8'd23;
b_mant0 = 8'd84; b_mant1 = 8'd208; b_mant2 = 8'd53; b_mant3 = 8'd218;
a_exp0 = 10'd679; a_exp1 = 10'd386; a_exp2 = 10'd816; a_exp3 = 10'd976;
b_exp0 = 10'd121; b_exp1 = 10'd369; b_exp2 = 10'd652; b_exp3 = 10'd613;
a_sign0 = 4'd10; a_sign1 = 4'd1; a_sign2 = 4'd2; a_sign3 = 4'd9;
b_sign0 = 4'd10; b_sign1 = 4'd12; b_sign2 = 4'd6; b_sign3 = 4'd8;
@(posedge clk_i);
shared_exps0 = 8'd139;
shared_exps1 = 8'd132;
rstn = 0;
@(posedge clk_i);
rstn = 1;
a_mant0 = 8'd101; a_mant1 = 8'd21; a_mant2 = 8'd60; a_mant3 = 8'd131;
b_mant0 = 8'd185; b_mant1 = 8'd139; b_mant2 = 8'd145; b_mant3 = 8'd73;
a_exp0 = 10'd200; a_exp1 = 10'd854; a_exp2 = 10'd744; a_exp3 = 10'd726;
b_exp0 = 10'd585; b_exp1 = 10'd266; b_exp2 = 10'd916; b_exp3 = 10'd54;
a_sign0 = 4'd2; a_sign1 = 4'd10; a_sign2 = 4'd11; a_sign3 = 4'd10;
b_sign0 = 4'd3; b_sign1 = 4'd9; b_sign2 = 4'd0; b_sign3 = 4'd14;
@(posedge clk_i);
a_mant0 = 8'd240; a_mant1 = 8'd77; a_mant2 = 8'd214; a_mant3 = 8'd125;
b_mant0 = 8'd196; b_mant1 = 8'd203; b_mant2 = 8'd143; b_mant3 = 8'd128;
a_exp0 = 10'd976; a_exp1 = 10'd854; a_exp2 = 10'd634; a_exp3 = 10'd568;
b_exp0 = 10'd660; b_exp1 = 10'd773; b_exp2 = 10'd332; b_exp3 = 10'd123;
a_sign0 = 4'd13; a_sign1 = 4'd1; a_sign2 = 4'd8; a_sign3 = 4'd8;
b_sign0 = 4'd4; b_sign1 = 4'd16; b_sign2 = 4'd5; b_sign3 = 4'd5;
@(posedge clk_i);
a_mant0 = 8'd41; a_mant1 = 8'd58; a_mant2 = 8'd89; a_mant3 = 8'd76;
b_mant0 = 8'd111; b_mant1 = 8'd233; b_mant2 = 8'd163; b_mant3 = 8'd136;
a_exp0 = 10'd904; a_exp1 = 10'd698; a_exp2 = 10'd240; a_exp3 = 10'd304;
b_exp0 = 10'd309; b_exp1 = 10'd490; b_exp2 = 10'd735; b_exp3 = 10'd16;
a_sign0 = 4'd2; a_sign1 = 4'd9; a_sign2 = 4'd2; a_sign3 = 4'd11;
b_sign0 = 4'd8; b_sign1 = 4'd14; b_sign2 = 4'd7; b_sign3 = 4'd1;
@(posedge clk_i);
a_mant0 = 8'd19; a_mant1 = 8'd32; a_mant2 = 8'd166; a_mant3 = 8'd185;
b_mant0 = 8'd34; b_mant1 = 8'd228; b_mant2 = 8'd149; b_mant3 = 8'd56;
a_exp0 = 10'd887; a_exp1 = 10'd432; a_exp2 = 10'd127; a_exp3 = 10'd413;
b_exp0 = 10'd336; b_exp1 = 10'd443; b_exp2 = 10'd261; b_exp3 = 10'd451;
a_sign0 = 4'd10; a_sign1 = 4'd5; a_sign2 = 4'd6; a_sign3 = 4'd16;
b_sign0 = 4'd6; b_sign1 = 4'd8; b_sign2 = 4'd12; b_sign3 = 4'd5;
@(posedge clk_i);
a_mant0 = 8'd241; a_mant1 = 8'd114; a_mant2 = 8'd217; a_mant3 = 8'd164;
b_mant0 = 8'd118; b_mant1 = 8'd174; b_mant2 = 8'd44; b_mant3 = 8'd145;
a_exp0 = 10'd389; a_exp1 = 10'd786; a_exp2 = 10'd45; a_exp3 = 10'd649;
b_exp0 = 10'd883; b_exp1 = 10'd667; b_exp2 = 10'd1001; b_exp3 = 10'd848;
a_sign0 = 4'd12; a_sign1 = 4'd14; a_sign2 = 4'd11; a_sign3 = 4'd9;
b_sign0 = 4'd13; b_sign1 = 4'd12; b_sign2 = 4'd14; b_sign3 = 4'd12;
@(posedge clk_i);
a_mant0 = 8'd222; a_mant1 = 8'd95; a_mant2 = 8'd166; a_mant3 = 8'd179;
b_mant0 = 8'd95; b_mant1 = 8'd82; b_mant2 = 8'd15; b_mant3 = 8'd239;
a_exp0 = 10'd248; a_exp1 = 10'd906; a_exp2 = 10'd461; a_exp3 = 10'd727;
b_exp0 = 10'd876; b_exp1 = 10'd740; b_exp2 = 10'd191; b_exp3 = 10'd561;
a_sign0 = 4'd16; a_sign1 = 4'd10; a_sign2 = 4'd11; a_sign3 = 4'd11;
b_sign0 = 4'd7; b_sign1 = 4'd9; b_sign2 = 4'd15; b_sign3 = 4'd4;
@(posedge clk_i);
a_mant0 = 8'd154; a_mant1 = 8'd241; a_mant2 = 8'd3; a_mant3 = 8'd6;
b_mant0 = 8'd236; b_mant1 = 8'd188; b_mant2 = 8'd202; b_mant3 = 8'd108;
a_exp0 = 10'd206; a_exp1 = 10'd630; a_exp2 = 10'd714; a_exp3 = 10'd380;
b_exp0 = 10'd721; b_exp1 = 10'd763; b_exp2 = 10'd439; b_exp3 = 10'd336;
a_sign0 = 4'd7; a_sign1 = 4'd1; a_sign2 = 4'd10; a_sign3 = 4'd4;
b_sign0 = 4'd0; b_sign1 = 4'd16; b_sign2 = 4'd7; b_sign3 = 4'd6;
@(posedge clk_i);
shared_exps0 = 8'd110;
shared_exps1 = 8'd131;
a_mant0 = 8'd115; a_mant1 = 8'd196; a_mant2 = 8'd88; a_mant3 = 8'd213;
b_mant0 = 8'd233; b_mant1 = 8'd3; b_mant2 = 8'd147; b_mant3 = 8'd170;
a_exp0 = 10'd425; a_exp1 = 10'd380; a_exp2 = 10'd1013; a_exp3 = 10'd1018;
b_exp0 = 10'd753; b_exp1 = 10'd343; b_exp2 = 10'd955; b_exp3 = 10'd627;
a_sign0 = 4'd15; a_sign1 = 4'd8; a_sign2 = 4'd10; a_sign3 = 4'd3;
b_sign0 = 4'd11; b_sign1 = 4'd10; b_sign2 = 4'd13; b_sign3 = 4'd16;
@(posedge clk_i);
a_mant0 = 8'd82; a_mant1 = 8'd23; a_mant2 = 8'd155; a_mant3 = 8'd7;
b_mant0 = 8'd153; b_mant1 = 8'd157; b_mant2 = 8'd20; b_mant3 = 8'd176;
a_exp0 = 10'd972; a_exp1 = 10'd398; a_exp2 = 10'd623; a_exp3 = 10'd59;
b_exp0 = 10'd578; b_exp1 = 10'd64; b_exp2 = 10'd287; b_exp3 = 10'd476;
a_sign0 = 4'd15; a_sign1 = 4'd9; a_sign2 = 4'd6; a_sign3 = 4'd2;
b_sign0 = 4'd4; b_sign1 = 4'd6; b_sign2 = 4'd6; b_sign3 = 4'd11;
@(posedge clk_i);
a_mant0 = 8'd49; a_mant1 = 8'd139; a_mant2 = 8'd103; a_mant3 = 8'd223;
b_mant0 = 8'd13; b_mant1 = 8'd35; b_mant2 = 8'd232; b_mant3 = 8'd191;
a_exp0 = 10'd901; a_exp1 = 10'd699; a_exp2 = 10'd491; a_exp3 = 10'd471;
b_exp0 = 10'd1013; b_exp1 = 10'd796; b_exp2 = 10'd1007; b_exp3 = 10'd373;
a_sign0 = 4'd8; a_sign1 = 4'd3; a_sign2 = 4'd10; a_sign3 = 4'd12;
b_sign0 = 4'd14; b_sign1 = 4'd6; b_sign2 = 4'd11; b_sign3 = 4'd8;
@(posedge clk_i);
a_mant0 = 8'd92; a_mant1 = 8'd91; a_mant2 = 8'd107; a_mant3 = 8'd73;
b_mant0 = 8'd242; b_mant1 = 8'd202; b_mant2 = 8'd186; b_mant3 = 8'd190;
a_exp0 = 10'd974; a_exp1 = 10'd197; a_exp2 = 10'd572; a_exp3 = 10'd20;
b_exp0 = 10'd58; b_exp1 = 10'd639; b_exp2 = 10'd237; b_exp3 = 10'd115;
a_sign0 = 4'd12; a_sign1 = 4'd0; a_sign2 = 4'd3; a_sign3 = 4'd15;
b_sign0 = 4'd5; b_sign1 = 4'd12; b_sign2 = 4'd8; b_sign3 = 4'd9;
@(posedge clk_i);
a_mant0 = 8'd196; a_mant1 = 8'd197; a_mant2 = 8'd11; a_mant3 = 8'd50;
b_mant0 = 8'd254; b_mant1 = 8'd221; b_mant2 = 8'd116; b_mant3 = 8'd211;
a_exp0 = 10'd334; a_exp1 = 10'd603; a_exp2 = 10'd710; a_exp3 = 10'd568;
b_exp0 = 10'd795; b_exp1 = 10'd60; b_exp2 = 10'd362; b_exp3 = 10'd678;
a_sign0 = 4'd12; a_sign1 = 4'd9; a_sign2 = 4'd5; a_sign3 = 4'd11;
b_sign0 = 4'd7; b_sign1 = 4'd2; b_sign2 = 4'd14; b_sign3 = 4'd9;
@(posedge clk_i);
a_mant0 = 8'd105; a_mant1 = 8'd11; a_mant2 = 8'd190; a_mant3 = 8'd189;
b_mant0 = 8'd58; b_mant1 = 8'd19; b_mant2 = 8'd122; b_mant3 = 8'd106;
a_exp0 = 10'd100; a_exp1 = 10'd150; a_exp2 = 10'd182; a_exp3 = 10'd283;
b_exp0 = 10'd925; b_exp1 = 10'd79; b_exp2 = 10'd69; b_exp3 = 10'd454;
a_sign0 = 4'd16; a_sign1 = 4'd5; a_sign2 = 4'd6; a_sign3 = 4'd8;
b_sign0 = 4'd2; b_sign1 = 4'd11; b_sign2 = 4'd16; b_sign3 = 4'd15;
@(posedge clk_i);
a_mant0 = 8'd75; a_mant1 = 8'd135; a_mant2 = 8'd2; a_mant3 = 8'd162;
b_mant0 = 8'd44; b_mant1 = 8'd222; b_mant2 = 8'd179; b_mant3 = 8'd33;
a_exp0 = 10'd679; a_exp1 = 10'd467; a_exp2 = 10'd813; a_exp3 = 10'd917;
b_exp0 = 10'd719; b_exp1 = 10'd856; b_exp2 = 10'd812; b_exp3 = 10'd327;
a_sign0 = 4'd2; a_sign1 = 4'd16; a_sign2 = 4'd7; a_sign3 = 4'd1;
b_sign0 = 4'd4; b_sign1 = 4'd16; b_sign2 = 4'd0; b_sign3 = 4'd15;
@(posedge clk_i);
a_mant0 = 8'd217; a_mant1 = 8'd228; a_mant2 = 8'd245; a_mant3 = 8'd198;
b_mant0 = 8'd77; b_mant1 = 8'd10; b_mant2 = 8'd249; b_mant3 = 8'd33;
a_exp0 = 10'd146; a_exp1 = 10'd859; a_exp2 = 10'd29; a_exp3 = 10'd404;
b_exp0 = 10'd508; b_exp1 = 10'd194; b_exp2 = 10'd314; b_exp3 = 10'd919;
a_sign0 = 4'd13; a_sign1 = 4'd12; a_sign2 = 4'd15; a_sign3 = 4'd0;
b_sign0 = 4'd13; b_sign1 = 4'd6; b_sign2 = 4'd12; b_sign3 = 4'd8;
@(posedge clk_i);
shared_exps0 = 8'd97;
shared_exps1 = 8'd100;
a_mant0 = 8'd4; a_mant1 = 8'd209; a_mant2 = 8'd41; a_mant3 = 8'd246;
b_mant0 = 8'd50; b_mant1 = 8'd44; b_mant2 = 8'd208; b_mant3 = 8'd169;
a_exp0 = 10'd366; a_exp1 = 10'd269; a_exp2 = 10'd274; a_exp3 = 10'd149;
b_exp0 = 10'd691; b_exp1 = 10'd60; b_exp2 = 10'd526; b_exp3 = 10'd277;
a_sign0 = 4'd7; a_sign1 = 4'd14; a_sign2 = 4'd12; a_sign3 = 4'd9;
b_sign0 = 4'd10; b_sign1 = 4'd8; b_sign2 = 4'd2; b_sign3 = 4'd14;
@(posedge clk_i);
a_mant0 = 8'd92; a_mant1 = 8'd159; a_mant2 = 8'd212; a_mant3 = 8'd214;
b_mant0 = 8'd238; b_mant1 = 8'd79; b_mant2 = 8'd182; b_mant3 = 8'd176;
a_exp0 = 10'd144; a_exp1 = 10'd535; a_exp2 = 10'd839; a_exp3 = 10'd626;
b_exp0 = 10'd954; b_exp1 = 10'd733; b_exp2 = 10'd554; b_exp3 = 10'd782;
a_sign0 = 4'd8; a_sign1 = 4'd3; a_sign2 = 4'd15; a_sign3 = 4'd16;
b_sign0 = 4'd16; b_sign1 = 4'd11; b_sign2 = 4'd10; b_sign3 = 4'd11;
@(posedge clk_i);
a_mant0 = 8'd100; a_mant1 = 8'd84; a_mant2 = 8'd252; a_mant3 = 8'd140;
b_mant0 = 8'd222; b_mant1 = 8'd243; b_mant2 = 8'd152; b_mant3 = 8'd241;
a_exp0 = 10'd166; a_exp1 = 10'd165; a_exp2 = 10'd693; a_exp3 = 10'd414;
b_exp0 = 10'd347; b_exp1 = 10'd829; b_exp2 = 10'd0; b_exp3 = 10'd992;
a_sign0 = 4'd6; a_sign1 = 4'd14; a_sign2 = 4'd14; a_sign3 = 4'd12;
b_sign0 = 4'd12; b_sign1 = 4'd0; b_sign2 = 4'd6; b_sign3 = 4'd15;
@(posedge clk_i);
a_mant0 = 8'd45; a_mant1 = 8'd59; a_mant2 = 8'd176; a_mant3 = 8'd41;
b_mant0 = 8'd27; b_mant1 = 8'd134; b_mant2 = 8'd76; b_mant3 = 8'd210;
a_exp0 = 10'd683; a_exp1 = 10'd154; a_exp2 = 10'd476; a_exp3 = 10'd411;
b_exp0 = 10'd729; b_exp1 = 10'd46; b_exp2 = 10'd819; b_exp3 = 10'd665;
a_sign0 = 4'd15; a_sign1 = 4'd0; a_sign2 = 4'd10; a_sign3 = 4'd15;
b_sign0 = 4'd13; b_sign1 = 4'd8; b_sign2 = 4'd2; b_sign3 = 4'd6;
@(posedge clk_i);
a_mant0 = 8'd148; a_mant1 = 8'd161; a_mant2 = 8'd220; a_mant3 = 8'd181;
b_mant0 = 8'd72; b_mant1 = 8'd241; b_mant2 = 8'd236; b_mant3 = 8'd185;
a_exp0 = 10'd416; a_exp1 = 10'd929; a_exp2 = 10'd316; a_exp3 = 10'd449;
b_exp0 = 10'd968; b_exp1 = 10'd760; b_exp2 = 10'd964; b_exp3 = 10'd639;
a_sign0 = 4'd7; a_sign1 = 4'd7; a_sign2 = 4'd3; a_sign3 = 4'd3;
b_sign0 = 4'd13; b_sign1 = 4'd12; b_sign2 = 4'd16; b_sign3 = 4'd16;
@(posedge clk_i);
a_mant0 = 8'd239; a_mant1 = 8'd1; a_mant2 = 8'd159; a_mant3 = 8'd245;
b_mant0 = 8'd10; b_mant1 = 8'd140; b_mant2 = 8'd105; b_mant3 = 8'd210;
a_exp0 = 10'd555; a_exp1 = 10'd534; a_exp2 = 10'd164; a_exp3 = 10'd438;
b_exp0 = 10'd761; b_exp1 = 10'd777; b_exp2 = 10'd12; b_exp3 = 10'd585;
a_sign0 = 4'd9; a_sign1 = 4'd6; a_sign2 = 4'd7; a_sign3 = 4'd0;
b_sign0 = 4'd14; b_sign1 = 4'd4; b_sign2 = 4'd11; b_sign3 = 4'd15;
@(posedge clk_i);
a_mant0 = 8'd32; a_mant1 = 8'd24; a_mant2 = 8'd35; a_mant3 = 8'd90;
b_mant0 = 8'd44; b_mant1 = 8'd248; b_mant2 = 8'd253; b_mant3 = 8'd90;
a_exp0 = 10'd370; a_exp1 = 10'd613; a_exp2 = 10'd291; a_exp3 = 10'd875;
b_exp0 = 10'd1017; b_exp1 = 10'd6; b_exp2 = 10'd290; b_exp3 = 10'd676;
a_sign0 = 4'd6; a_sign1 = 4'd5; a_sign2 = 4'd2; a_sign3 = 4'd7;
b_sign0 = 4'd2; b_sign1 = 4'd7; b_sign2 = 4'd6; b_sign3 = 4'd1;
@(posedge clk_i);
a_mant0 = 8'd40; a_mant1 = 8'd113; a_mant2 = 8'd165; a_mant3 = 8'd246;
b_mant0 = 8'd11; b_mant1 = 8'd58; b_mant2 = 8'd167; b_mant3 = 8'd202;
a_exp0 = 10'd917; a_exp1 = 10'd522; a_exp2 = 10'd472; a_exp3 = 10'd104;
b_exp0 = 10'd718; b_exp1 = 10'd71; b_exp2 = 10'd214; b_exp3 = 10'd802;
a_sign0 = 4'd10; a_sign1 = 4'd11; a_sign2 = 4'd3; a_sign3 = 4'd16;
b_sign0 = 4'd4; b_sign1 = 4'd6; b_sign2 = 4'd6; b_sign3 = 4'd15;
@(posedge clk_i);
shared_exps0 = 8'd127;
shared_exps1 = 8'd112;
a_mant0 = 8'd49; a_mant1 = 8'd195; a_mant2 = 8'd123; a_mant3 = 8'd111;
b_mant0 = 8'd202; b_mant1 = 8'd97; b_mant2 = 8'd76; b_mant3 = 8'd39;
a_exp0 = 10'd303; a_exp1 = 10'd810; a_exp2 = 10'd29; a_exp3 = 10'd21;
b_exp0 = 10'd713; b_exp1 = 10'd353; b_exp2 = 10'd703; b_exp3 = 10'd646;
a_sign0 = 4'd2; a_sign1 = 4'd16; a_sign2 = 4'd13; a_sign3 = 4'd14;
b_sign0 = 4'd1; b_sign1 = 4'd6; b_sign2 = 4'd9; b_sign3 = 4'd14;
@(posedge clk_i);
a_mant0 = 8'd215; a_mant1 = 8'd79; a_mant2 = 8'd82; a_mant3 = 8'd175;
b_mant0 = 8'd9; b_mant1 = 8'd3; b_mant2 = 8'd174; b_mant3 = 8'd192;
a_exp0 = 10'd706; a_exp1 = 10'd624; a_exp2 = 10'd552; a_exp3 = 10'd693;
b_exp0 = 10'd776; b_exp1 = 10'd815; b_exp2 = 10'd745; b_exp3 = 10'd484;
a_sign0 = 4'd13; a_sign1 = 4'd16; a_sign2 = 4'd1; a_sign3 = 4'd13;
b_sign0 = 4'd2; b_sign1 = 4'd10; b_sign2 = 4'd3; b_sign3 = 4'd13;
@(posedge clk_i);
a_mant0 = 8'd51; a_mant1 = 8'd74; a_mant2 = 8'd49; a_mant3 = 8'd174;
b_mant0 = 8'd115; b_mant1 = 8'd71; b_mant2 = 8'd210; b_mant3 = 8'd109;
a_exp0 = 10'd582; a_exp1 = 10'd929; a_exp2 = 10'd875; a_exp3 = 10'd726;
b_exp0 = 10'd478; b_exp1 = 10'd575; b_exp2 = 10'd788; b_exp3 = 10'd639;
a_sign0 = 4'd9; a_sign1 = 4'd14; a_sign2 = 4'd8; a_sign3 = 4'd16;
b_sign0 = 4'd4; b_sign1 = 4'd10; b_sign2 = 4'd10; b_sign3 = 4'd5;
@(posedge clk_i);
a_mant0 = 8'd19; a_mant1 = 8'd178; a_mant2 = 8'd220; a_mant3 = 8'd198;
b_mant0 = 8'd126; b_mant1 = 8'd249; b_mant2 = 8'd33; b_mant3 = 8'd44;
a_exp0 = 10'd223; a_exp1 = 10'd556; a_exp2 = 10'd709; a_exp3 = 10'd287;
b_exp0 = 10'd772; b_exp1 = 10'd316; b_exp2 = 10'd182; b_exp3 = 10'd58;
a_sign0 = 4'd15; a_sign1 = 4'd10; a_sign2 = 4'd13; a_sign3 = 4'd13;
b_sign0 = 4'd15; b_sign1 = 4'd10; b_sign2 = 4'd10; b_sign3 = 4'd7;
@(posedge clk_i);
a_mant0 = 8'd60; a_mant1 = 8'd182; a_mant2 = 8'd87; a_mant3 = 8'd205;
b_mant0 = 8'd18; b_mant1 = 8'd115; b_mant2 = 8'd233; b_mant3 = 8'd65;
a_exp0 = 10'd590; a_exp1 = 10'd331; a_exp2 = 10'd406; a_exp3 = 10'd331;
b_exp0 = 10'd732; b_exp1 = 10'd454; b_exp2 = 10'd371; b_exp3 = 10'd226;
a_sign0 = 4'd3; a_sign1 = 4'd0; a_sign2 = 4'd14; a_sign3 = 4'd14;
b_sign0 = 4'd9; b_sign1 = 4'd3; b_sign2 = 4'd7; b_sign3 = 4'd4;
@(posedge clk_i);
a_mant0 = 8'd81; a_mant1 = 8'd3; a_mant2 = 8'd133; a_mant3 = 8'd252;
b_mant0 = 8'd130; b_mant1 = 8'd186; b_mant2 = 8'd67; b_mant3 = 8'd130;
a_exp0 = 10'd447; a_exp1 = 10'd436; a_exp2 = 10'd1015; a_exp3 = 10'd962;
b_exp0 = 10'd582; b_exp1 = 10'd373; b_exp2 = 10'd787; b_exp3 = 10'd1016;
a_sign0 = 4'd6; a_sign1 = 4'd11; a_sign2 = 4'd13; a_sign3 = 4'd2;
b_sign0 = 4'd14; b_sign1 = 4'd13; b_sign2 = 4'd10; b_sign3 = 4'd7;
@(posedge clk_i);
a_mant0 = 8'd182; a_mant1 = 8'd142; a_mant2 = 8'd124; a_mant3 = 8'd182;
b_mant0 = 8'd76; b_mant1 = 8'd132; b_mant2 = 8'd113; b_mant3 = 8'd60;
a_exp0 = 10'd13; a_exp1 = 10'd945; a_exp2 = 10'd352; a_exp3 = 10'd530;
b_exp0 = 10'd491; b_exp1 = 10'd308; b_exp2 = 10'd323; b_exp3 = 10'd385;
a_sign0 = 4'd2; a_sign1 = 4'd13; a_sign2 = 4'd14; a_sign3 = 4'd1;
b_sign0 = 4'd16; b_sign1 = 4'd13; b_sign2 = 4'd12; b_sign3 = 4'd7;
@(posedge clk_i);
a_mant0 = 8'd38; a_mant1 = 8'd79; a_mant2 = 8'd213; a_mant3 = 8'd39;
b_mant0 = 8'd80; b_mant1 = 8'd159; b_mant2 = 8'd114; b_mant3 = 8'd241;
a_exp0 = 10'd695; a_exp1 = 10'd662; a_exp2 = 10'd588; a_exp3 = 10'd661;
b_exp0 = 10'd591; b_exp1 = 10'd472; b_exp2 = 10'd672; b_exp3 = 10'd434;
a_sign0 = 4'd8; a_sign1 = 4'd8; a_sign2 = 4'd9; a_sign3 = 4'd12;
b_sign0 = 4'd1; b_sign1 = 4'd8; b_sign2 = 4'd16; b_sign3 = 4'd8;
@(posedge clk_i);
shared_exps0 = 8'd116;
shared_exps1 = 8'd130;
rstn = 0;
@(posedge clk_i);
rstn = 1;
a_mant0 = 8'd0; a_mant1 = 8'd171; a_mant2 = 8'd213; a_mant3 = 8'd145;
b_mant0 = 8'd96; b_mant1 = 8'd129; b_mant2 = 8'd68; b_mant3 = 8'd117;
a_exp0 = 10'd241; a_exp1 = 10'd200; a_exp2 = 10'd261; a_exp3 = 10'd261;
b_exp0 = 10'd642; b_exp1 = 10'd176; b_exp2 = 10'd519; b_exp3 = 10'd322;
a_sign0 = 4'd6; a_sign1 = 4'd15; a_sign2 = 4'd6; a_sign3 = 4'd7;
b_sign0 = 4'd1; b_sign1 = 4'd6; b_sign2 = 4'd16; b_sign3 = 4'd13;
@(posedge clk_i);
a_mant0 = 8'd50; a_mant1 = 8'd97; a_mant2 = 8'd222; a_mant3 = 8'd149;
b_mant0 = 8'd171; b_mant1 = 8'd71; b_mant2 = 8'd74; b_mant3 = 8'd52;
a_exp0 = 10'd415; a_exp1 = 10'd272; a_exp2 = 10'd806; a_exp3 = 10'd208;
b_exp0 = 10'd430; b_exp1 = 10'd513; b_exp2 = 10'd168; b_exp3 = 10'd238;
a_sign0 = 4'd2; a_sign1 = 4'd5; a_sign2 = 4'd15; a_sign3 = 4'd11;
b_sign0 = 4'd3; b_sign1 = 4'd0; b_sign2 = 4'd11; b_sign3 = 4'd12;
@(posedge clk_i);
a_mant0 = 8'd214; a_mant1 = 8'd163; a_mant2 = 8'd61; a_mant3 = 8'd144;
b_mant0 = 8'd217; b_mant1 = 8'd12; b_mant2 = 8'd148; b_mant3 = 8'd155;
a_exp0 = 10'd756; a_exp1 = 10'd206; a_exp2 = 10'd326; a_exp3 = 10'd553;
b_exp0 = 10'd193; b_exp1 = 10'd944; b_exp2 = 10'd821; b_exp3 = 10'd117;
a_sign0 = 4'd5; a_sign1 = 4'd3; a_sign2 = 4'd15; a_sign3 = 4'd5;
b_sign0 = 4'd15; b_sign1 = 4'd7; b_sign2 = 4'd3; b_sign3 = 4'd7;
@(posedge clk_i);
a_mant0 = 8'd20; a_mant1 = 8'd246; a_mant2 = 8'd67; a_mant3 = 8'd117;
b_mant0 = 8'd28; b_mant1 = 8'd35; b_mant2 = 8'd243; b_mant3 = 8'd186;
a_exp0 = 10'd565; a_exp1 = 10'd66; a_exp2 = 10'd564; a_exp3 = 10'd621;
b_exp0 = 10'd776; b_exp1 = 10'd731; b_exp2 = 10'd671; b_exp3 = 10'd328;
a_sign0 = 4'd8; a_sign1 = 4'd4; a_sign2 = 4'd0; a_sign3 = 4'd9;
b_sign0 = 4'd10; b_sign1 = 4'd15; b_sign2 = 4'd13; b_sign3 = 4'd13;
@(posedge clk_i);
a_mant0 = 8'd77; a_mant1 = 8'd166; a_mant2 = 8'd28; a_mant3 = 8'd21;
b_mant0 = 8'd119; b_mant1 = 8'd145; b_mant2 = 8'd185; b_mant3 = 8'd155;
a_exp0 = 10'd629; a_exp1 = 10'd546; a_exp2 = 10'd345; a_exp3 = 10'd181;
b_exp0 = 10'd365; b_exp1 = 10'd111; b_exp2 = 10'd599; b_exp3 = 10'd812;
a_sign0 = 4'd10; a_sign1 = 4'd10; a_sign2 = 4'd11; a_sign3 = 4'd1;
b_sign0 = 4'd8; b_sign1 = 4'd1; b_sign2 = 4'd0; b_sign3 = 4'd13;
@(posedge clk_i);
a_mant0 = 8'd128; a_mant1 = 8'd12; a_mant2 = 8'd51; a_mant3 = 8'd104;
b_mant0 = 8'd178; b_mant1 = 8'd242; b_mant2 = 8'd8; b_mant3 = 8'd156;
a_exp0 = 10'd612; a_exp1 = 10'd200; a_exp2 = 10'd611; a_exp3 = 10'd580;
b_exp0 = 10'd829; b_exp1 = 10'd982; b_exp2 = 10'd89; b_exp3 = 10'd534;
a_sign0 = 4'd3; a_sign1 = 4'd2; a_sign2 = 4'd8; a_sign3 = 4'd11;
b_sign0 = 4'd14; b_sign1 = 4'd16; b_sign2 = 4'd12; b_sign3 = 4'd11;
@(posedge clk_i);
a_mant0 = 8'd75; a_mant1 = 8'd209; a_mant2 = 8'd27; a_mant3 = 8'd2;
b_mant0 = 8'd11; b_mant1 = 8'd7; b_mant2 = 8'd207; b_mant3 = 8'd6;
a_exp0 = 10'd378; a_exp1 = 10'd216; a_exp2 = 10'd751; a_exp3 = 10'd56;
b_exp0 = 10'd753; b_exp1 = 10'd373; b_exp2 = 10'd544; b_exp3 = 10'd715;
a_sign0 = 4'd15; a_sign1 = 4'd13; a_sign2 = 4'd14; a_sign3 = 4'd10;
b_sign0 = 4'd10; b_sign1 = 4'd11; b_sign2 = 4'd7; b_sign3 = 4'd7;
@(posedge clk_i);
shared_exps0 = 8'd149;
shared_exps1 = 8'd126;
a_mant0 = 8'd207; a_mant1 = 8'd4; a_mant2 = 8'd90; a_mant3 = 8'd152;
b_mant0 = 8'd79; b_mant1 = 8'd13; b_mant2 = 8'd255; b_mant3 = 8'd112;
a_exp0 = 10'd253; a_exp1 = 10'd368; a_exp2 = 10'd643; a_exp3 = 10'd497;
b_exp0 = 10'd946; b_exp1 = 10'd121; b_exp2 = 10'd63; b_exp3 = 10'd33;
a_sign0 = 4'd9; a_sign1 = 4'd12; a_sign2 = 4'd16; a_sign3 = 4'd3;
b_sign0 = 4'd9; b_sign1 = 4'd6; b_sign2 = 4'd0; b_sign3 = 4'd7;
@(posedge clk_i);
a_mant0 = 8'd9; a_mant1 = 8'd11; a_mant2 = 8'd159; a_mant3 = 8'd229;
b_mant0 = 8'd36; b_mant1 = 8'd119; b_mant2 = 8'd171; b_mant3 = 8'd143;
a_exp0 = 10'd132; a_exp1 = 10'd29; a_exp2 = 10'd824; a_exp3 = 10'd727;
b_exp0 = 10'd155; b_exp1 = 10'd15; b_exp2 = 10'd445; b_exp3 = 10'd732;
a_sign0 = 4'd6; a_sign1 = 4'd6; a_sign2 = 4'd2; a_sign3 = 4'd7;
b_sign0 = 4'd2; b_sign1 = 4'd3; b_sign2 = 4'd1; b_sign3 = 4'd13;
@(posedge clk_i);
a_mant0 = 8'd183; a_mant1 = 8'd46; a_mant2 = 8'd163; a_mant3 = 8'd33;
b_mant0 = 8'd138; b_mant1 = 8'd206; b_mant2 = 8'd107; b_mant3 = 8'd112;
a_exp0 = 10'd366; a_exp1 = 10'd783; a_exp2 = 10'd917; a_exp3 = 10'd542;
b_exp0 = 10'd348; b_exp1 = 10'd352; b_exp2 = 10'd503; b_exp3 = 10'd832;
a_sign0 = 4'd0; a_sign1 = 4'd8; a_sign2 = 4'd11; a_sign3 = 4'd14;
b_sign0 = 4'd12; b_sign1 = 4'd11; b_sign2 = 4'd15; b_sign3 = 4'd13;
@(posedge clk_i);
a_mant0 = 8'd56; a_mant1 = 8'd191; a_mant2 = 8'd230; a_mant3 = 8'd57;
b_mant0 = 8'd150; b_mant1 = 8'd172; b_mant2 = 8'd192; b_mant3 = 8'd112;
a_exp0 = 10'd151; a_exp1 = 10'd754; a_exp2 = 10'd580; a_exp3 = 10'd577;
b_exp0 = 10'd140; b_exp1 = 10'd454; b_exp2 = 10'd532; b_exp3 = 10'd940;
a_sign0 = 4'd9; a_sign1 = 4'd0; a_sign2 = 4'd5; a_sign3 = 4'd10;
b_sign0 = 4'd11; b_sign1 = 4'd9; b_sign2 = 4'd14; b_sign3 = 4'd14;
@(posedge clk_i);
a_mant0 = 8'd115; a_mant1 = 8'd45; a_mant2 = 8'd3; a_mant3 = 8'd252;
b_mant0 = 8'd154; b_mant1 = 8'd64; b_mant2 = 8'd52; b_mant3 = 8'd192;
a_exp0 = 10'd123; a_exp1 = 10'd787; a_exp2 = 10'd601; a_exp3 = 10'd443;
b_exp0 = 10'd256; b_exp1 = 10'd709; b_exp2 = 10'd362; b_exp3 = 10'd734;
a_sign0 = 4'd16; a_sign1 = 4'd4; a_sign2 = 4'd6; a_sign3 = 4'd11;
b_sign0 = 4'd14; b_sign1 = 4'd4; b_sign2 = 4'd0; b_sign3 = 4'd2;
@(posedge clk_i);
a_mant0 = 8'd217; a_mant1 = 8'd242; a_mant2 = 8'd14; a_mant3 = 8'd137;
b_mant0 = 8'd80; b_mant1 = 8'd178; b_mant2 = 8'd146; b_mant3 = 8'd22;
a_exp0 = 10'd382; a_exp1 = 10'd888; a_exp2 = 10'd380; a_exp3 = 10'd90;
b_exp0 = 10'd501; b_exp1 = 10'd229; b_exp2 = 10'd894; b_exp3 = 10'd683;
a_sign0 = 4'd10; a_sign1 = 4'd4; a_sign2 = 4'd14; a_sign3 = 4'd13;
b_sign0 = 4'd6; b_sign1 = 4'd16; b_sign2 = 4'd1; b_sign3 = 4'd5;
@(posedge clk_i);
a_mant0 = 8'd179; a_mant1 = 8'd180; a_mant2 = 8'd5; a_mant3 = 8'd113;
b_mant0 = 8'd44; b_mant1 = 8'd132; b_mant2 = 8'd120; b_mant3 = 8'd183;
a_exp0 = 10'd599; a_exp1 = 10'd300; a_exp2 = 10'd737; a_exp3 = 10'd274;
b_exp0 = 10'd275; b_exp1 = 10'd399; b_exp2 = 10'd763; b_exp3 = 10'd183;
a_sign0 = 4'd15; a_sign1 = 4'd16; a_sign2 = 4'd6; a_sign3 = 4'd11;
b_sign0 = 4'd10; b_sign1 = 4'd9; b_sign2 = 4'd9; b_sign3 = 4'd4;
@(posedge clk_i);
a_mant0 = 8'd109; a_mant1 = 8'd33; a_mant2 = 8'd60; a_mant3 = 8'd39;
b_mant0 = 8'd240; b_mant1 = 8'd88; b_mant2 = 8'd196; b_mant3 = 8'd75;
a_exp0 = 10'd0; a_exp1 = 10'd289; a_exp2 = 10'd485; a_exp3 = 10'd653;
b_exp0 = 10'd351; b_exp1 = 10'd202; b_exp2 = 10'd820; b_exp3 = 10'd654;
a_sign0 = 4'd0; a_sign1 = 4'd3; a_sign2 = 4'd10; a_sign3 = 4'd10;
b_sign0 = 4'd10; b_sign1 = 4'd4; b_sign2 = 4'd6; b_sign3 = 4'd6;
@(posedge clk_i);
shared_exps0 = 8'd119;
shared_exps1 = 8'd127;
a_mant0 = 8'd126; a_mant1 = 8'd0; a_mant2 = 8'd119; a_mant3 = 8'd195;
b_mant0 = 8'd135; b_mant1 = 8'd163; b_mant2 = 8'd218; b_mant3 = 8'd210;
a_exp0 = 10'd547; a_exp1 = 10'd330; a_exp2 = 10'd298; a_exp3 = 10'd611;
b_exp0 = 10'd392; b_exp1 = 10'd992; b_exp2 = 10'd134; b_exp3 = 10'd7;
a_sign0 = 4'd0; a_sign1 = 4'd4; a_sign2 = 4'd4; a_sign3 = 4'd5;
b_sign0 = 4'd0; b_sign1 = 4'd9; b_sign2 = 4'd1; b_sign3 = 4'd10;
@(posedge clk_i);
a_mant0 = 8'd35; a_mant1 = 8'd226; a_mant2 = 8'd206; a_mant3 = 8'd150;
b_mant0 = 8'd146; b_mant1 = 8'd201; b_mant2 = 8'd26; b_mant3 = 8'd145;
a_exp0 = 10'd637; a_exp1 = 10'd664; a_exp2 = 10'd755; a_exp3 = 10'd50;
b_exp0 = 10'd35; b_exp1 = 10'd498; b_exp2 = 10'd364; b_exp3 = 10'd804;
a_sign0 = 4'd0; a_sign1 = 4'd3; a_sign2 = 4'd11; a_sign3 = 4'd6;
b_sign0 = 4'd14; b_sign1 = 4'd1; b_sign2 = 4'd2; b_sign3 = 4'd9;
@(posedge clk_i);
a_mant0 = 8'd67; a_mant1 = 8'd162; a_mant2 = 8'd255; a_mant3 = 8'd248;
b_mant0 = 8'd157; b_mant1 = 8'd104; b_mant2 = 8'd40; b_mant3 = 8'd172;
a_exp0 = 10'd910; a_exp1 = 10'd122; a_exp2 = 10'd254; a_exp3 = 10'd297;
b_exp0 = 10'd632; b_exp1 = 10'd173; b_exp2 = 10'd6; b_exp3 = 10'd560;
a_sign0 = 4'd11; a_sign1 = 4'd10; a_sign2 = 4'd4; a_sign3 = 4'd3;
b_sign0 = 4'd14; b_sign1 = 4'd12; b_sign2 = 4'd3; b_sign3 = 4'd14;
@(posedge clk_i);
a_mant0 = 8'd239; a_mant1 = 8'd12; a_mant2 = 8'd195; a_mant3 = 8'd162;
b_mant0 = 8'd187; b_mant1 = 8'd142; b_mant2 = 8'd101; b_mant3 = 8'd70;
a_exp0 = 10'd44; a_exp1 = 10'd930; a_exp2 = 10'd440; a_exp3 = 10'd637;
b_exp0 = 10'd422; b_exp1 = 10'd364; b_exp2 = 10'd213; b_exp3 = 10'd842;
a_sign0 = 4'd9; a_sign1 = 4'd11; a_sign2 = 4'd8; a_sign3 = 4'd10;
b_sign0 = 4'd13; b_sign1 = 4'd14; b_sign2 = 4'd5; b_sign3 = 4'd4;
@(posedge clk_i);
a_mant0 = 8'd162; a_mant1 = 8'd209; a_mant2 = 8'd253; a_mant3 = 8'd125;
b_mant0 = 8'd37; b_mant1 = 8'd18; b_mant2 = 8'd231; b_mant3 = 8'd31;
a_exp0 = 10'd1013; a_exp1 = 10'd796; a_exp2 = 10'd997; a_exp3 = 10'd362;
b_exp0 = 10'd311; b_exp1 = 10'd565; b_exp2 = 10'd692; b_exp3 = 10'd923;
a_sign0 = 4'd16; a_sign1 = 4'd12; a_sign2 = 4'd15; a_sign3 = 4'd14;
b_sign0 = 4'd8; b_sign1 = 4'd14; b_sign2 = 4'd3; b_sign3 = 4'd12;
@(posedge clk_i);
a_mant0 = 8'd240; a_mant1 = 8'd67; a_mant2 = 8'd182; a_mant3 = 8'd126;
b_mant0 = 8'd126; b_mant1 = 8'd105; b_mant2 = 8'd25; b_mant3 = 8'd57;
a_exp0 = 10'd37; a_exp1 = 10'd346; a_exp2 = 10'd234; a_exp3 = 10'd237;
b_exp0 = 10'd793; b_exp1 = 10'd640; b_exp2 = 10'd166; b_exp3 = 10'd454;
a_sign0 = 4'd9; a_sign1 = 4'd1; a_sign2 = 4'd14; a_sign3 = 4'd1;
b_sign0 = 4'd13; b_sign1 = 4'd5; b_sign2 = 4'd12; b_sign3 = 4'd3;
@(posedge clk_i);
a_mant0 = 8'd137; a_mant1 = 8'd9; a_mant2 = 8'd27; a_mant3 = 8'd1;
b_mant0 = 8'd228; b_mant1 = 8'd224; b_mant2 = 8'd117; b_mant3 = 8'd53;
a_exp0 = 10'd166; a_exp1 = 10'd265; a_exp2 = 10'd763; a_exp3 = 10'd690;
b_exp0 = 10'd483; b_exp1 = 10'd993; b_exp2 = 10'd981; b_exp3 = 10'd459;
a_sign0 = 4'd11; a_sign1 = 4'd16; a_sign2 = 4'd8; a_sign3 = 4'd5;
b_sign0 = 4'd14; b_sign1 = 4'd11; b_sign2 = 4'd0; b_sign3 = 4'd0;
@(posedge clk_i);
a_mant0 = 8'd99; a_mant1 = 8'd100; a_mant2 = 8'd229; a_mant3 = 8'd241;
b_mant0 = 8'd163; b_mant1 = 8'd179; b_mant2 = 8'd85; b_mant3 = 8'd254;
a_exp0 = 10'd781; a_exp1 = 10'd996; a_exp2 = 10'd841; a_exp3 = 10'd17;
b_exp0 = 10'd913; b_exp1 = 10'd140; b_exp2 = 10'd472; b_exp3 = 10'd1000;
a_sign0 = 4'd2; a_sign1 = 4'd8; a_sign2 = 4'd0; a_sign3 = 4'd3;
b_sign0 = 4'd11; b_sign1 = 4'd7; b_sign2 = 4'd10; b_sign3 = 4'd12;
@(posedge clk_i);
shared_exps0 = 8'd101;
shared_exps1 = 8'd146;
a_mant0 = 8'd227; a_mant1 = 8'd106; a_mant2 = 8'd143; a_mant3 = 8'd65;
b_mant0 = 8'd220; b_mant1 = 8'd105; b_mant2 = 8'd231; b_mant3 = 8'd135;
a_exp0 = 10'd975; a_exp1 = 10'd566; a_exp2 = 10'd293; a_exp3 = 10'd605;
b_exp0 = 10'd613; b_exp1 = 10'd930; b_exp2 = 10'd799; b_exp3 = 10'd293;
a_sign0 = 4'd11; a_sign1 = 4'd10; a_sign2 = 4'd16; a_sign3 = 4'd16;
b_sign0 = 4'd5; b_sign1 = 4'd5; b_sign2 = 4'd8; b_sign3 = 4'd3;
@(posedge clk_i);
a_mant0 = 8'd212; a_mant1 = 8'd225; a_mant2 = 8'd89; a_mant3 = 8'd234;
b_mant0 = 8'd12; b_mant1 = 8'd139; b_mant2 = 8'd88; b_mant3 = 8'd189;
a_exp0 = 10'd463; a_exp1 = 10'd643; a_exp2 = 10'd938; a_exp3 = 10'd610;
b_exp0 = 10'd668; b_exp1 = 10'd341; b_exp2 = 10'd964; b_exp3 = 10'd314;
a_sign0 = 4'd12; a_sign1 = 4'd10; a_sign2 = 4'd10; a_sign3 = 4'd4;
b_sign0 = 4'd16; b_sign1 = 4'd9; b_sign2 = 4'd9; b_sign3 = 4'd2;
@(posedge clk_i);
a_mant0 = 8'd21; a_mant1 = 8'd165; a_mant2 = 8'd3; a_mant3 = 8'd52;
b_mant0 = 8'd119; b_mant1 = 8'd63; b_mant2 = 8'd86; b_mant3 = 8'd130;
a_exp0 = 10'd544; a_exp1 = 10'd983; a_exp2 = 10'd1001; a_exp3 = 10'd912;
b_exp0 = 10'd277; b_exp1 = 10'd992; b_exp2 = 10'd919; b_exp3 = 10'd319;
a_sign0 = 4'd16; a_sign1 = 4'd9; a_sign2 = 4'd14; a_sign3 = 4'd6;
b_sign0 = 4'd10; b_sign1 = 4'd1; b_sign2 = 4'd11; b_sign3 = 4'd2;
@(posedge clk_i);
a_mant0 = 8'd75; a_mant1 = 8'd87; a_mant2 = 8'd216; a_mant3 = 8'd222;
b_mant0 = 8'd81; b_mant1 = 8'd149; b_mant2 = 8'd126; b_mant3 = 8'd66;
a_exp0 = 10'd138; a_exp1 = 10'd97; a_exp2 = 10'd260; a_exp3 = 10'd81;
b_exp0 = 10'd932; b_exp1 = 10'd834; b_exp2 = 10'd883; b_exp3 = 10'd375;
a_sign0 = 4'd10; a_sign1 = 4'd6; a_sign2 = 4'd10; a_sign3 = 4'd8;
b_sign0 = 4'd11; b_sign1 = 4'd10; b_sign2 = 4'd11; b_sign3 = 4'd3;
@(posedge clk_i);
a_mant0 = 8'd207; a_mant1 = 8'd14; a_mant2 = 8'd95; a_mant3 = 8'd133;
b_mant0 = 8'd43; b_mant1 = 8'd117; b_mant2 = 8'd238; b_mant3 = 8'd155;
a_exp0 = 10'd341; a_exp1 = 10'd1006; a_exp2 = 10'd436; a_exp3 = 10'd533;
b_exp0 = 10'd801; b_exp1 = 10'd660; b_exp2 = 10'd230; b_exp3 = 10'd262;
a_sign0 = 4'd3; a_sign1 = 4'd12; a_sign2 = 4'd8; a_sign3 = 4'd11;
b_sign0 = 4'd1; b_sign1 = 4'd10; b_sign2 = 4'd15; b_sign3 = 4'd13;
@(posedge clk_i);
a_mant0 = 8'd79; a_mant1 = 8'd53; a_mant2 = 8'd140; a_mant3 = 8'd13;
b_mant0 = 8'd46; b_mant1 = 8'd177; b_mant2 = 8'd6; b_mant3 = 8'd134;
a_exp0 = 10'd152; a_exp1 = 10'd420; a_exp2 = 10'd610; a_exp3 = 10'd486;
b_exp0 = 10'd880; b_exp1 = 10'd382; b_exp2 = 10'd250; b_exp3 = 10'd895;
a_sign0 = 4'd5; a_sign1 = 4'd7; a_sign2 = 4'd12; a_sign3 = 4'd13;
b_sign0 = 4'd4; b_sign1 = 4'd13; b_sign2 = 4'd13; b_sign3 = 4'd10;
@(posedge clk_i);
a_mant0 = 8'd88; a_mant1 = 8'd11; a_mant2 = 8'd166; a_mant3 = 8'd50;
b_mant0 = 8'd230; b_mant1 = 8'd98; b_mant2 = 8'd171; b_mant3 = 8'd6;
a_exp0 = 10'd41; a_exp1 = 10'd346; a_exp2 = 10'd274; a_exp3 = 10'd136;
b_exp0 = 10'd234; b_exp1 = 10'd151; b_exp2 = 10'd41; b_exp3 = 10'd822;
a_sign0 = 4'd2; a_sign1 = 4'd13; a_sign2 = 4'd3; a_sign3 = 4'd8;
b_sign0 = 4'd10; b_sign1 = 4'd6; b_sign2 = 4'd14; b_sign3 = 4'd11;
@(posedge clk_i);
a_mant0 = 8'd73; a_mant1 = 8'd255; a_mant2 = 8'd125; a_mant3 = 8'd57;
b_mant0 = 8'd31; b_mant1 = 8'd3; b_mant2 = 8'd172; b_mant3 = 8'd43;
a_exp0 = 10'd340; a_exp1 = 10'd371; a_exp2 = 10'd820; a_exp3 = 10'd762;
b_exp0 = 10'd48; b_exp1 = 10'd55; b_exp2 = 10'd216; b_exp3 = 10'd760;
a_sign0 = 4'd0; a_sign1 = 4'd9; a_sign2 = 4'd4; a_sign3 = 4'd1;
b_sign0 = 4'd12; b_sign1 = 4'd13; b_sign2 = 4'd4; b_sign3 = 4'd11;
@(posedge clk_i);
shared_exps0 = 8'd136;
shared_exps1 = 8'd121;
rstn = 0;
@(posedge clk_i);
rstn = 1;
a_mant0 = 8'd60; a_mant1 = 8'd95; a_mant2 = 8'd171; a_mant3 = 8'd131;
b_mant0 = 8'd39; b_mant1 = 8'd175; b_mant2 = 8'd133; b_mant3 = 8'd125;
a_exp0 = 10'd886; a_exp1 = 10'd192; a_exp2 = 10'd759; a_exp3 = 10'd732;
b_exp0 = 10'd963; b_exp1 = 10'd18; b_exp2 = 10'd746; b_exp3 = 10'd447;
a_sign0 = 4'd14; a_sign1 = 4'd1; a_sign2 = 4'd7; a_sign3 = 4'd11;
b_sign0 = 4'd0; b_sign1 = 4'd14; b_sign2 = 4'd11; b_sign3 = 4'd3;
@(posedge clk_i);
a_mant0 = 8'd205; a_mant1 = 8'd56; a_mant2 = 8'd33; a_mant3 = 8'd222;
b_mant0 = 8'd59; b_mant1 = 8'd252; b_mant2 = 8'd27; b_mant3 = 8'd47;
a_exp0 = 10'd619; a_exp1 = 10'd423; a_exp2 = 10'd286; a_exp3 = 10'd151;
b_exp0 = 10'd575; b_exp1 = 10'd606; b_exp2 = 10'd7; b_exp3 = 10'd580;
a_sign0 = 4'd11; a_sign1 = 4'd12; a_sign2 = 4'd13; a_sign3 = 4'd9;
b_sign0 = 4'd3; b_sign1 = 4'd14; b_sign2 = 4'd11; b_sign3 = 4'd5;
@(posedge clk_i);
a_mant0 = 8'd68; a_mant1 = 8'd145; a_mant2 = 8'd86; a_mant3 = 8'd21;
b_mant0 = 8'd23; b_mant1 = 8'd135; b_mant2 = 8'd19; b_mant3 = 8'd66;
a_exp0 = 10'd562; a_exp1 = 10'd146; a_exp2 = 10'd420; a_exp3 = 10'd925;
b_exp0 = 10'd218; b_exp1 = 10'd453; b_exp2 = 10'd345; b_exp3 = 10'd726;
a_sign0 = 4'd1; a_sign1 = 4'd6; a_sign2 = 4'd3; a_sign3 = 4'd16;
b_sign0 = 4'd7; b_sign1 = 4'd2; b_sign2 = 4'd4; b_sign3 = 4'd0;
@(posedge clk_i);
a_mant0 = 8'd71; a_mant1 = 8'd72; a_mant2 = 8'd226; a_mant3 = 8'd207;
b_mant0 = 8'd139; b_mant1 = 8'd47; b_mant2 = 8'd113; b_mant3 = 8'd234;
a_exp0 = 10'd204; a_exp1 = 10'd804; a_exp2 = 10'd142; a_exp3 = 10'd155;
b_exp0 = 10'd453; b_exp1 = 10'd119; b_exp2 = 10'd956; b_exp3 = 10'd302;
a_sign0 = 4'd3; a_sign1 = 4'd14; a_sign2 = 4'd1; a_sign3 = 4'd1;
b_sign0 = 4'd12; b_sign1 = 4'd0; b_sign2 = 4'd14; b_sign3 = 4'd3;
@(posedge clk_i);
a_mant0 = 8'd26; a_mant1 = 8'd78; a_mant2 = 8'd237; a_mant3 = 8'd94;
b_mant0 = 8'd151; b_mant1 = 8'd65; b_mant2 = 8'd239; b_mant3 = 8'd101;
a_exp0 = 10'd905; a_exp1 = 10'd43; a_exp2 = 10'd623; a_exp3 = 10'd743;
b_exp0 = 10'd36; b_exp1 = 10'd300; b_exp2 = 10'd539; b_exp3 = 10'd648;
a_sign0 = 4'd5; a_sign1 = 4'd15; a_sign2 = 4'd6; a_sign3 = 4'd6;
b_sign0 = 4'd11; b_sign1 = 4'd7; b_sign2 = 4'd0; b_sign3 = 4'd14;
@(posedge clk_i);
a_mant0 = 8'd45; a_mant1 = 8'd28; a_mant2 = 8'd29; a_mant3 = 8'd93;
b_mant0 = 8'd106; b_mant1 = 8'd202; b_mant2 = 8'd205; b_mant3 = 8'd188;
a_exp0 = 10'd950; a_exp1 = 10'd427; a_exp2 = 10'd111; a_exp3 = 10'd229;
b_exp0 = 10'd454; b_exp1 = 10'd453; b_exp2 = 10'd756; b_exp3 = 10'd989;
a_sign0 = 4'd10; a_sign1 = 4'd13; a_sign2 = 4'd14; a_sign3 = 4'd5;
b_sign0 = 4'd13; b_sign1 = 4'd12; b_sign2 = 4'd9; b_sign3 = 4'd15;
@(posedge clk_i);
a_mant0 = 8'd164; a_mant1 = 8'd190; a_mant2 = 8'd203; a_mant3 = 8'd141;
b_mant0 = 8'd243; b_mant1 = 8'd1; b_mant2 = 8'd103; b_mant3 = 8'd35;
a_exp0 = 10'd129; a_exp1 = 10'd95; a_exp2 = 10'd837; a_exp3 = 10'd114;
b_exp0 = 10'd595; b_exp1 = 10'd673; b_exp2 = 10'd67; b_exp3 = 10'd297;
a_sign0 = 4'd5; a_sign1 = 4'd7; a_sign2 = 4'd9; a_sign3 = 4'd5;
b_sign0 = 4'd8; b_sign1 = 4'd3; b_sign2 = 4'd13; b_sign3 = 4'd7;
@(posedge clk_i);
shared_exps0 = 8'd114;
shared_exps1 = 8'd127;
a_mant0 = 8'd51; a_mant1 = 8'd37; a_mant2 = 8'd228; a_mant3 = 8'd91;
b_mant0 = 8'd182; b_mant1 = 8'd70; b_mant2 = 8'd48; b_mant3 = 8'd55;
a_exp0 = 10'd78; a_exp1 = 10'd812; a_exp2 = 10'd377; a_exp3 = 10'd938;
b_exp0 = 10'd87; b_exp1 = 10'd376; b_exp2 = 10'd830; b_exp3 = 10'd317;
a_sign0 = 4'd0; a_sign1 = 4'd13; a_sign2 = 4'd9; a_sign3 = 4'd8;
b_sign0 = 4'd10; b_sign1 = 4'd6; b_sign2 = 4'd3; b_sign3 = 4'd14;
@(posedge clk_i);
a_mant0 = 8'd71; a_mant1 = 8'd56; a_mant2 = 8'd190; a_mant3 = 8'd223;
b_mant0 = 8'd197; b_mant1 = 8'd228; b_mant2 = 8'd146; b_mant3 = 8'd187;
a_exp0 = 10'd510; a_exp1 = 10'd742; a_exp2 = 10'd126; a_exp3 = 10'd327;
b_exp0 = 10'd63; b_exp1 = 10'd550; b_exp2 = 10'd509; b_exp3 = 10'd507;
a_sign0 = 4'd9; a_sign1 = 4'd0; a_sign2 = 4'd0; a_sign3 = 4'd11;
b_sign0 = 4'd9; b_sign1 = 4'd1; b_sign2 = 4'd5; b_sign3 = 4'd15;
@(posedge clk_i);
a_mant0 = 8'd60; a_mant1 = 8'd160; a_mant2 = 8'd236; a_mant3 = 8'd82;
b_mant0 = 8'd143; b_mant1 = 8'd90; b_mant2 = 8'd157; b_mant3 = 8'd210;
a_exp0 = 10'd687; a_exp1 = 10'd868; a_exp2 = 10'd426; a_exp3 = 10'd722;
b_exp0 = 10'd581; b_exp1 = 10'd291; b_exp2 = 10'd921; b_exp3 = 10'd573;
a_sign0 = 4'd14; a_sign1 = 4'd3; a_sign2 = 4'd11; a_sign3 = 4'd2;
b_sign0 = 4'd7; b_sign1 = 4'd16; b_sign2 = 4'd4; b_sign3 = 4'd12;
@(posedge clk_i);
a_mant0 = 8'd238; a_mant1 = 8'd232; a_mant2 = 8'd251; a_mant3 = 8'd189;
b_mant0 = 8'd66; b_mant1 = 8'd203; b_mant2 = 8'd78; b_mant3 = 8'd126;
a_exp0 = 10'd207; a_exp1 = 10'd221; a_exp2 = 10'd37; a_exp3 = 10'd99;
b_exp0 = 10'd521; b_exp1 = 10'd770; b_exp2 = 10'd916; b_exp3 = 10'd792;
a_sign0 = 4'd5; a_sign1 = 4'd14; a_sign2 = 4'd6; a_sign3 = 4'd15;
b_sign0 = 4'd3; b_sign1 = 4'd2; b_sign2 = 4'd11; b_sign3 = 4'd7;
@(posedge clk_i);
a_mant0 = 8'd117; a_mant1 = 8'd131; a_mant2 = 8'd202; a_mant3 = 8'd74;
b_mant0 = 8'd157; b_mant1 = 8'd224; b_mant2 = 8'd112; b_mant3 = 8'd17;
a_exp0 = 10'd437; a_exp1 = 10'd539; a_exp2 = 10'd216; a_exp3 = 10'd452;
b_exp0 = 10'd297; b_exp1 = 10'd812; b_exp2 = 10'd255; b_exp3 = 10'd336;
a_sign0 = 4'd10; a_sign1 = 4'd10; a_sign2 = 4'd4; a_sign3 = 4'd2;
b_sign0 = 4'd15; b_sign1 = 4'd15; b_sign2 = 4'd5; b_sign3 = 4'd3;
@(posedge clk_i);
a_mant0 = 8'd60; a_mant1 = 8'd41; a_mant2 = 8'd167; a_mant3 = 8'd174;
b_mant0 = 8'd7; b_mant1 = 8'd142; b_mant2 = 8'd150; b_mant3 = 8'd32;
a_exp0 = 10'd1001; a_exp1 = 10'd230; a_exp2 = 10'd372; a_exp3 = 10'd83;
b_exp0 = 10'd559; b_exp1 = 10'd276; b_exp2 = 10'd639; b_exp3 = 10'd491;
a_sign0 = 4'd8; a_sign1 = 4'd14; a_sign2 = 4'd2; a_sign3 = 4'd13;
b_sign0 = 4'd10; b_sign1 = 4'd11; b_sign2 = 4'd13; b_sign3 = 4'd1;
@(posedge clk_i);
a_mant0 = 8'd107; a_mant1 = 8'd63; a_mant2 = 8'd148; a_mant3 = 8'd126;
b_mant0 = 8'd236; b_mant1 = 8'd191; b_mant2 = 8'd8; b_mant3 = 8'd4;
a_exp0 = 10'd762; a_exp1 = 10'd666; a_exp2 = 10'd207; a_exp3 = 10'd339;
b_exp0 = 10'd512; b_exp1 = 10'd859; b_exp2 = 10'd215; b_exp3 = 10'd650;
a_sign0 = 4'd3; a_sign1 = 4'd7; a_sign2 = 4'd4; a_sign3 = 4'd7;
b_sign0 = 4'd13; b_sign1 = 4'd8; b_sign2 = 4'd2; b_sign3 = 4'd10;
@(posedge clk_i);
a_mant0 = 8'd221; a_mant1 = 8'd11; a_mant2 = 8'd151; a_mant3 = 8'd3;
b_mant0 = 8'd90; b_mant1 = 8'd220; b_mant2 = 8'd86; b_mant3 = 8'd35;
a_exp0 = 10'd581; a_exp1 = 10'd865; a_exp2 = 10'd377; a_exp3 = 10'd16;
b_exp0 = 10'd225; b_exp1 = 10'd619; b_exp2 = 10'd175; b_exp3 = 10'd317;
a_sign0 = 4'd13; a_sign1 = 4'd16; a_sign2 = 4'd11; a_sign3 = 4'd14;
b_sign0 = 4'd16; b_sign1 = 4'd13; b_sign2 = 4'd4; b_sign3 = 4'd7;
@(posedge clk_i);
shared_exps0 = 8'd143;
shared_exps1 = 8'd117;
a_mant0 = 8'd247; a_mant1 = 8'd255; a_mant2 = 8'd244; a_mant3 = 8'd147;
b_mant0 = 8'd59; b_mant1 = 8'd3; b_mant2 = 8'd168; b_mant3 = 8'd86;
a_exp0 = 10'd320; a_exp1 = 10'd922; a_exp2 = 10'd6; a_exp3 = 10'd718;
b_exp0 = 10'd992; b_exp1 = 10'd387; b_exp2 = 10'd335; b_exp3 = 10'd141;
a_sign0 = 4'd8; a_sign1 = 4'd16; a_sign2 = 4'd15; a_sign3 = 4'd2;
b_sign0 = 4'd9; b_sign1 = 4'd5; b_sign2 = 4'd16; b_sign3 = 4'd1;
@(posedge clk_i);
a_mant0 = 8'd237; a_mant1 = 8'd120; a_mant2 = 8'd189; a_mant3 = 8'd54;
b_mant0 = 8'd194; b_mant1 = 8'd74; b_mant2 = 8'd188; b_mant3 = 8'd104;
a_exp0 = 10'd383; a_exp1 = 10'd537; a_exp2 = 10'd672; a_exp3 = 10'd959;
b_exp0 = 10'd604; b_exp1 = 10'd558; b_exp2 = 10'd609; b_exp3 = 10'd312;
a_sign0 = 4'd11; a_sign1 = 4'd4; a_sign2 = 4'd12; a_sign3 = 4'd7;
b_sign0 = 4'd4; b_sign1 = 4'd6; b_sign2 = 4'd12; b_sign3 = 4'd8;
@(posedge clk_i);
a_mant0 = 8'd9; a_mant1 = 8'd137; a_mant2 = 8'd189; a_mant3 = 8'd160;
b_mant0 = 8'd175; b_mant1 = 8'd15; b_mant2 = 8'd147; b_mant3 = 8'd230;
a_exp0 = 10'd719; a_exp1 = 10'd848; a_exp2 = 10'd534; a_exp3 = 10'd0;
b_exp0 = 10'd1022; b_exp1 = 10'd997; b_exp2 = 10'd566; b_exp3 = 10'd992;
a_sign0 = 4'd2; a_sign1 = 4'd13; a_sign2 = 4'd10; a_sign3 = 4'd0;
b_sign0 = 4'd2; b_sign1 = 4'd16; b_sign2 = 4'd8; b_sign3 = 4'd4;
@(posedge clk_i);
a_mant0 = 8'd248; a_mant1 = 8'd111; a_mant2 = 8'd83; a_mant3 = 8'd139;
b_mant0 = 8'd20; b_mant1 = 8'd200; b_mant2 = 8'd235; b_mant3 = 8'd171;
a_exp0 = 10'd11; a_exp1 = 10'd100; a_exp2 = 10'd329; a_exp3 = 10'd907;
b_exp0 = 10'd457; b_exp1 = 10'd978; b_exp2 = 10'd487; b_exp3 = 10'd4;
a_sign0 = 4'd7; a_sign1 = 4'd7; a_sign2 = 4'd9; a_sign3 = 4'd0;
b_sign0 = 4'd14; b_sign1 = 4'd10; b_sign2 = 4'd2; b_sign3 = 4'd13;
@(posedge clk_i);
a_mant0 = 8'd168; a_mant1 = 8'd16; a_mant2 = 8'd43; a_mant3 = 8'd94;
b_mant0 = 8'd18; b_mant1 = 8'd218; b_mant2 = 8'd217; b_mant3 = 8'd89;
a_exp0 = 10'd770; a_exp1 = 10'd959; a_exp2 = 10'd365; a_exp3 = 10'd733;
b_exp0 = 10'd885; b_exp1 = 10'd934; b_exp2 = 10'd985; b_exp3 = 10'd288;
a_sign0 = 4'd11; a_sign1 = 4'd9; a_sign2 = 4'd13; a_sign3 = 4'd9;
b_sign0 = 4'd14; b_sign1 = 4'd12; b_sign2 = 4'd12; b_sign3 = 4'd14;
@(posedge clk_i);
a_mant0 = 8'd127; a_mant1 = 8'd222; a_mant2 = 8'd199; a_mant3 = 8'd202;
b_mant0 = 8'd184; b_mant1 = 8'd162; b_mant2 = 8'd70; b_mant3 = 8'd122;
a_exp0 = 10'd765; a_exp1 = 10'd462; a_exp2 = 10'd870; a_exp3 = 10'd636;
b_exp0 = 10'd557; b_exp1 = 10'd563; b_exp2 = 10'd36; b_exp3 = 10'd712;
a_sign0 = 4'd3; a_sign1 = 4'd14; a_sign2 = 4'd10; a_sign3 = 4'd13;
b_sign0 = 4'd5; b_sign1 = 4'd14; b_sign2 = 4'd5; b_sign3 = 4'd6;
@(posedge clk_i);
a_mant0 = 8'd243; a_mant1 = 8'd87; a_mant2 = 8'd213; a_mant3 = 8'd13;
b_mant0 = 8'd237; b_mant1 = 8'd141; b_mant2 = 8'd59; b_mant3 = 8'd74;
a_exp0 = 10'd82; a_exp1 = 10'd102; a_exp2 = 10'd52; a_exp3 = 10'd304;
b_exp0 = 10'd536; b_exp1 = 10'd957; b_exp2 = 10'd160; b_exp3 = 10'd356;
a_sign0 = 4'd4; a_sign1 = 4'd8; a_sign2 = 4'd16; a_sign3 = 4'd3;
b_sign0 = 4'd15; b_sign1 = 4'd15; b_sign2 = 4'd15; b_sign3 = 4'd0;
@(posedge clk_i);
a_mant0 = 8'd111; a_mant1 = 8'd143; a_mant2 = 8'd73; a_mant3 = 8'd100;
b_mant0 = 8'd20; b_mant1 = 8'd227; b_mant2 = 8'd167; b_mant3 = 8'd101;
a_exp0 = 10'd509; a_exp1 = 10'd855; a_exp2 = 10'd848; a_exp3 = 10'd265;
b_exp0 = 10'd990; b_exp1 = 10'd826; b_exp2 = 10'd832; b_exp3 = 10'd756;
a_sign0 = 4'd11; a_sign1 = 4'd9; a_sign2 = 4'd15; a_sign3 = 4'd11;
b_sign0 = 4'd12; b_sign1 = 4'd12; b_sign2 = 4'd4; b_sign3 = 4'd15;
@(posedge clk_i);
shared_exps0 = 8'd110;
shared_exps1 = 8'd128;
a_mant0 = 8'd30; a_mant1 = 8'd183; a_mant2 = 8'd112; a_mant3 = 8'd152;
b_mant0 = 8'd72; b_mant1 = 8'd24; b_mant2 = 8'd134; b_mant3 = 8'd91;
a_exp0 = 10'd179; a_exp1 = 10'd861; a_exp2 = 10'd74; a_exp3 = 10'd130;
b_exp0 = 10'd41; b_exp1 = 10'd972; b_exp2 = 10'd105; b_exp3 = 10'd468;
a_sign0 = 4'd15; a_sign1 = 4'd15; a_sign2 = 4'd2; a_sign3 = 4'd13;
b_sign0 = 4'd7; b_sign1 = 4'd7; b_sign2 = 4'd3; b_sign3 = 4'd13;
@(posedge clk_i);
a_mant0 = 8'd220; a_mant1 = 8'd245; a_mant2 = 8'd145; a_mant3 = 8'd122;
b_mant0 = 8'd109; b_mant1 = 8'd126; b_mant2 = 8'd65; b_mant3 = 8'd138;
a_exp0 = 10'd197; a_exp1 = 10'd855; a_exp2 = 10'd756; a_exp3 = 10'd285;
b_exp0 = 10'd1015; b_exp1 = 10'd262; b_exp2 = 10'd881; b_exp3 = 10'd984;
a_sign0 = 4'd2; a_sign1 = 4'd8; a_sign2 = 4'd4; a_sign3 = 4'd9;
b_sign0 = 4'd9; b_sign1 = 4'd10; b_sign2 = 4'd0; b_sign3 = 4'd13;
@(posedge clk_i);
a_mant0 = 8'd111; a_mant1 = 8'd127; a_mant2 = 8'd253; a_mant3 = 8'd192;
b_mant0 = 8'd148; b_mant1 = 8'd68; b_mant2 = 8'd102; b_mant3 = 8'd182;
a_exp0 = 10'd707; a_exp1 = 10'd691; a_exp2 = 10'd147; a_exp3 = 10'd101;
b_exp0 = 10'd640; b_exp1 = 10'd253; b_exp2 = 10'd887; b_exp3 = 10'd501;
a_sign0 = 4'd10; a_sign1 = 4'd5; a_sign2 = 4'd15; a_sign3 = 4'd5;
b_sign0 = 4'd11; b_sign1 = 4'd6; b_sign2 = 4'd7; b_sign3 = 4'd7;
@(posedge clk_i);
a_mant0 = 8'd7; a_mant1 = 8'd242; a_mant2 = 8'd240; a_mant3 = 8'd117;
b_mant0 = 8'd208; b_mant1 = 8'd206; b_mant2 = 8'd24; b_mant3 = 8'd48;
a_exp0 = 10'd508; a_exp1 = 10'd648; a_exp2 = 10'd893; a_exp3 = 10'd992;
b_exp0 = 10'd738; b_exp1 = 10'd459; b_exp2 = 10'd933; b_exp3 = 10'd767;
a_sign0 = 4'd11; a_sign1 = 4'd4; a_sign2 = 4'd16; a_sign3 = 4'd1;
b_sign0 = 4'd5; b_sign1 = 4'd9; b_sign2 = 4'd14; b_sign3 = 4'd11;
@(posedge clk_i);
a_mant0 = 8'd228; a_mant1 = 8'd238; a_mant2 = 8'd34; a_mant3 = 8'd152;
b_mant0 = 8'd119; b_mant1 = 8'd125; b_mant2 = 8'd187; b_mant3 = 8'd138;
a_exp0 = 10'd454; a_exp1 = 10'd434; a_exp2 = 10'd974; a_exp3 = 10'd869;
b_exp0 = 10'd670; b_exp1 = 10'd691; b_exp2 = 10'd400; b_exp3 = 10'd1012;
a_sign0 = 4'd8; a_sign1 = 4'd4; a_sign2 = 4'd11; a_sign3 = 4'd16;
b_sign0 = 4'd9; b_sign1 = 4'd7; b_sign2 = 4'd5; b_sign3 = 4'd10;
@(posedge clk_i);
a_mant0 = 8'd31; a_mant1 = 8'd23; a_mant2 = 8'd212; a_mant3 = 8'd206;
b_mant0 = 8'd112; b_mant1 = 8'd158; b_mant2 = 8'd222; b_mant3 = 8'd44;
a_exp0 = 10'd1021; a_exp1 = 10'd45; a_exp2 = 10'd368; a_exp3 = 10'd205;
b_exp0 = 10'd644; b_exp1 = 10'd923; b_exp2 = 10'd618; b_exp3 = 10'd317;
a_sign0 = 4'd14; a_sign1 = 4'd12; a_sign2 = 4'd12; a_sign3 = 4'd16;
b_sign0 = 4'd4; b_sign1 = 4'd7; b_sign2 = 4'd7; b_sign3 = 4'd3;
@(posedge clk_i);
a_mant0 = 8'd61; a_mant1 = 8'd157; a_mant2 = 8'd128; a_mant3 = 8'd218;
b_mant0 = 8'd151; b_mant1 = 8'd225; b_mant2 = 8'd82; b_mant3 = 8'd225;
a_exp0 = 10'd542; a_exp1 = 10'd956; a_exp2 = 10'd153; a_exp3 = 10'd798;
b_exp0 = 10'd1014; b_exp1 = 10'd428; b_exp2 = 10'd275; b_exp3 = 10'd339;
a_sign0 = 4'd15; a_sign1 = 4'd10; a_sign2 = 4'd8; a_sign3 = 4'd11;
b_sign0 = 4'd16; b_sign1 = 4'd6; b_sign2 = 4'd5; b_sign3 = 4'd8;
@(posedge clk_i);
a_mant0 = 8'd83; a_mant1 = 8'd249; a_mant2 = 8'd21; a_mant3 = 8'd114;
b_mant0 = 8'd205; b_mant1 = 8'd39; b_mant2 = 8'd68; b_mant3 = 8'd133;
a_exp0 = 10'd727; a_exp1 = 10'd365; a_exp2 = 10'd558; a_exp3 = 10'd958;
b_exp0 = 10'd306; b_exp1 = 10'd725; b_exp2 = 10'd0; b_exp3 = 10'd412;
a_sign0 = 4'd12; a_sign1 = 4'd16; a_sign2 = 4'd12; a_sign3 = 4'd13;
b_sign0 = 4'd8; b_sign1 = 4'd9; b_sign2 = 4'd9; b_sign3 = 4'd3;
@(posedge clk_i);
shared_exps0 = 8'd107;
shared_exps1 = 8'd103;
rstn = 0;
@(posedge clk_i);
rstn = 1;
a_mant0 = 8'd44; a_mant1 = 8'd37; a_mant2 = 8'd50; a_mant3 = 8'd26;
b_mant0 = 8'd118; b_mant1 = 8'd224; b_mant2 = 8'd133; b_mant3 = 8'd50;
a_exp0 = 10'd165; a_exp1 = 10'd518; a_exp2 = 10'd731; a_exp3 = 10'd909;
b_exp0 = 10'd836; b_exp1 = 10'd166; b_exp2 = 10'd989; b_exp3 = 10'd350;
a_sign0 = 4'd14; a_sign1 = 4'd14; a_sign2 = 4'd1; a_sign3 = 4'd0;
b_sign0 = 4'd7; b_sign1 = 4'd2; b_sign2 = 4'd8; b_sign3 = 4'd1;
@(posedge clk_i);
a_mant0 = 8'd189; a_mant1 = 8'd147; a_mant2 = 8'd159; a_mant3 = 8'd153;
b_mant0 = 8'd94; b_mant1 = 8'd173; b_mant2 = 8'd125; b_mant3 = 8'd206;
a_exp0 = 10'd1012; a_exp1 = 10'd617; a_exp2 = 10'd63; a_exp3 = 10'd396;
b_exp0 = 10'd782; b_exp1 = 10'd596; b_exp2 = 10'd122; b_exp3 = 10'd671;
a_sign0 = 4'd0; a_sign1 = 4'd12; a_sign2 = 4'd9; a_sign3 = 4'd16;
b_sign0 = 4'd3; b_sign1 = 4'd1; b_sign2 = 4'd11; b_sign3 = 4'd15;
@(posedge clk_i);
a_mant0 = 8'd144; a_mant1 = 8'd137; a_mant2 = 8'd117; a_mant3 = 8'd223;
b_mant0 = 8'd105; b_mant1 = 8'd88; b_mant2 = 8'd229; b_mant3 = 8'd85;
a_exp0 = 10'd52; a_exp1 = 10'd250; a_exp2 = 10'd588; a_exp3 = 10'd116;
b_exp0 = 10'd843; b_exp1 = 10'd726; b_exp2 = 10'd673; b_exp3 = 10'd240;
a_sign0 = 4'd3; a_sign1 = 4'd15; a_sign2 = 4'd1; a_sign3 = 4'd1;
b_sign0 = 4'd14; b_sign1 = 4'd9; b_sign2 = 4'd13; b_sign3 = 4'd15;
@(posedge clk_i);
a_mant0 = 8'd116; a_mant1 = 8'd104; a_mant2 = 8'd49; a_mant3 = 8'd157;
b_mant0 = 8'd115; b_mant1 = 8'd205; b_mant2 = 8'd113; b_mant3 = 8'd84;
a_exp0 = 10'd102; a_exp1 = 10'd229; a_exp2 = 10'd557; a_exp3 = 10'd131;
b_exp0 = 10'd160; b_exp1 = 10'd521; b_exp2 = 10'd178; b_exp3 = 10'd910;
a_sign0 = 4'd3; a_sign1 = 4'd8; a_sign2 = 4'd9; a_sign3 = 4'd11;
b_sign0 = 4'd1; b_sign1 = 4'd2; b_sign2 = 4'd15; b_sign3 = 4'd8;
@(posedge clk_i);
a_mant0 = 8'd233; a_mant1 = 8'd221; a_mant2 = 8'd143; a_mant3 = 8'd199;
b_mant0 = 8'd89; b_mant1 = 8'd228; b_mant2 = 8'd228; b_mant3 = 8'd121;
a_exp0 = 10'd338; a_exp1 = 10'd780; a_exp2 = 10'd294; a_exp3 = 10'd740;
b_exp0 = 10'd485; b_exp1 = 10'd904; b_exp2 = 10'd410; b_exp3 = 10'd515;
a_sign0 = 4'd13; a_sign1 = 4'd13; a_sign2 = 4'd15; a_sign3 = 4'd11;
b_sign0 = 4'd4; b_sign1 = 4'd0; b_sign2 = 4'd13; b_sign3 = 4'd12;
@(posedge clk_i);
a_mant0 = 8'd4; a_mant1 = 8'd107; a_mant2 = 8'd210; a_mant3 = 8'd152;
b_mant0 = 8'd167; b_mant1 = 8'd163; b_mant2 = 8'd25; b_mant3 = 8'd127;
a_exp0 = 10'd412; a_exp1 = 10'd913; a_exp2 = 10'd114; a_exp3 = 10'd27;
b_exp0 = 10'd829; b_exp1 = 10'd399; b_exp2 = 10'd499; b_exp3 = 10'd307;
a_sign0 = 4'd10; a_sign1 = 4'd9; a_sign2 = 4'd15; a_sign3 = 4'd14;
b_sign0 = 4'd3; b_sign1 = 4'd10; b_sign2 = 4'd13; b_sign3 = 4'd16;
@(posedge clk_i);
a_mant0 = 8'd243; a_mant1 = 8'd3; a_mant2 = 8'd92; a_mant3 = 8'd209;
b_mant0 = 8'd37; b_mant1 = 8'd193; b_mant2 = 8'd242; b_mant3 = 8'd253;
a_exp0 = 10'd990; a_exp1 = 10'd178; a_exp2 = 10'd631; a_exp3 = 10'd421;
b_exp0 = 10'd184; b_exp1 = 10'd499; b_exp2 = 10'd374; b_exp3 = 10'd665;
a_sign0 = 4'd6; a_sign1 = 4'd7; a_sign2 = 4'd7; a_sign3 = 4'd8;
b_sign0 = 4'd1; b_sign1 = 4'd11; b_sign2 = 4'd1; b_sign3 = 4'd8;
@(posedge clk_i);
shared_exps0 = 8'd116;
shared_exps1 = 8'd132;
a_mant0 = 8'd31; a_mant1 = 8'd163; a_mant2 = 8'd0; a_mant3 = 8'd133;
b_mant0 = 8'd239; b_mant1 = 8'd63; b_mant2 = 8'd48; b_mant3 = 8'd162;
a_exp0 = 10'd966; a_exp1 = 10'd399; a_exp2 = 10'd390; a_exp3 = 10'd243;
b_exp0 = 10'd536; b_exp1 = 10'd306; b_exp2 = 10'd136; b_exp3 = 10'd576;
a_sign0 = 4'd16; a_sign1 = 4'd10; a_sign2 = 4'd4; a_sign3 = 4'd10;
b_sign0 = 4'd5; b_sign1 = 4'd0; b_sign2 = 4'd4; b_sign3 = 4'd8;
@(posedge clk_i);
a_mant0 = 8'd26; a_mant1 = 8'd188; a_mant2 = 8'd145; a_mant3 = 8'd228;
b_mant0 = 8'd64; b_mant1 = 8'd59; b_mant2 = 8'd135; b_mant3 = 8'd88;
a_exp0 = 10'd755; a_exp1 = 10'd464; a_exp2 = 10'd354; a_exp3 = 10'd676;
b_exp0 = 10'd689; b_exp1 = 10'd69; b_exp2 = 10'd769; b_exp3 = 10'd445;
a_sign0 = 4'd2; a_sign1 = 4'd4; a_sign2 = 4'd6; a_sign3 = 4'd8;
b_sign0 = 4'd12; b_sign1 = 4'd16; b_sign2 = 4'd12; b_sign3 = 4'd0;
@(posedge clk_i);
a_mant0 = 8'd99; a_mant1 = 8'd51; a_mant2 = 8'd135; a_mant3 = 8'd213;
b_mant0 = 8'd143; b_mant1 = 8'd45; b_mant2 = 8'd100; b_mant3 = 8'd117;
a_exp0 = 10'd494; a_exp1 = 10'd508; a_exp2 = 10'd997; a_exp3 = 10'd652;
b_exp0 = 10'd717; b_exp1 = 10'd225; b_exp2 = 10'd750; b_exp3 = 10'd344;
a_sign0 = 4'd4; a_sign1 = 4'd11; a_sign2 = 4'd5; a_sign3 = 4'd6;
b_sign0 = 4'd2; b_sign1 = 4'd9; b_sign2 = 4'd8; b_sign3 = 4'd1;
@(posedge clk_i);
a_mant0 = 8'd35; a_mant1 = 8'd19; a_mant2 = 8'd221; a_mant3 = 8'd200;
b_mant0 = 8'd149; b_mant1 = 8'd164; b_mant2 = 8'd97; b_mant3 = 8'd60;
a_exp0 = 10'd670; a_exp1 = 10'd363; a_exp2 = 10'd936; a_exp3 = 10'd311;
b_exp0 = 10'd887; b_exp1 = 10'd263; b_exp2 = 10'd930; b_exp3 = 10'd940;
a_sign0 = 4'd15; a_sign1 = 4'd12; a_sign2 = 4'd4; a_sign3 = 4'd12;
b_sign0 = 4'd14; b_sign1 = 4'd9; b_sign2 = 4'd1; b_sign3 = 4'd3;
@(posedge clk_i);
a_mant0 = 8'd119; a_mant1 = 8'd134; a_mant2 = 8'd159; a_mant3 = 8'd5;
b_mant0 = 8'd174; b_mant1 = 8'd216; b_mant2 = 8'd60; b_mant3 = 8'd27;
a_exp0 = 10'd141; a_exp1 = 10'd411; a_exp2 = 10'd778; a_exp3 = 10'd475;
b_exp0 = 10'd1017; b_exp1 = 10'd1015; b_exp2 = 10'd178; b_exp3 = 10'd732;
a_sign0 = 4'd2; a_sign1 = 4'd15; a_sign2 = 4'd1; a_sign3 = 4'd15;
b_sign0 = 4'd13; b_sign1 = 4'd2; b_sign2 = 4'd10; b_sign3 = 4'd12;
@(posedge clk_i);
a_mant0 = 8'd239; a_mant1 = 8'd179; a_mant2 = 8'd85; a_mant3 = 8'd152;
b_mant0 = 8'd224; b_mant1 = 8'd27; b_mant2 = 8'd75; b_mant3 = 8'd158;
a_exp0 = 10'd607; a_exp1 = 10'd170; a_exp2 = 10'd723; a_exp3 = 10'd90;
b_exp0 = 10'd254; b_exp1 = 10'd499; b_exp2 = 10'd157; b_exp3 = 10'd181;
a_sign0 = 4'd15; a_sign1 = 4'd14; a_sign2 = 4'd4; a_sign3 = 4'd9;
b_sign0 = 4'd9; b_sign1 = 4'd6; b_sign2 = 4'd16; b_sign3 = 4'd11;
@(posedge clk_i);
a_mant0 = 8'd163; a_mant1 = 8'd63; a_mant2 = 8'd227; a_mant3 = 8'd241;
b_mant0 = 8'd90; b_mant1 = 8'd62; b_mant2 = 8'd153; b_mant3 = 8'd9;
a_exp0 = 10'd181; a_exp1 = 10'd458; a_exp2 = 10'd454; a_exp3 = 10'd795;
b_exp0 = 10'd703; b_exp1 = 10'd448; b_exp2 = 10'd628; b_exp3 = 10'd926;
a_sign0 = 4'd0; a_sign1 = 4'd2; a_sign2 = 4'd12; a_sign3 = 4'd11;
b_sign0 = 4'd6; b_sign1 = 4'd8; b_sign2 = 4'd13; b_sign3 = 4'd0;
@(posedge clk_i);
a_mant0 = 8'd109; a_mant1 = 8'd28; a_mant2 = 8'd20; a_mant3 = 8'd18;
b_mant0 = 8'd17; b_mant1 = 8'd45; b_mant2 = 8'd30; b_mant3 = 8'd191;
a_exp0 = 10'd1002; a_exp1 = 10'd501; a_exp2 = 10'd5; a_exp3 = 10'd427;
b_exp0 = 10'd247; b_exp1 = 10'd539; b_exp2 = 10'd608; b_exp3 = 10'd573;
a_sign0 = 4'd5; a_sign1 = 4'd4; a_sign2 = 4'd12; a_sign3 = 4'd2;
b_sign0 = 4'd12; b_sign1 = 4'd7; b_sign2 = 4'd9; b_sign3 = 4'd14;
@(posedge clk_i);
shared_exps0 = 8'd121;
shared_exps1 = 8'd101;
a_mant0 = 8'd46; a_mant1 = 8'd175; a_mant2 = 8'd223; a_mant3 = 8'd181;
b_mant0 = 8'd66; b_mant1 = 8'd71; b_mant2 = 8'd159; b_mant3 = 8'd12;
a_exp0 = 10'd3; a_exp1 = 10'd11; a_exp2 = 10'd175; a_exp3 = 10'd131;
b_exp0 = 10'd309; b_exp1 = 10'd735; b_exp2 = 10'd70; b_exp3 = 10'd203;
a_sign0 = 4'd14; a_sign1 = 4'd6; a_sign2 = 4'd7; a_sign3 = 4'd16;
b_sign0 = 4'd10; b_sign1 = 4'd9; b_sign2 = 4'd5; b_sign3 = 4'd5;
@(posedge clk_i);
a_mant0 = 8'd246; a_mant1 = 8'd236; a_mant2 = 8'd197; a_mant3 = 8'd4;
b_mant0 = 8'd200; b_mant1 = 8'd15; b_mant2 = 8'd208; b_mant3 = 8'd16;
a_exp0 = 10'd409; a_exp1 = 10'd357; a_exp2 = 10'd454; a_exp3 = 10'd836;
b_exp0 = 10'd379; b_exp1 = 10'd220; b_exp2 = 10'd4; b_exp3 = 10'd747;
a_sign0 = 4'd12; a_sign1 = 4'd8; a_sign2 = 4'd7; a_sign3 = 4'd11;
b_sign0 = 4'd0; b_sign1 = 4'd16; b_sign2 = 4'd5; b_sign3 = 4'd3;
@(posedge clk_i);
a_mant0 = 8'd42; a_mant1 = 8'd161; a_mant2 = 8'd50; a_mant3 = 8'd164;
b_mant0 = 8'd74; b_mant1 = 8'd192; b_mant2 = 8'd251; b_mant3 = 8'd13;
a_exp0 = 10'd44; a_exp1 = 10'd745; a_exp2 = 10'd771; a_exp3 = 10'd356;
b_exp0 = 10'd1011; b_exp1 = 10'd119; b_exp2 = 10'd583; b_exp3 = 10'd208;
a_sign0 = 4'd13; a_sign1 = 4'd13; a_sign2 = 4'd15; a_sign3 = 4'd8;
b_sign0 = 4'd4; b_sign1 = 4'd1; b_sign2 = 4'd8; b_sign3 = 4'd8;
@(posedge clk_i);
a_mant0 = 8'd104; a_mant1 = 8'd29; a_mant2 = 8'd221; a_mant3 = 8'd220;
b_mant0 = 8'd53; b_mant1 = 8'd63; b_mant2 = 8'd12; b_mant3 = 8'd91;
a_exp0 = 10'd356; a_exp1 = 10'd1001; a_exp2 = 10'd768; a_exp3 = 10'd341;
b_exp0 = 10'd457; b_exp1 = 10'd223; b_exp2 = 10'd329; b_exp3 = 10'd538;
a_sign0 = 4'd16; a_sign1 = 4'd4; a_sign2 = 4'd14; a_sign3 = 4'd8;
b_sign0 = 4'd3; b_sign1 = 4'd0; b_sign2 = 4'd10; b_sign3 = 4'd10;
@(posedge clk_i);
a_mant0 = 8'd123; a_mant1 = 8'd167; a_mant2 = 8'd110; a_mant3 = 8'd33;
b_mant0 = 8'd211; b_mant1 = 8'd120; b_mant2 = 8'd111; b_mant3 = 8'd85;
a_exp0 = 10'd988; a_exp1 = 10'd530; a_exp2 = 10'd428; a_exp3 = 10'd393;
b_exp0 = 10'd1001; b_exp1 = 10'd494; b_exp2 = 10'd554; b_exp3 = 10'd807;
a_sign0 = 4'd1; a_sign1 = 4'd9; a_sign2 = 4'd11; a_sign3 = 4'd13;
b_sign0 = 4'd1; b_sign1 = 4'd1; b_sign2 = 4'd8; b_sign3 = 4'd15;
@(posedge clk_i);
a_mant0 = 8'd226; a_mant1 = 8'd32; a_mant2 = 8'd74; a_mant3 = 8'd222;
b_mant0 = 8'd15; b_mant1 = 8'd116; b_mant2 = 8'd49; b_mant3 = 8'd94;
a_exp0 = 10'd110; a_exp1 = 10'd177; a_exp2 = 10'd527; a_exp3 = 10'd421;
b_exp0 = 10'd813; b_exp1 = 10'd996; b_exp2 = 10'd1009; b_exp3 = 10'd813;
a_sign0 = 4'd2; a_sign1 = 4'd8; a_sign2 = 4'd5; a_sign3 = 4'd15;
b_sign0 = 4'd16; b_sign1 = 4'd11; b_sign2 = 4'd14; b_sign3 = 4'd7;
@(posedge clk_i);
a_mant0 = 8'd78; a_mant1 = 8'd160; a_mant2 = 8'd228; a_mant3 = 8'd83;
b_mant0 = 8'd198; b_mant1 = 8'd23; b_mant2 = 8'd101; b_mant3 = 8'd33;
a_exp0 = 10'd231; a_exp1 = 10'd379; a_exp2 = 10'd887; a_exp3 = 10'd802;
b_exp0 = 10'd810; b_exp1 = 10'd796; b_exp2 = 10'd1006; b_exp3 = 10'd400;
a_sign0 = 4'd16; a_sign1 = 4'd5; a_sign2 = 4'd2; a_sign3 = 4'd0;
b_sign0 = 4'd2; b_sign1 = 4'd2; b_sign2 = 4'd4; b_sign3 = 4'd10;
@(posedge clk_i);
a_mant0 = 8'd230; a_mant1 = 8'd173; a_mant2 = 8'd82; a_mant3 = 8'd146;
b_mant0 = 8'd64; b_mant1 = 8'd70; b_mant2 = 8'd225; b_mant3 = 8'd132;
a_exp0 = 10'd312; a_exp1 = 10'd576; a_exp2 = 10'd803; a_exp3 = 10'd850;
b_exp0 = 10'd618; b_exp1 = 10'd590; b_exp2 = 10'd393; b_exp3 = 10'd3;
a_sign0 = 4'd5; a_sign1 = 4'd4; a_sign2 = 4'd16; a_sign3 = 4'd8;
b_sign0 = 4'd6; b_sign1 = 4'd11; b_sign2 = 4'd0; b_sign3 = 4'd8;
@(posedge clk_i);
shared_exps0 = 8'd148;
shared_exps1 = 8'd114;
a_mant0 = 8'd10; a_mant1 = 8'd102; a_mant2 = 8'd159; a_mant3 = 8'd106;
b_mant0 = 8'd58; b_mant1 = 8'd71; b_mant2 = 8'd149; b_mant3 = 8'd122;
a_exp0 = 10'd524; a_exp1 = 10'd485; a_exp2 = 10'd684; a_exp3 = 10'd948;
b_exp0 = 10'd560; b_exp1 = 10'd84; b_exp2 = 10'd974; b_exp3 = 10'd856;
a_sign0 = 4'd0; a_sign1 = 4'd14; a_sign2 = 4'd15; a_sign3 = 4'd3;
b_sign0 = 4'd1; b_sign1 = 4'd13; b_sign2 = 4'd13; b_sign3 = 4'd13;
@(posedge clk_i);
a_mant0 = 8'd24; a_mant1 = 8'd225; a_mant2 = 8'd202; a_mant3 = 8'd90;
b_mant0 = 8'd234; b_mant1 = 8'd125; b_mant2 = 8'd183; b_mant3 = 8'd46;
a_exp0 = 10'd308; a_exp1 = 10'd208; a_exp2 = 10'd254; a_exp3 = 10'd111;
b_exp0 = 10'd65; b_exp1 = 10'd40; b_exp2 = 10'd73; b_exp3 = 10'd621;
a_sign0 = 4'd9; a_sign1 = 4'd7; a_sign2 = 4'd10; a_sign3 = 4'd8;
b_sign0 = 4'd14; b_sign1 = 4'd15; b_sign2 = 4'd0; b_sign3 = 4'd8;
@(posedge clk_i);
a_mant0 = 8'd253; a_mant1 = 8'd76; a_mant2 = 8'd89; a_mant3 = 8'd105;
b_mant0 = 8'd180; b_mant1 = 8'd0; b_mant2 = 8'd251; b_mant3 = 8'd94;
a_exp0 = 10'd979; a_exp1 = 10'd922; a_exp2 = 10'd525; a_exp3 = 10'd819;
b_exp0 = 10'd656; b_exp1 = 10'd116; b_exp2 = 10'd346; b_exp3 = 10'd756;
a_sign0 = 4'd9; a_sign1 = 4'd12; a_sign2 = 4'd14; a_sign3 = 4'd3;
b_sign0 = 4'd10; b_sign1 = 4'd2; b_sign2 = 4'd13; b_sign3 = 4'd7;
@(posedge clk_i);
a_mant0 = 8'd87; a_mant1 = 8'd172; a_mant2 = 8'd169; a_mant3 = 8'd48;
b_mant0 = 8'd188; b_mant1 = 8'd72; b_mant2 = 8'd43; b_mant3 = 8'd205;
a_exp0 = 10'd430; a_exp1 = 10'd695; a_exp2 = 10'd605; a_exp3 = 10'd840;
b_exp0 = 10'd150; b_exp1 = 10'd546; b_exp2 = 10'd472; b_exp3 = 10'd362;
a_sign0 = 4'd12; a_sign1 = 4'd9; a_sign2 = 4'd1; a_sign3 = 4'd14;
b_sign0 = 4'd4; b_sign1 = 4'd12; b_sign2 = 4'd3; b_sign3 = 4'd7;
@(posedge clk_i);
a_mant0 = 8'd149; a_mant1 = 8'd1; a_mant2 = 8'd97; a_mant3 = 8'd66;
b_mant0 = 8'd130; b_mant1 = 8'd74; b_mant2 = 8'd240; b_mant3 = 8'd239;
a_exp0 = 10'd792; a_exp1 = 10'd502; a_exp2 = 10'd596; a_exp3 = 10'd350;
b_exp0 = 10'd846; b_exp1 = 10'd294; b_exp2 = 10'd195; b_exp3 = 10'd1;
a_sign0 = 4'd11; a_sign1 = 4'd3; a_sign2 = 4'd4; a_sign3 = 4'd8;
b_sign0 = 4'd4; b_sign1 = 4'd7; b_sign2 = 4'd10; b_sign3 = 4'd2;
@(posedge clk_i);
a_mant0 = 8'd212; a_mant1 = 8'd176; a_mant2 = 8'd208; a_mant3 = 8'd153;
b_mant0 = 8'd3; b_mant1 = 8'd209; b_mant2 = 8'd93; b_mant3 = 8'd106;
a_exp0 = 10'd70; a_exp1 = 10'd134; a_exp2 = 10'd432; a_exp3 = 10'd544;
b_exp0 = 10'd450; b_exp1 = 10'd503; b_exp2 = 10'd699; b_exp3 = 10'd290;
a_sign0 = 4'd13; a_sign1 = 4'd14; a_sign2 = 4'd7; a_sign3 = 4'd16;
b_sign0 = 4'd8; b_sign1 = 4'd16; b_sign2 = 4'd0; b_sign3 = 4'd3;
@(posedge clk_i);
a_mant0 = 8'd146; a_mant1 = 8'd219; a_mant2 = 8'd195; a_mant3 = 8'd115;
b_mant0 = 8'd236; b_mant1 = 8'd142; b_mant2 = 8'd233; b_mant3 = 8'd26;
a_exp0 = 10'd131; a_exp1 = 10'd905; a_exp2 = 10'd773; a_exp3 = 10'd415;
b_exp0 = 10'd244; b_exp1 = 10'd326; b_exp2 = 10'd704; b_exp3 = 10'd461;
a_sign0 = 4'd0; a_sign1 = 4'd1; a_sign2 = 4'd11; a_sign3 = 4'd13;
b_sign0 = 4'd5; b_sign1 = 4'd16; b_sign2 = 4'd3; b_sign3 = 4'd16;
@(posedge clk_i);
a_mant0 = 8'd135; a_mant1 = 8'd142; a_mant2 = 8'd64; a_mant3 = 8'd219;
b_mant0 = 8'd132; b_mant1 = 8'd164; b_mant2 = 8'd59; b_mant3 = 8'd107;
a_exp0 = 10'd648; a_exp1 = 10'd248; a_exp2 = 10'd355; a_exp3 = 10'd999;
b_exp0 = 10'd91; b_exp1 = 10'd57; b_exp2 = 10'd949; b_exp3 = 10'd317;
a_sign0 = 4'd15; a_sign1 = 4'd14; a_sign2 = 4'd6; a_sign3 = 4'd5;
b_sign0 = 4'd4; b_sign1 = 4'd9; b_sign2 = 4'd6; b_sign3 = 4'd1;
@(posedge clk_i);
shared_exps0 = 8'd136;
shared_exps1 = 8'd144;
rstn = 0;
@(posedge clk_i);
rstn = 1;
a_mant0 = 8'd90; a_mant1 = 8'd159; a_mant2 = 8'd122; a_mant3 = 8'd190;
b_mant0 = 8'd113; b_mant1 = 8'd131; b_mant2 = 8'd143; b_mant3 = 8'd19;
a_exp0 = 10'd297; a_exp1 = 10'd72; a_exp2 = 10'd449; a_exp3 = 10'd679;
b_exp0 = 10'd1007; b_exp1 = 10'd338; b_exp2 = 10'd843; b_exp3 = 10'd732;
a_sign0 = 4'd3; a_sign1 = 4'd6; a_sign2 = 4'd11; a_sign3 = 4'd14;
b_sign0 = 4'd10; b_sign1 = 4'd13; b_sign2 = 4'd5; b_sign3 = 4'd9;
@(posedge clk_i);
a_mant0 = 8'd84; a_mant1 = 8'd41; a_mant2 = 8'd140; a_mant3 = 8'd186;
b_mant0 = 8'd107; b_mant1 = 8'd126; b_mant2 = 8'd191; b_mant3 = 8'd248;
a_exp0 = 10'd387; a_exp1 = 10'd390; a_exp2 = 10'd506; a_exp3 = 10'd373;
b_exp0 = 10'd654; b_exp1 = 10'd49; b_exp2 = 10'd527; b_exp3 = 10'd60;
a_sign0 = 4'd14; a_sign1 = 4'd0; a_sign2 = 4'd6; a_sign3 = 4'd2;
b_sign0 = 4'd2; b_sign1 = 4'd5; b_sign2 = 4'd10; b_sign3 = 4'd2;
@(posedge clk_i);
a_mant0 = 8'd60; a_mant1 = 8'd162; a_mant2 = 8'd96; a_mant3 = 8'd111;
b_mant0 = 8'd172; b_mant1 = 8'd173; b_mant2 = 8'd140; b_mant3 = 8'd174;
a_exp0 = 10'd763; a_exp1 = 10'd590; a_exp2 = 10'd497; a_exp3 = 10'd453;
b_exp0 = 10'd583; b_exp1 = 10'd597; b_exp2 = 10'd68; b_exp3 = 10'd201;
a_sign0 = 4'd9; a_sign1 = 4'd8; a_sign2 = 4'd5; a_sign3 = 4'd12;
b_sign0 = 4'd14; b_sign1 = 4'd11; b_sign2 = 4'd5; b_sign3 = 4'd1;
@(posedge clk_i);
a_mant0 = 8'd166; a_mant1 = 8'd21; a_mant2 = 8'd183; a_mant3 = 8'd189;
b_mant0 = 8'd78; b_mant1 = 8'd17; b_mant2 = 8'd84; b_mant3 = 8'd150;
a_exp0 = 10'd997; a_exp1 = 10'd835; a_exp2 = 10'd724; a_exp3 = 10'd166;
b_exp0 = 10'd650; b_exp1 = 10'd100; b_exp2 = 10'd311; b_exp3 = 10'd332;
a_sign0 = 4'd14; a_sign1 = 4'd2; a_sign2 = 4'd16; a_sign3 = 4'd0;
b_sign0 = 4'd12; b_sign1 = 4'd15; b_sign2 = 4'd9; b_sign3 = 4'd10;
@(posedge clk_i);
a_mant0 = 8'd84; a_mant1 = 8'd38; a_mant2 = 8'd179; a_mant3 = 8'd226;
b_mant0 = 8'd108; b_mant1 = 8'd185; b_mant2 = 8'd244; b_mant3 = 8'd162;
a_exp0 = 10'd769; a_exp1 = 10'd87; a_exp2 = 10'd769; a_exp3 = 10'd413;
b_exp0 = 10'd352; b_exp1 = 10'd546; b_exp2 = 10'd417; b_exp3 = 10'd439;
a_sign0 = 4'd2; a_sign1 = 4'd14; a_sign2 = 4'd5; a_sign3 = 4'd7;
b_sign0 = 4'd13; b_sign1 = 4'd2; b_sign2 = 4'd6; b_sign3 = 4'd16;
@(posedge clk_i);
a_mant0 = 8'd63; a_mant1 = 8'd131; a_mant2 = 8'd191; a_mant3 = 8'd160;
b_mant0 = 8'd160; b_mant1 = 8'd204; b_mant2 = 8'd221; b_mant3 = 8'd71;
a_exp0 = 10'd112; a_exp1 = 10'd854; a_exp2 = 10'd934; a_exp3 = 10'd532;
b_exp0 = 10'd288; b_exp1 = 10'd21; b_exp2 = 10'd903; b_exp3 = 10'd106;
a_sign0 = 4'd12; a_sign1 = 4'd7; a_sign2 = 4'd16; a_sign3 = 4'd10;
b_sign0 = 4'd2; b_sign1 = 4'd12; b_sign2 = 4'd0; b_sign3 = 4'd3;
@(posedge clk_i);
a_mant0 = 8'd42; a_mant1 = 8'd66; a_mant2 = 8'd145; a_mant3 = 8'd227;
b_mant0 = 8'd240; b_mant1 = 8'd29; b_mant2 = 8'd227; b_mant3 = 8'd225;
a_exp0 = 10'd454; a_exp1 = 10'd725; a_exp2 = 10'd398; a_exp3 = 10'd302;
b_exp0 = 10'd706; b_exp1 = 10'd265; b_exp2 = 10'd1021; b_exp3 = 10'd836;
a_sign0 = 4'd8; a_sign1 = 4'd16; a_sign2 = 4'd14; a_sign3 = 4'd13;
b_sign0 = 4'd5; b_sign1 = 4'd13; b_sign2 = 4'd3; b_sign3 = 4'd6;
@(posedge clk_i);
shared_exps0 = 8'd140;
shared_exps1 = 8'd99;
a_mant0 = 8'd58; a_mant1 = 8'd146; a_mant2 = 8'd151; a_mant3 = 8'd249;
b_mant0 = 8'd102; b_mant1 = 8'd128; b_mant2 = 8'd200; b_mant3 = 8'd255;
a_exp0 = 10'd412; a_exp1 = 10'd301; a_exp2 = 10'd134; a_exp3 = 10'd402;
b_exp0 = 10'd1019; b_exp1 = 10'd292; b_exp2 = 10'd586; b_exp3 = 10'd508;
a_sign0 = 4'd11; a_sign1 = 4'd1; a_sign2 = 4'd10; a_sign3 = 4'd0;
b_sign0 = 4'd8; b_sign1 = 4'd10; b_sign2 = 4'd2; b_sign3 = 4'd5;
@(posedge clk_i);
a_mant0 = 8'd170; a_mant1 = 8'd52; a_mant2 = 8'd231; a_mant3 = 8'd69;
b_mant0 = 8'd48; b_mant1 = 8'd137; b_mant2 = 8'd65; b_mant3 = 8'd149;
a_exp0 = 10'd771; a_exp1 = 10'd42; a_exp2 = 10'd386; a_exp3 = 10'd457;
b_exp0 = 10'd413; b_exp1 = 10'd393; b_exp2 = 10'd933; b_exp3 = 10'd809;
a_sign0 = 4'd12; a_sign1 = 4'd0; a_sign2 = 4'd6; a_sign3 = 4'd2;
b_sign0 = 4'd10; b_sign1 = 4'd1; b_sign2 = 4'd2; b_sign3 = 4'd11;
@(posedge clk_i);
a_mant0 = 8'd211; a_mant1 = 8'd146; a_mant2 = 8'd220; a_mant3 = 8'd63;
b_mant0 = 8'd32; b_mant1 = 8'd67; b_mant2 = 8'd94; b_mant3 = 8'd31;
a_exp0 = 10'd922; a_exp1 = 10'd110; a_exp2 = 10'd307; a_exp3 = 10'd477;
b_exp0 = 10'd877; b_exp1 = 10'd10; b_exp2 = 10'd193; b_exp3 = 10'd234;
a_sign0 = 4'd16; a_sign1 = 4'd7; a_sign2 = 4'd12; a_sign3 = 4'd0;
b_sign0 = 4'd5; b_sign1 = 4'd16; b_sign2 = 4'd15; b_sign3 = 4'd10;
@(posedge clk_i);
a_mant0 = 8'd56; a_mant1 = 8'd104; a_mant2 = 8'd89; a_mant3 = 8'd174;
b_mant0 = 8'd19; b_mant1 = 8'd99; b_mant2 = 8'd24; b_mant3 = 8'd98;
a_exp0 = 10'd981; a_exp1 = 10'd378; a_exp2 = 10'd897; a_exp3 = 10'd927;
b_exp0 = 10'd262; b_exp1 = 10'd585; b_exp2 = 10'd528; b_exp3 = 10'd734;
a_sign0 = 4'd9; a_sign1 = 4'd16; a_sign2 = 4'd6; a_sign3 = 4'd9;
b_sign0 = 4'd16; b_sign1 = 4'd14; b_sign2 = 4'd12; b_sign3 = 4'd10;
@(posedge clk_i);
a_mant0 = 8'd184; a_mant1 = 8'd201; a_mant2 = 8'd62; a_mant3 = 8'd82;
b_mant0 = 8'd242; b_mant1 = 8'd99; b_mant2 = 8'd151; b_mant3 = 8'd214;
a_exp0 = 10'd835; a_exp1 = 10'd761; a_exp2 = 10'd198; a_exp3 = 10'd793;
b_exp0 = 10'd855; b_exp1 = 10'd985; b_exp2 = 10'd998; b_exp3 = 10'd633;
a_sign0 = 4'd3; a_sign1 = 4'd2; a_sign2 = 4'd5; a_sign3 = 4'd1;
b_sign0 = 4'd8; b_sign1 = 4'd3; b_sign2 = 4'd11; b_sign3 = 4'd15;
@(posedge clk_i);
a_mant0 = 8'd79; a_mant1 = 8'd190; a_mant2 = 8'd28; a_mant3 = 8'd39;
b_mant0 = 8'd11; b_mant1 = 8'd104; b_mant2 = 8'd217; b_mant3 = 8'd15;
a_exp0 = 10'd165; a_exp1 = 10'd83; a_exp2 = 10'd34; a_exp3 = 10'd653;
b_exp0 = 10'd469; b_exp1 = 10'd109; b_exp2 = 10'd476; b_exp3 = 10'd829;
a_sign0 = 4'd6; a_sign1 = 4'd16; a_sign2 = 4'd12; a_sign3 = 4'd0;
b_sign0 = 4'd4; b_sign1 = 4'd4; b_sign2 = 4'd9; b_sign3 = 4'd15;
@(posedge clk_i);
a_mant0 = 8'd175; a_mant1 = 8'd59; a_mant2 = 8'd54; a_mant3 = 8'd148;
b_mant0 = 8'd17; b_mant1 = 8'd184; b_mant2 = 8'd76; b_mant3 = 8'd195;
a_exp0 = 10'd126; a_exp1 = 10'd377; a_exp2 = 10'd476; a_exp3 = 10'd630;
b_exp0 = 10'd530; b_exp1 = 10'd538; b_exp2 = 10'd55; b_exp3 = 10'd508;
a_sign0 = 4'd4; a_sign1 = 4'd10; a_sign2 = 4'd9; a_sign3 = 4'd5;
b_sign0 = 4'd4; b_sign1 = 4'd4; b_sign2 = 4'd7; b_sign3 = 4'd3;
@(posedge clk_i);
a_mant0 = 8'd16; a_mant1 = 8'd84; a_mant2 = 8'd124; a_mant3 = 8'd151;
b_mant0 = 8'd83; b_mant1 = 8'd3; b_mant2 = 8'd17; b_mant3 = 8'd191;
a_exp0 = 10'd887; a_exp1 = 10'd695; a_exp2 = 10'd582; a_exp3 = 10'd10;
b_exp0 = 10'd441; b_exp1 = 10'd699; b_exp2 = 10'd32; b_exp3 = 10'd12;
a_sign0 = 4'd16; a_sign1 = 4'd12; a_sign2 = 4'd8; a_sign3 = 4'd11;
b_sign0 = 4'd1; b_sign1 = 4'd5; b_sign2 = 4'd12; b_sign3 = 4'd8;
@(posedge clk_i);
shared_exps0 = 8'd143;
shared_exps1 = 8'd130;
a_mant0 = 8'd213; a_mant1 = 8'd10; a_mant2 = 8'd155; a_mant3 = 8'd156;
b_mant0 = 8'd82; b_mant1 = 8'd250; b_mant2 = 8'd197; b_mant3 = 8'd44;
a_exp0 = 10'd317; a_exp1 = 10'd807; a_exp2 = 10'd489; a_exp3 = 10'd556;
b_exp0 = 10'd908; b_exp1 = 10'd552; b_exp2 = 10'd476; b_exp3 = 10'd916;
a_sign0 = 4'd2; a_sign1 = 4'd2; a_sign2 = 4'd13; a_sign3 = 4'd14;
b_sign0 = 4'd2; b_sign1 = 4'd16; b_sign2 = 4'd2; b_sign3 = 4'd9;
@(posedge clk_i);
a_mant0 = 8'd164; a_mant1 = 8'd10; a_mant2 = 8'd82; a_mant3 = 8'd233;
b_mant0 = 8'd60; b_mant1 = 8'd240; b_mant2 = 8'd132; b_mant3 = 8'd45;
a_exp0 = 10'd607; a_exp1 = 10'd285; a_exp2 = 10'd916; a_exp3 = 10'd262;
b_exp0 = 10'd130; b_exp1 = 10'd578; b_exp2 = 10'd92; b_exp3 = 10'd336;
a_sign0 = 4'd7; a_sign1 = 4'd14; a_sign2 = 4'd3; a_sign3 = 4'd10;
b_sign0 = 4'd11; b_sign1 = 4'd13; b_sign2 = 4'd9; b_sign3 = 4'd2;
@(posedge clk_i);
a_mant0 = 8'd47; a_mant1 = 8'd9; a_mant2 = 8'd153; a_mant3 = 8'd103;
b_mant0 = 8'd202; b_mant1 = 8'd27; b_mant2 = 8'd60; b_mant3 = 8'd125;
a_exp0 = 10'd882; a_exp1 = 10'd508; a_exp2 = 10'd869; a_exp3 = 10'd44;
b_exp0 = 10'd911; b_exp1 = 10'd554; b_exp2 = 10'd35; b_exp3 = 10'd120;
a_sign0 = 4'd2; a_sign1 = 4'd10; a_sign2 = 4'd8; a_sign3 = 4'd10;
b_sign0 = 4'd15; b_sign1 = 4'd14; b_sign2 = 4'd13; b_sign3 = 4'd8;
@(posedge clk_i);
a_mant0 = 8'd85; a_mant1 = 8'd209; a_mant2 = 8'd151; a_mant3 = 8'd106;
b_mant0 = 8'd39; b_mant1 = 8'd41; b_mant2 = 8'd91; b_mant3 = 8'd192;
a_exp0 = 10'd977; a_exp1 = 10'd958; a_exp2 = 10'd686; a_exp3 = 10'd221;
b_exp0 = 10'd529; b_exp1 = 10'd409; b_exp2 = 10'd649; b_exp3 = 10'd148;
a_sign0 = 4'd6; a_sign1 = 4'd2; a_sign2 = 4'd1; a_sign3 = 4'd13;
b_sign0 = 4'd8; b_sign1 = 4'd0; b_sign2 = 4'd1; b_sign3 = 4'd1;
@(posedge clk_i);
a_mant0 = 8'd151; a_mant1 = 8'd118; a_mant2 = 8'd6; a_mant3 = 8'd210;
b_mant0 = 8'd162; b_mant1 = 8'd131; b_mant2 = 8'd29; b_mant3 = 8'd0;
a_exp0 = 10'd745; a_exp1 = 10'd890; a_exp2 = 10'd129; a_exp3 = 10'd478;
b_exp0 = 10'd375; b_exp1 = 10'd565; b_exp2 = 10'd150; b_exp3 = 10'd466;
a_sign0 = 4'd6; a_sign1 = 4'd2; a_sign2 = 4'd0; a_sign3 = 4'd8;
b_sign0 = 4'd12; b_sign1 = 4'd11; b_sign2 = 4'd10; b_sign3 = 4'd13;
@(posedge clk_i);
a_mant0 = 8'd96; a_mant1 = 8'd111; a_mant2 = 8'd171; a_mant3 = 8'd14;
b_mant0 = 8'd109; b_mant1 = 8'd182; b_mant2 = 8'd141; b_mant3 = 8'd4;
a_exp0 = 10'd824; a_exp1 = 10'd457; a_exp2 = 10'd343; a_exp3 = 10'd636;
b_exp0 = 10'd202; b_exp1 = 10'd226; b_exp2 = 10'd216; b_exp3 = 10'd640;
a_sign0 = 4'd13; a_sign1 = 4'd12; a_sign2 = 4'd15; a_sign3 = 4'd16;
b_sign0 = 4'd15; b_sign1 = 4'd8; b_sign2 = 4'd4; b_sign3 = 4'd11;
@(posedge clk_i);
a_mant0 = 8'd160; a_mant1 = 8'd247; a_mant2 = 8'd8; a_mant3 = 8'd123;
b_mant0 = 8'd231; b_mant1 = 8'd115; b_mant2 = 8'd77; b_mant3 = 8'd34;
a_exp0 = 10'd591; a_exp1 = 10'd137; a_exp2 = 10'd1005; a_exp3 = 10'd797;
b_exp0 = 10'd250; b_exp1 = 10'd343; b_exp2 = 10'd650; b_exp3 = 10'd721;
a_sign0 = 4'd7; a_sign1 = 4'd1; a_sign2 = 4'd12; a_sign3 = 4'd3;
b_sign0 = 4'd8; b_sign1 = 4'd4; b_sign2 = 4'd10; b_sign3 = 4'd13;
@(posedge clk_i);
a_mant0 = 8'd36; a_mant1 = 8'd194; a_mant2 = 8'd79; a_mant3 = 8'd90;
b_mant0 = 8'd76; b_mant1 = 8'd123; b_mant2 = 8'd30; b_mant3 = 8'd158;
a_exp0 = 10'd628; a_exp1 = 10'd27; a_exp2 = 10'd624; a_exp3 = 10'd254;
b_exp0 = 10'd550; b_exp1 = 10'd416; b_exp2 = 10'd879; b_exp3 = 10'd4;
a_sign0 = 4'd12; a_sign1 = 4'd5; a_sign2 = 4'd12; a_sign3 = 4'd14;
b_sign0 = 4'd7; b_sign1 = 4'd2; b_sign2 = 4'd12; b_sign3 = 4'd9;
@(posedge clk_i);
shared_exps0 = 8'd139;
shared_exps1 = 8'd132;
a_mant0 = 8'd197; a_mant1 = 8'd149; a_mant2 = 8'd114; a_mant3 = 8'd29;
b_mant0 = 8'd133; b_mant1 = 8'd45; b_mant2 = 8'd157; b_mant3 = 8'd191;
a_exp0 = 10'd559; a_exp1 = 10'd654; a_exp2 = 10'd1015; a_exp3 = 10'd556;
b_exp0 = 10'd399; b_exp1 = 10'd662; b_exp2 = 10'd230; b_exp3 = 10'd776;
a_sign0 = 4'd1; a_sign1 = 4'd0; a_sign2 = 4'd14; a_sign3 = 4'd8;
b_sign0 = 4'd7; b_sign1 = 4'd4; b_sign2 = 4'd10; b_sign3 = 4'd1;
@(posedge clk_i);
a_mant0 = 8'd108; a_mant1 = 8'd12; a_mant2 = 8'd28; a_mant3 = 8'd22;
b_mant0 = 8'd212; b_mant1 = 8'd191; b_mant2 = 8'd119; b_mant3 = 8'd246;
a_exp0 = 10'd821; a_exp1 = 10'd635; a_exp2 = 10'd185; a_exp3 = 10'd263;
b_exp0 = 10'd783; b_exp1 = 10'd273; b_exp2 = 10'd352; b_exp3 = 10'd865;
a_sign0 = 4'd10; a_sign1 = 4'd12; a_sign2 = 4'd8; a_sign3 = 4'd16;
b_sign0 = 4'd3; b_sign1 = 4'd1; b_sign2 = 4'd5; b_sign3 = 4'd9;
@(posedge clk_i);
a_mant0 = 8'd97; a_mant1 = 8'd163; a_mant2 = 8'd216; a_mant3 = 8'd79;
b_mant0 = 8'd214; b_mant1 = 8'd164; b_mant2 = 8'd119; b_mant3 = 8'd9;
a_exp0 = 10'd732; a_exp1 = 10'd938; a_exp2 = 10'd193; a_exp3 = 10'd155;
b_exp0 = 10'd611; b_exp1 = 10'd43; b_exp2 = 10'd66; b_exp3 = 10'd1010;
a_sign0 = 4'd16; a_sign1 = 4'd13; a_sign2 = 4'd16; a_sign3 = 4'd10;
b_sign0 = 4'd6; b_sign1 = 4'd7; b_sign2 = 4'd9; b_sign3 = 4'd4;
@(posedge clk_i);
a_mant0 = 8'd178; a_mant1 = 8'd23; a_mant2 = 8'd198; a_mant3 = 8'd187;
b_mant0 = 8'd149; b_mant1 = 8'd82; b_mant2 = 8'd7; b_mant3 = 8'd3;
a_exp0 = 10'd115; a_exp1 = 10'd569; a_exp2 = 10'd635; a_exp3 = 10'd686;
b_exp0 = 10'd134; b_exp1 = 10'd791; b_exp2 = 10'd359; b_exp3 = 10'd556;
a_sign0 = 4'd6; a_sign1 = 4'd8; a_sign2 = 4'd5; a_sign3 = 4'd8;
b_sign0 = 4'd12; b_sign1 = 4'd5; b_sign2 = 4'd7; b_sign3 = 4'd3;
@(posedge clk_i);
a_mant0 = 8'd238; a_mant1 = 8'd252; a_mant2 = 8'd25; a_mant3 = 8'd132;
b_mant0 = 8'd208; b_mant1 = 8'd77; b_mant2 = 8'd120; b_mant3 = 8'd66;
a_exp0 = 10'd378; a_exp1 = 10'd440; a_exp2 = 10'd924; a_exp3 = 10'd307;
b_exp0 = 10'd748; b_exp1 = 10'd906; b_exp2 = 10'd206; b_exp3 = 10'd662;
a_sign0 = 4'd13; a_sign1 = 4'd6; a_sign2 = 4'd5; a_sign3 = 4'd8;
b_sign0 = 4'd1; b_sign1 = 4'd0; b_sign2 = 4'd9; b_sign3 = 4'd11;
@(posedge clk_i);
a_mant0 = 8'd222; a_mant1 = 8'd103; a_mant2 = 8'd166; a_mant3 = 8'd42;
b_mant0 = 8'd27; b_mant1 = 8'd113; b_mant2 = 8'd161; b_mant3 = 8'd48;
a_exp0 = 10'd903; a_exp1 = 10'd1004; a_exp2 = 10'd129; a_exp3 = 10'd415;
b_exp0 = 10'd685; b_exp1 = 10'd172; b_exp2 = 10'd832; b_exp3 = 10'd987;
a_sign0 = 4'd11; a_sign1 = 4'd13; a_sign2 = 4'd4; a_sign3 = 4'd7;
b_sign0 = 4'd1; b_sign1 = 4'd12; b_sign2 = 4'd1; b_sign3 = 4'd4;
@(posedge clk_i);
a_mant0 = 8'd134; a_mant1 = 8'd82; a_mant2 = 8'd98; a_mant3 = 8'd13;
b_mant0 = 8'd8; b_mant1 = 8'd229; b_mant2 = 8'd90; b_mant3 = 8'd155;
a_exp0 = 10'd197; a_exp1 = 10'd619; a_exp2 = 10'd386; a_exp3 = 10'd410;
b_exp0 = 10'd4; b_exp1 = 10'd815; b_exp2 = 10'd678; b_exp3 = 10'd81;
a_sign0 = 4'd16; a_sign1 = 4'd16; a_sign2 = 4'd15; a_sign3 = 4'd13;
b_sign0 = 4'd12; b_sign1 = 4'd12; b_sign2 = 4'd7; b_sign3 = 4'd7;
@(posedge clk_i);
a_mant0 = 8'd101; a_mant1 = 8'd69; a_mant2 = 8'd215; a_mant3 = 8'd149;
b_mant0 = 8'd170; b_mant1 = 8'd115; b_mant2 = 8'd116; b_mant3 = 8'd53;
a_exp0 = 10'd826; a_exp1 = 10'd684; a_exp2 = 10'd176; a_exp3 = 10'd849;
b_exp0 = 10'd589; b_exp1 = 10'd107; b_exp2 = 10'd805; b_exp3 = 10'd514;
a_sign0 = 4'd9; a_sign1 = 4'd2; a_sign2 = 4'd11; a_sign3 = 4'd9;
b_sign0 = 4'd14; b_sign1 = 4'd0; b_sign2 = 4'd6; b_sign3 = 4'd7;
@(posedge clk_i);
shared_exps0 = 8'd99;
shared_exps1 = 8'd129;
rstn = 0;
@(posedge clk_i);
rstn = 1;
a_mant0 = 8'd188; a_mant1 = 8'd82; a_mant2 = 8'd22; a_mant3 = 8'd8;
b_mant0 = 8'd124; b_mant1 = 8'd76; b_mant2 = 8'd117; b_mant3 = 8'd224;
a_exp0 = 10'd895; a_exp1 = 10'd272; a_exp2 = 10'd90; a_exp3 = 10'd603;
b_exp0 = 10'd721; b_exp1 = 10'd606; b_exp2 = 10'd420; b_exp3 = 10'd555;
a_sign0 = 4'd0; a_sign1 = 4'd5; a_sign2 = 4'd10; a_sign3 = 4'd0;
b_sign0 = 4'd14; b_sign1 = 4'd6; b_sign2 = 4'd16; b_sign3 = 4'd9;
@(posedge clk_i);
a_mant0 = 8'd195; a_mant1 = 8'd161; a_mant2 = 8'd249; a_mant3 = 8'd195;
b_mant0 = 8'd203; b_mant1 = 8'd242; b_mant2 = 8'd56; b_mant3 = 8'd169;
a_exp0 = 10'd614; a_exp1 = 10'd396; a_exp2 = 10'd901; a_exp3 = 10'd836;
b_exp0 = 10'd476; b_exp1 = 10'd667; b_exp2 = 10'd175; b_exp3 = 10'd160;
a_sign0 = 4'd10; a_sign1 = 4'd4; a_sign2 = 4'd0; a_sign3 = 4'd10;
b_sign0 = 4'd12; b_sign1 = 4'd4; b_sign2 = 4'd11; b_sign3 = 4'd16;
@(posedge clk_i);
a_mant0 = 8'd50; a_mant1 = 8'd112; a_mant2 = 8'd245; a_mant3 = 8'd24;
b_mant0 = 8'd195; b_mant1 = 8'd127; b_mant2 = 8'd43; b_mant3 = 8'd106;
a_exp0 = 10'd795; a_exp1 = 10'd240; a_exp2 = 10'd578; a_exp3 = 10'd672;
b_exp0 = 10'd774; b_exp1 = 10'd30; b_exp2 = 10'd948; b_exp3 = 10'd28;
a_sign0 = 4'd12; a_sign1 = 4'd3; a_sign2 = 4'd0; a_sign3 = 4'd16;
b_sign0 = 4'd5; b_sign1 = 4'd13; b_sign2 = 4'd10; b_sign3 = 4'd16;
@(posedge clk_i);
a_mant0 = 8'd127; a_mant1 = 8'd40; a_mant2 = 8'd15; a_mant3 = 8'd238;
b_mant0 = 8'd186; b_mant1 = 8'd32; b_mant2 = 8'd99; b_mant3 = 8'd148;
a_exp0 = 10'd662; a_exp1 = 10'd915; a_exp2 = 10'd264; a_exp3 = 10'd316;
b_exp0 = 10'd659; b_exp1 = 10'd405; b_exp2 = 10'd989; b_exp3 = 10'd988;
a_sign0 = 4'd15; a_sign1 = 4'd8; a_sign2 = 4'd14; a_sign3 = 4'd0;
b_sign0 = 4'd12; b_sign1 = 4'd0; b_sign2 = 4'd8; b_sign3 = 4'd14;
@(posedge clk_i);
a_mant0 = 8'd255; a_mant1 = 8'd117; a_mant2 = 8'd103; a_mant3 = 8'd250;
b_mant0 = 8'd71; b_mant1 = 8'd150; b_mant2 = 8'd217; b_mant3 = 8'd156;
a_exp0 = 10'd266; a_exp1 = 10'd877; a_exp2 = 10'd601; a_exp3 = 10'd648;
b_exp0 = 10'd995; b_exp1 = 10'd437; b_exp2 = 10'd73; b_exp3 = 10'd445;
a_sign0 = 4'd2; a_sign1 = 4'd0; a_sign2 = 4'd5; a_sign3 = 4'd13;
b_sign0 = 4'd2; b_sign1 = 4'd1; b_sign2 = 4'd4; b_sign3 = 4'd11;
@(posedge clk_i);
a_mant0 = 8'd90; a_mant1 = 8'd229; a_mant2 = 8'd194; a_mant3 = 8'd54;
b_mant0 = 8'd169; b_mant1 = 8'd14; b_mant2 = 8'd157; b_mant3 = 8'd85;
a_exp0 = 10'd928; a_exp1 = 10'd523; a_exp2 = 10'd786; a_exp3 = 10'd622;
b_exp0 = 10'd767; b_exp1 = 10'd140; b_exp2 = 10'd481; b_exp3 = 10'd230;
a_sign0 = 4'd6; a_sign1 = 4'd13; a_sign2 = 4'd0; a_sign3 = 4'd10;
b_sign0 = 4'd3; b_sign1 = 4'd16; b_sign2 = 4'd14; b_sign3 = 4'd14;
@(posedge clk_i);
a_mant0 = 8'd220; a_mant1 = 8'd207; a_mant2 = 8'd29; a_mant3 = 8'd251;
b_mant0 = 8'd6; b_mant1 = 8'd71; b_mant2 = 8'd40; b_mant3 = 8'd191;
a_exp0 = 10'd894; a_exp1 = 10'd360; a_exp2 = 10'd162; a_exp3 = 10'd52;
b_exp0 = 10'd919; b_exp1 = 10'd583; b_exp2 = 10'd7; b_exp3 = 10'd417;
a_sign0 = 4'd1; a_sign1 = 4'd2; a_sign2 = 4'd14; a_sign3 = 4'd5;
b_sign0 = 4'd4; b_sign1 = 4'd6; b_sign2 = 4'd10; b_sign3 = 4'd8;
@(posedge clk_i);
shared_exps0 = 8'd138;
shared_exps1 = 8'd128;
a_mant0 = 8'd217; a_mant1 = 8'd97; a_mant2 = 8'd134; a_mant3 = 8'd41;
b_mant0 = 8'd46; b_mant1 = 8'd212; b_mant2 = 8'd59; b_mant3 = 8'd220;
a_exp0 = 10'd201; a_exp1 = 10'd342; a_exp2 = 10'd1015; a_exp3 = 10'd408;
b_exp0 = 10'd722; b_exp1 = 10'd100; b_exp2 = 10'd805; b_exp3 = 10'd793;
a_sign0 = 4'd11; a_sign1 = 4'd9; a_sign2 = 4'd6; a_sign3 = 4'd7;
b_sign0 = 4'd12; b_sign1 = 4'd6; b_sign2 = 4'd14; b_sign3 = 4'd4;
@(posedge clk_i);
a_mant0 = 8'd238; a_mant1 = 8'd87; a_mant2 = 8'd1; a_mant3 = 8'd200;
b_mant0 = 8'd243; b_mant1 = 8'd47; b_mant2 = 8'd76; b_mant3 = 8'd166;
a_exp0 = 10'd922; a_exp1 = 10'd604; a_exp2 = 10'd270; a_exp3 = 10'd522;
b_exp0 = 10'd350; b_exp1 = 10'd75; b_exp2 = 10'd524; b_exp3 = 10'd115;
a_sign0 = 4'd12; a_sign1 = 4'd5; a_sign2 = 4'd14; a_sign3 = 4'd4;
b_sign0 = 4'd13; b_sign1 = 4'd6; b_sign2 = 4'd6; b_sign3 = 4'd15;
@(posedge clk_i);
a_mant0 = 8'd70; a_mant1 = 8'd169; a_mant2 = 8'd154; a_mant3 = 8'd57;
b_mant0 = 8'd188; b_mant1 = 8'd179; b_mant2 = 8'd207; b_mant3 = 8'd211;
a_exp0 = 10'd568; a_exp1 = 10'd682; a_exp2 = 10'd347; a_exp3 = 10'd641;
b_exp0 = 10'd80; b_exp1 = 10'd285; b_exp2 = 10'd329; b_exp3 = 10'd508;
a_sign0 = 4'd1; a_sign1 = 4'd12; a_sign2 = 4'd15; a_sign3 = 4'd4;
b_sign0 = 4'd12; b_sign1 = 4'd0; b_sign2 = 4'd12; b_sign3 = 4'd14;
@(posedge clk_i);
a_mant0 = 8'd225; a_mant1 = 8'd142; a_mant2 = 8'd241; a_mant3 = 8'd194;
b_mant0 = 8'd70; b_mant1 = 8'd200; b_mant2 = 8'd37; b_mant3 = 8'd255;
a_exp0 = 10'd746; a_exp1 = 10'd375; a_exp2 = 10'd151; a_exp3 = 10'd479;
b_exp0 = 10'd462; b_exp1 = 10'd505; b_exp2 = 10'd274; b_exp3 = 10'd996;
a_sign0 = 4'd16; a_sign1 = 4'd1; a_sign2 = 4'd15; a_sign3 = 4'd5;
b_sign0 = 4'd11; b_sign1 = 4'd15; b_sign2 = 4'd13; b_sign3 = 4'd9;
@(posedge clk_i);
a_mant0 = 8'd97; a_mant1 = 8'd153; a_mant2 = 8'd55; a_mant3 = 8'd75;
b_mant0 = 8'd227; b_mant1 = 8'd35; b_mant2 = 8'd242; b_mant3 = 8'd111;
a_exp0 = 10'd735; a_exp1 = 10'd428; a_exp2 = 10'd480; a_exp3 = 10'd1016;
b_exp0 = 10'd159; b_exp1 = 10'd512; b_exp2 = 10'd481; b_exp3 = 10'd900;
a_sign0 = 4'd4; a_sign1 = 4'd12; a_sign2 = 4'd9; a_sign3 = 4'd8;
b_sign0 = 4'd3; b_sign1 = 4'd11; b_sign2 = 4'd5; b_sign3 = 4'd15;
@(posedge clk_i);
a_mant0 = 8'd87; a_mant1 = 8'd250; a_mant2 = 8'd88; a_mant3 = 8'd137;
b_mant0 = 8'd137; b_mant1 = 8'd190; b_mant2 = 8'd104; b_mant3 = 8'd89;
a_exp0 = 10'd757; a_exp1 = 10'd815; a_exp2 = 10'd173; a_exp3 = 10'd207;
b_exp0 = 10'd236; b_exp1 = 10'd840; b_exp2 = 10'd172; b_exp3 = 10'd982;
a_sign0 = 4'd12; a_sign1 = 4'd15; a_sign2 = 4'd13; a_sign3 = 4'd8;
b_sign0 = 4'd16; b_sign1 = 4'd7; b_sign2 = 4'd6; b_sign3 = 4'd12;
@(posedge clk_i);
a_mant0 = 8'd69; a_mant1 = 8'd55; a_mant2 = 8'd188; a_mant3 = 8'd199;
b_mant0 = 8'd89; b_mant1 = 8'd200; b_mant2 = 8'd166; b_mant3 = 8'd198;
a_exp0 = 10'd67; a_exp1 = 10'd382; a_exp2 = 10'd565; a_exp3 = 10'd829;
b_exp0 = 10'd545; b_exp1 = 10'd879; b_exp2 = 10'd584; b_exp3 = 10'd951;
a_sign0 = 4'd11; a_sign1 = 4'd3; a_sign2 = 4'd4; a_sign3 = 4'd0;
b_sign0 = 4'd0; b_sign1 = 4'd4; b_sign2 = 4'd7; b_sign3 = 4'd15;
@(posedge clk_i);
a_mant0 = 8'd224; a_mant1 = 8'd178; a_mant2 = 8'd188; a_mant3 = 8'd56;
b_mant0 = 8'd186; b_mant1 = 8'd124; b_mant2 = 8'd20; b_mant3 = 8'd111;
a_exp0 = 10'd770; a_exp1 = 10'd505; a_exp2 = 10'd714; a_exp3 = 10'd382;
b_exp0 = 10'd220; b_exp1 = 10'd750; b_exp2 = 10'd254; b_exp3 = 10'd586;
a_sign0 = 4'd3; a_sign1 = 4'd9; a_sign2 = 4'd5; a_sign3 = 4'd9;
b_sign0 = 4'd0; b_sign1 = 4'd1; b_sign2 = 4'd6; b_sign3 = 4'd9;
@(posedge clk_i);
shared_exps0 = 8'd120;
shared_exps1 = 8'd151;
a_mant0 = 8'd13; a_mant1 = 8'd120; a_mant2 = 8'd198; a_mant3 = 8'd43;
b_mant0 = 8'd39; b_mant1 = 8'd83; b_mant2 = 8'd222; b_mant3 = 8'd169;
a_exp0 = 10'd347; a_exp1 = 10'd704; a_exp2 = 10'd823; a_exp3 = 10'd662;
b_exp0 = 10'd762; b_exp1 = 10'd581; b_exp2 = 10'd451; b_exp3 = 10'd496;
a_sign0 = 4'd6; a_sign1 = 4'd1; a_sign2 = 4'd16; a_sign3 = 4'd5;
b_sign0 = 4'd14; b_sign1 = 4'd12; b_sign2 = 4'd16; b_sign3 = 4'd14;
@(posedge clk_i);
a_mant0 = 8'd53; a_mant1 = 8'd91; a_mant2 = 8'd14; a_mant3 = 8'd159;
b_mant0 = 8'd107; b_mant1 = 8'd164; b_mant2 = 8'd243; b_mant3 = 8'd182;
a_exp0 = 10'd451; a_exp1 = 10'd934; a_exp2 = 10'd467; a_exp3 = 10'd242;
b_exp0 = 10'd190; b_exp1 = 10'd115; b_exp2 = 10'd876; b_exp3 = 10'd609;
a_sign0 = 4'd0; a_sign1 = 4'd11; a_sign2 = 4'd6; a_sign3 = 4'd4;
b_sign0 = 4'd7; b_sign1 = 4'd9; b_sign2 = 4'd14; b_sign3 = 4'd10;
@(posedge clk_i);
a_mant0 = 8'd113; a_mant1 = 8'd92; a_mant2 = 8'd66; a_mant3 = 8'd154;
b_mant0 = 8'd174; b_mant1 = 8'd194; b_mant2 = 8'd126; b_mant3 = 8'd77;
a_exp0 = 10'd527; a_exp1 = 10'd516; a_exp2 = 10'd536; a_exp3 = 10'd946;
b_exp0 = 10'd828; b_exp1 = 10'd35; b_exp2 = 10'd947; b_exp3 = 10'd656;
a_sign0 = 4'd9; a_sign1 = 4'd8; a_sign2 = 4'd10; a_sign3 = 4'd3;
b_sign0 = 4'd0; b_sign1 = 4'd9; b_sign2 = 4'd15; b_sign3 = 4'd3;
@(posedge clk_i);
a_mant0 = 8'd107; a_mant1 = 8'd152; a_mant2 = 8'd174; a_mant3 = 8'd135;
b_mant0 = 8'd124; b_mant1 = 8'd244; b_mant2 = 8'd38; b_mant3 = 8'd150;
a_exp0 = 10'd710; a_exp1 = 10'd19; a_exp2 = 10'd731; a_exp3 = 10'd704;
b_exp0 = 10'd139; b_exp1 = 10'd1008; b_exp2 = 10'd614; b_exp3 = 10'd969;
a_sign0 = 4'd16; a_sign1 = 4'd13; a_sign2 = 4'd13; a_sign3 = 4'd13;
b_sign0 = 4'd5; b_sign1 = 4'd0; b_sign2 = 4'd3; b_sign3 = 4'd15;
@(posedge clk_i);
a_mant0 = 8'd140; a_mant1 = 8'd248; a_mant2 = 8'd159; a_mant3 = 8'd45;
b_mant0 = 8'd200; b_mant1 = 8'd107; b_mant2 = 8'd82; b_mant3 = 8'd246;
a_exp0 = 10'd176; a_exp1 = 10'd676; a_exp2 = 10'd866; a_exp3 = 10'd611;
b_exp0 = 10'd705; b_exp1 = 10'd798; b_exp2 = 10'd720; b_exp3 = 10'd585;
a_sign0 = 4'd12; a_sign1 = 4'd8; a_sign2 = 4'd3; a_sign3 = 4'd6;
b_sign0 = 4'd7; b_sign1 = 4'd13; b_sign2 = 4'd5; b_sign3 = 4'd7;
@(posedge clk_i);
a_mant0 = 8'd16; a_mant1 = 8'd11; a_mant2 = 8'd231; a_mant3 = 8'd87;
b_mant0 = 8'd10; b_mant1 = 8'd193; b_mant2 = 8'd112; b_mant3 = 8'd131;
a_exp0 = 10'd166; a_exp1 = 10'd862; a_exp2 = 10'd480; a_exp3 = 10'd121;
b_exp0 = 10'd318; b_exp1 = 10'd52; b_exp2 = 10'd80; b_exp3 = 10'd712;
a_sign0 = 4'd4; a_sign1 = 4'd2; a_sign2 = 4'd5; a_sign3 = 4'd3;
b_sign0 = 4'd8; b_sign1 = 4'd9; b_sign2 = 4'd5; b_sign3 = 4'd14;
@(posedge clk_i);
a_mant0 = 8'd55; a_mant1 = 8'd142; a_mant2 = 8'd150; a_mant3 = 8'd188;
b_mant0 = 8'd9; b_mant1 = 8'd182; b_mant2 = 8'd251; b_mant3 = 8'd67;
a_exp0 = 10'd343; a_exp1 = 10'd562; a_exp2 = 10'd710; a_exp3 = 10'd793;
b_exp0 = 10'd195; b_exp1 = 10'd681; b_exp2 = 10'd911; b_exp3 = 10'd684;
a_sign0 = 4'd8; a_sign1 = 4'd12; a_sign2 = 4'd15; a_sign3 = 4'd0;
b_sign0 = 4'd8; b_sign1 = 4'd16; b_sign2 = 4'd8; b_sign3 = 4'd9;
@(posedge clk_i);
a_mant0 = 8'd193; a_mant1 = 8'd151; a_mant2 = 8'd254; a_mant3 = 8'd65;
b_mant0 = 8'd226; b_mant1 = 8'd3; b_mant2 = 8'd82; b_mant3 = 8'd202;
a_exp0 = 10'd796; a_exp1 = 10'd776; a_exp2 = 10'd624; a_exp3 = 10'd157;
b_exp0 = 10'd375; b_exp1 = 10'd15; b_exp2 = 10'd332; b_exp3 = 10'd420;
a_sign0 = 4'd11; a_sign1 = 4'd0; a_sign2 = 4'd11; a_sign3 = 4'd11;
b_sign0 = 4'd9; b_sign1 = 4'd7; b_sign2 = 4'd5; b_sign3 = 4'd15;
@(posedge clk_i);
shared_exps0 = 8'd130;
shared_exps1 = 8'd95;
a_mant0 = 8'd89; a_mant1 = 8'd23; a_mant2 = 8'd203; a_mant3 = 8'd46;
b_mant0 = 8'd174; b_mant1 = 8'd232; b_mant2 = 8'd122; b_mant3 = 8'd239;
a_exp0 = 10'd154; a_exp1 = 10'd673; a_exp2 = 10'd1006; a_exp3 = 10'd765;
b_exp0 = 10'd363; b_exp1 = 10'd839; b_exp2 = 10'd738; b_exp3 = 10'd953;
a_sign0 = 4'd3; a_sign1 = 4'd1; a_sign2 = 4'd13; a_sign3 = 4'd7;
b_sign0 = 4'd5; b_sign1 = 4'd0; b_sign2 = 4'd12; b_sign3 = 4'd13;
@(posedge clk_i);
a_mant0 = 8'd105; a_mant1 = 8'd52; a_mant2 = 8'd249; a_mant3 = 8'd39;
b_mant0 = 8'd128; b_mant1 = 8'd14; b_mant2 = 8'd170; b_mant3 = 8'd25;
a_exp0 = 10'd873; a_exp1 = 10'd503; a_exp2 = 10'd546; a_exp3 = 10'd670;
b_exp0 = 10'd265; b_exp1 = 10'd674; b_exp2 = 10'd534; b_exp3 = 10'd436;
a_sign0 = 4'd11; a_sign1 = 4'd1; a_sign2 = 4'd10; a_sign3 = 4'd8;
b_sign0 = 4'd3; b_sign1 = 4'd3; b_sign2 = 4'd15; b_sign3 = 4'd2;
@(posedge clk_i);
a_mant0 = 8'd97; a_mant1 = 8'd219; a_mant2 = 8'd42; a_mant3 = 8'd246;
b_mant0 = 8'd231; b_mant1 = 8'd183; b_mant2 = 8'd86; b_mant3 = 8'd193;
a_exp0 = 10'd537; a_exp1 = 10'd738; a_exp2 = 10'd26; a_exp3 = 10'd641;
b_exp0 = 10'd30; b_exp1 = 10'd524; b_exp2 = 10'd495; b_exp3 = 10'd707;
a_sign0 = 4'd15; a_sign1 = 4'd9; a_sign2 = 4'd12; a_sign3 = 4'd9;
b_sign0 = 4'd6; b_sign1 = 4'd3; b_sign2 = 4'd6; b_sign3 = 4'd4;
@(posedge clk_i);
a_mant0 = 8'd202; a_mant1 = 8'd244; a_mant2 = 8'd144; a_mant3 = 8'd173;
b_mant0 = 8'd227; b_mant1 = 8'd92; b_mant2 = 8'd207; b_mant3 = 8'd225;
a_exp0 = 10'd485; a_exp1 = 10'd803; a_exp2 = 10'd186; a_exp3 = 10'd626;
b_exp0 = 10'd97; b_exp1 = 10'd522; b_exp2 = 10'd257; b_exp3 = 10'd567;
a_sign0 = 4'd16; a_sign1 = 4'd3; a_sign2 = 4'd14; a_sign3 = 4'd3;
b_sign0 = 4'd7; b_sign1 = 4'd9; b_sign2 = 4'd6; b_sign3 = 4'd4;
@(posedge clk_i);
a_mant0 = 8'd97; a_mant1 = 8'd123; a_mant2 = 8'd51; a_mant3 = 8'd148;
b_mant0 = 8'd71; b_mant1 = 8'd156; b_mant2 = 8'd169; b_mant3 = 8'd183;
a_exp0 = 10'd962; a_exp1 = 10'd358; a_exp2 = 10'd865; a_exp3 = 10'd263;
b_exp0 = 10'd398; b_exp1 = 10'd223; b_exp2 = 10'd472; b_exp3 = 10'd715;
a_sign0 = 4'd1; a_sign1 = 4'd16; a_sign2 = 4'd6; a_sign3 = 4'd1;
b_sign0 = 4'd13; b_sign1 = 4'd15; b_sign2 = 4'd9; b_sign3 = 4'd8;
@(posedge clk_i);
a_mant0 = 8'd66; a_mant1 = 8'd212; a_mant2 = 8'd124; a_mant3 = 8'd236;
b_mant0 = 8'd122; b_mant1 = 8'd209; b_mant2 = 8'd100; b_mant3 = 8'd140;
a_exp0 = 10'd268; a_exp1 = 10'd236; a_exp2 = 10'd806; a_exp3 = 10'd911;
b_exp0 = 10'd181; b_exp1 = 10'd500; b_exp2 = 10'd166; b_exp3 = 10'd791;
a_sign0 = 4'd12; a_sign1 = 4'd12; a_sign2 = 4'd13; a_sign3 = 4'd3;
b_sign0 = 4'd0; b_sign1 = 4'd15; b_sign2 = 4'd1; b_sign3 = 4'd8;
@(posedge clk_i);
a_mant0 = 8'd179; a_mant1 = 8'd80; a_mant2 = 8'd72; a_mant3 = 8'd120;
b_mant0 = 8'd120; b_mant1 = 8'd206; b_mant2 = 8'd144; b_mant3 = 8'd11;
a_exp0 = 10'd346; a_exp1 = 10'd752; a_exp2 = 10'd760; a_exp3 = 10'd52;
b_exp0 = 10'd7; b_exp1 = 10'd715; b_exp2 = 10'd349; b_exp3 = 10'd537;
a_sign0 = 4'd2; a_sign1 = 4'd7; a_sign2 = 4'd7; a_sign3 = 4'd15;
b_sign0 = 4'd12; b_sign1 = 4'd5; b_sign2 = 4'd3; b_sign3 = 4'd5;
@(posedge clk_i);
a_mant0 = 8'd166; a_mant1 = 8'd37; a_mant2 = 8'd168; a_mant3 = 8'd27;
b_mant0 = 8'd89; b_mant1 = 8'd44; b_mant2 = 8'd251; b_mant3 = 8'd82;
a_exp0 = 10'd81; a_exp1 = 10'd267; a_exp2 = 10'd801; a_exp3 = 10'd966;
b_exp0 = 10'd654; b_exp1 = 10'd119; b_exp2 = 10'd184; b_exp3 = 10'd384;
a_sign0 = 4'd1; a_sign1 = 4'd9; a_sign2 = 4'd6; a_sign3 = 4'd3;
b_sign0 = 4'd10; b_sign1 = 4'd12; b_sign2 = 4'd8; b_sign3 = 4'd10;
@(posedge clk_i);
shared_exps0 = 8'd138;
shared_exps1 = 8'd131;
rstn = 0;
@(posedge clk_i);
rstn = 1;
a_mant0 = 8'd65; a_mant1 = 8'd159; a_mant2 = 8'd34; a_mant3 = 8'd110;
b_mant0 = 8'd158; b_mant1 = 8'd186; b_mant2 = 8'd134; b_mant3 = 8'd223;
a_exp0 = 10'd775; a_exp1 = 10'd797; a_exp2 = 10'd303; a_exp3 = 10'd482;
b_exp0 = 10'd551; b_exp1 = 10'd484; b_exp2 = 10'd771; b_exp3 = 10'd723;
a_sign0 = 4'd8; a_sign1 = 4'd9; a_sign2 = 4'd16; a_sign3 = 4'd16;
b_sign0 = 4'd13; b_sign1 = 4'd11; b_sign2 = 4'd3; b_sign3 = 4'd4;
@(posedge clk_i);
a_mant0 = 8'd72; a_mant1 = 8'd222; a_mant2 = 8'd250; a_mant3 = 8'd53;
b_mant0 = 8'd15; b_mant1 = 8'd166; b_mant2 = 8'd50; b_mant3 = 8'd245;
a_exp0 = 10'd608; a_exp1 = 10'd163; a_exp2 = 10'd639; a_exp3 = 10'd478;
b_exp0 = 10'd75; b_exp1 = 10'd132; b_exp2 = 10'd331; b_exp3 = 10'd236;
a_sign0 = 4'd5; a_sign1 = 4'd3; a_sign2 = 4'd0; a_sign3 = 4'd11;
b_sign0 = 4'd10; b_sign1 = 4'd13; b_sign2 = 4'd8; b_sign3 = 4'd10;
@(posedge clk_i);
a_mant0 = 8'd148; a_mant1 = 8'd151; a_mant2 = 8'd20; a_mant3 = 8'd218;
b_mant0 = 8'd100; b_mant1 = 8'd211; b_mant2 = 8'd70; b_mant3 = 8'd21;
a_exp0 = 10'd130; a_exp1 = 10'd862; a_exp2 = 10'd108; a_exp3 = 10'd63;
b_exp0 = 10'd747; b_exp1 = 10'd15; b_exp2 = 10'd317; b_exp3 = 10'd759;
a_sign0 = 4'd14; a_sign1 = 4'd3; a_sign2 = 4'd13; a_sign3 = 4'd6;
b_sign0 = 4'd6; b_sign1 = 4'd16; b_sign2 = 4'd3; b_sign3 = 4'd2;
@(posedge clk_i);
a_mant0 = 8'd74; a_mant1 = 8'd190; a_mant2 = 8'd192; a_mant3 = 8'd93;
b_mant0 = 8'd204; b_mant1 = 8'd24; b_mant2 = 8'd50; b_mant3 = 8'd140;
a_exp0 = 10'd956; a_exp1 = 10'd149; a_exp2 = 10'd17; a_exp3 = 10'd114;
b_exp0 = 10'd426; b_exp1 = 10'd733; b_exp2 = 10'd299; b_exp3 = 10'd370;
a_sign0 = 4'd11; a_sign1 = 4'd8; a_sign2 = 4'd16; a_sign3 = 4'd11;
b_sign0 = 4'd9; b_sign1 = 4'd1; b_sign2 = 4'd12; b_sign3 = 4'd2;
@(posedge clk_i);
a_mant0 = 8'd81; a_mant1 = 8'd203; a_mant2 = 8'd111; a_mant3 = 8'd56;
b_mant0 = 8'd218; b_mant1 = 8'd3; b_mant2 = 8'd71; b_mant3 = 8'd19;
a_exp0 = 10'd931; a_exp1 = 10'd406; a_exp2 = 10'd67; a_exp3 = 10'd335;
b_exp0 = 10'd461; b_exp1 = 10'd1009; b_exp2 = 10'd895; b_exp3 = 10'd569;
a_sign0 = 4'd6; a_sign1 = 4'd4; a_sign2 = 4'd3; a_sign3 = 4'd16;
b_sign0 = 4'd11; b_sign1 = 4'd3; b_sign2 = 4'd12; b_sign3 = 4'd14;
@(posedge clk_i);
a_mant0 = 8'd205; a_mant1 = 8'd111; a_mant2 = 8'd67; a_mant3 = 8'd238;
b_mant0 = 8'd125; b_mant1 = 8'd180; b_mant2 = 8'd253; b_mant3 = 8'd167;
a_exp0 = 10'd556; a_exp1 = 10'd608; a_exp2 = 10'd651; a_exp3 = 10'd530;
b_exp0 = 10'd1018; b_exp1 = 10'd172; b_exp2 = 10'd95; b_exp3 = 10'd668;
a_sign0 = 4'd9; a_sign1 = 4'd1; a_sign2 = 4'd7; a_sign3 = 4'd15;
b_sign0 = 4'd13; b_sign1 = 4'd15; b_sign2 = 4'd16; b_sign3 = 4'd15;
@(posedge clk_i);
a_mant0 = 8'd189; a_mant1 = 8'd149; a_mant2 = 8'd34; a_mant3 = 8'd106;
b_mant0 = 8'd164; b_mant1 = 8'd185; b_mant2 = 8'd118; b_mant3 = 8'd59;
a_exp0 = 10'd681; a_exp1 = 10'd664; a_exp2 = 10'd145; a_exp3 = 10'd898;
b_exp0 = 10'd339; b_exp1 = 10'd38; b_exp2 = 10'd0; b_exp3 = 10'd436;
a_sign0 = 4'd2; a_sign1 = 4'd3; a_sign2 = 4'd7; a_sign3 = 4'd10;
b_sign0 = 4'd16; b_sign1 = 4'd12; b_sign2 = 4'd8; b_sign3 = 4'd11;
@(posedge clk_i);
shared_exps0 = 8'd122;
shared_exps1 = 8'd123;
a_mant0 = 8'd222; a_mant1 = 8'd254; a_mant2 = 8'd123; a_mant3 = 8'd154;
b_mant0 = 8'd116; b_mant1 = 8'd218; b_mant2 = 8'd234; b_mant3 = 8'd25;
a_exp0 = 10'd128; a_exp1 = 10'd692; a_exp2 = 10'd977; a_exp3 = 10'd830;
b_exp0 = 10'd672; b_exp1 = 10'd75; b_exp2 = 10'd43; b_exp3 = 10'd780;
a_sign0 = 4'd5; a_sign1 = 4'd9; a_sign2 = 4'd10; a_sign3 = 4'd14;
b_sign0 = 4'd0; b_sign1 = 4'd3; b_sign2 = 4'd14; b_sign3 = 4'd1;
@(posedge clk_i);
a_mant0 = 8'd33; a_mant1 = 8'd80; a_mant2 = 8'd87; a_mant3 = 8'd37;
b_mant0 = 8'd91; b_mant1 = 8'd179; b_mant2 = 8'd65; b_mant3 = 8'd14;
a_exp0 = 10'd1; a_exp1 = 10'd436; a_exp2 = 10'd178; a_exp3 = 10'd815;
b_exp0 = 10'd189; b_exp1 = 10'd849; b_exp2 = 10'd259; b_exp3 = 10'd380;
a_sign0 = 4'd5; a_sign1 = 4'd16; a_sign2 = 4'd6; a_sign3 = 4'd3;
b_sign0 = 4'd3; b_sign1 = 4'd1; b_sign2 = 4'd8; b_sign3 = 4'd11;
@(posedge clk_i);
a_mant0 = 8'd162; a_mant1 = 8'd168; a_mant2 = 8'd45; a_mant3 = 8'd62;
b_mant0 = 8'd1; b_mant1 = 8'd182; b_mant2 = 8'd85; b_mant3 = 8'd219;
a_exp0 = 10'd515; a_exp1 = 10'd227; a_exp2 = 10'd132; a_exp3 = 10'd474;
b_exp0 = 10'd318; b_exp1 = 10'd320; b_exp2 = 10'd785; b_exp3 = 10'd288;
a_sign0 = 4'd14; a_sign1 = 4'd0; a_sign2 = 4'd12; a_sign3 = 4'd0;
b_sign0 = 4'd9; b_sign1 = 4'd3; b_sign2 = 4'd13; b_sign3 = 4'd16;
@(posedge clk_i);
a_mant0 = 8'd15; a_mant1 = 8'd102; a_mant2 = 8'd151; a_mant3 = 8'd138;
b_mant0 = 8'd206; b_mant1 = 8'd77; b_mant2 = 8'd116; b_mant3 = 8'd20;
a_exp0 = 10'd774; a_exp1 = 10'd784; a_exp2 = 10'd614; a_exp3 = 10'd628;
b_exp0 = 10'd607; b_exp1 = 10'd234; b_exp2 = 10'd1020; b_exp3 = 10'd816;
a_sign0 = 4'd6; a_sign1 = 4'd0; a_sign2 = 4'd7; a_sign3 = 4'd12;
b_sign0 = 4'd15; b_sign1 = 4'd15; b_sign2 = 4'd10; b_sign3 = 4'd10;
@(posedge clk_i);
a_mant0 = 8'd247; a_mant1 = 8'd139; a_mant2 = 8'd68; a_mant3 = 8'd171;
b_mant0 = 8'd241; b_mant1 = 8'd108; b_mant2 = 8'd195; b_mant3 = 8'd198;
a_exp0 = 10'd94; a_exp1 = 10'd482; a_exp2 = 10'd1021; a_exp3 = 10'd613;
b_exp0 = 10'd984; b_exp1 = 10'd592; b_exp2 = 10'd837; b_exp3 = 10'd129;
a_sign0 = 4'd15; a_sign1 = 4'd14; a_sign2 = 4'd14; a_sign3 = 4'd1;
b_sign0 = 4'd0; b_sign1 = 4'd16; b_sign2 = 4'd14; b_sign3 = 4'd6;
@(posedge clk_i);
a_mant0 = 8'd67; a_mant1 = 8'd88; a_mant2 = 8'd12; a_mant3 = 8'd5;
b_mant0 = 8'd122; b_mant1 = 8'd65; b_mant2 = 8'd36; b_mant3 = 8'd162;
a_exp0 = 10'd161; a_exp1 = 10'd83; a_exp2 = 10'd631; a_exp3 = 10'd873;
b_exp0 = 10'd148; b_exp1 = 10'd179; b_exp2 = 10'd958; b_exp3 = 10'd758;
a_sign0 = 4'd0; a_sign1 = 4'd0; a_sign2 = 4'd12; a_sign3 = 4'd7;
b_sign0 = 4'd6; b_sign1 = 4'd7; b_sign2 = 4'd11; b_sign3 = 4'd9;
@(posedge clk_i);
a_mant0 = 8'd44; a_mant1 = 8'd218; a_mant2 = 8'd128; a_mant3 = 8'd149;
b_mant0 = 8'd23; b_mant1 = 8'd91; b_mant2 = 8'd48; b_mant3 = 8'd252;
a_exp0 = 10'd912; a_exp1 = 10'd479; a_exp2 = 10'd794; a_exp3 = 10'd670;
b_exp0 = 10'd430; b_exp1 = 10'd120; b_exp2 = 10'd270; b_exp3 = 10'd280;
a_sign0 = 4'd5; a_sign1 = 4'd12; a_sign2 = 4'd6; a_sign3 = 4'd3;
b_sign0 = 4'd11; b_sign1 = 4'd12; b_sign2 = 4'd8; b_sign3 = 4'd15;
@(posedge clk_i);
a_mant0 = 8'd182; a_mant1 = 8'd85; a_mant2 = 8'd152; a_mant3 = 8'd231;
b_mant0 = 8'd195; b_mant1 = 8'd126; b_mant2 = 8'd206; b_mant3 = 8'd112;
a_exp0 = 10'd471; a_exp1 = 10'd955; a_exp2 = 10'd685; a_exp3 = 10'd991;
b_exp0 = 10'd105; b_exp1 = 10'd156; b_exp2 = 10'd274; b_exp3 = 10'd79;
a_sign0 = 4'd7; a_sign1 = 4'd2; a_sign2 = 4'd2; a_sign3 = 4'd0;
b_sign0 = 4'd8; b_sign1 = 4'd13; b_sign2 = 4'd7; b_sign3 = 4'd10;
@(posedge clk_i);
shared_exps0 = 8'd126;
shared_exps1 = 8'd115;
a_mant0 = 8'd223; a_mant1 = 8'd172; a_mant2 = 8'd167; a_mant3 = 8'd254;
b_mant0 = 8'd81; b_mant1 = 8'd253; b_mant2 = 8'd46; b_mant3 = 8'd16;
a_exp0 = 10'd995; a_exp1 = 10'd68; a_exp2 = 10'd644; a_exp3 = 10'd1010;
b_exp0 = 10'd678; b_exp1 = 10'd1015; b_exp2 = 10'd242; b_exp3 = 10'd104;
a_sign0 = 4'd15; a_sign1 = 4'd0; a_sign2 = 4'd4; a_sign3 = 4'd4;
b_sign0 = 4'd2; b_sign1 = 4'd1; b_sign2 = 4'd15; b_sign3 = 4'd4;
@(posedge clk_i);
a_mant0 = 8'd185; a_mant1 = 8'd244; a_mant2 = 8'd32; a_mant3 = 8'd223;
b_mant0 = 8'd182; b_mant1 = 8'd202; b_mant2 = 8'd136; b_mant3 = 8'd109;
a_exp0 = 10'd598; a_exp1 = 10'd694; a_exp2 = 10'd765; a_exp3 = 10'd349;
b_exp0 = 10'd208; b_exp1 = 10'd217; b_exp2 = 10'd527; b_exp3 = 10'd471;
a_sign0 = 4'd2; a_sign1 = 4'd1; a_sign2 = 4'd2; a_sign3 = 4'd7;
b_sign0 = 4'd9; b_sign1 = 4'd0; b_sign2 = 4'd10; b_sign3 = 4'd11;
@(posedge clk_i);
a_mant0 = 8'd80; a_mant1 = 8'd82; a_mant2 = 8'd83; a_mant3 = 8'd110;
b_mant0 = 8'd95; b_mant1 = 8'd147; b_mant2 = 8'd118; b_mant3 = 8'd199;
a_exp0 = 10'd400; a_exp1 = 10'd219; a_exp2 = 10'd18; a_exp3 = 10'd287;
b_exp0 = 10'd91; b_exp1 = 10'd999; b_exp2 = 10'd382; b_exp3 = 10'd547;
a_sign0 = 4'd7; a_sign1 = 4'd9; a_sign2 = 4'd4; a_sign3 = 4'd3;
b_sign0 = 4'd4; b_sign1 = 4'd16; b_sign2 = 4'd0; b_sign3 = 4'd0;
@(posedge clk_i);
a_mant0 = 8'd36; a_mant1 = 8'd101; a_mant2 = 8'd197; a_mant3 = 8'd144;
b_mant0 = 8'd144; b_mant1 = 8'd113; b_mant2 = 8'd246; b_mant3 = 8'd75;
a_exp0 = 10'd974; a_exp1 = 10'd78; a_exp2 = 10'd596; a_exp3 = 10'd88;
b_exp0 = 10'd815; b_exp1 = 10'd866; b_exp2 = 10'd587; b_exp3 = 10'd726;
a_sign0 = 4'd12; a_sign1 = 4'd16; a_sign2 = 4'd12; a_sign3 = 4'd0;
b_sign0 = 4'd7; b_sign1 = 4'd6; b_sign2 = 4'd14; b_sign3 = 4'd11;
@(posedge clk_i);
a_mant0 = 8'd46; a_mant1 = 8'd172; a_mant2 = 8'd228; a_mant3 = 8'd165;
b_mant0 = 8'd174; b_mant1 = 8'd77; b_mant2 = 8'd237; b_mant3 = 8'd213;
a_exp0 = 10'd420; a_exp1 = 10'd419; a_exp2 = 10'd500; a_exp3 = 10'd399;
b_exp0 = 10'd576; b_exp1 = 10'd943; b_exp2 = 10'd367; b_exp3 = 10'd958;
a_sign0 = 4'd1; a_sign1 = 4'd8; a_sign2 = 4'd0; a_sign3 = 4'd5;
b_sign0 = 4'd14; b_sign1 = 4'd6; b_sign2 = 4'd5; b_sign3 = 4'd5;
@(posedge clk_i);
a_mant0 = 8'd127; a_mant1 = 8'd190; a_mant2 = 8'd155; a_mant3 = 8'd217;
b_mant0 = 8'd190; b_mant1 = 8'd153; b_mant2 = 8'd101; b_mant3 = 8'd101;
a_exp0 = 10'd546; a_exp1 = 10'd461; a_exp2 = 10'd600; a_exp3 = 10'd607;
b_exp0 = 10'd412; b_exp1 = 10'd106; b_exp2 = 10'd534; b_exp3 = 10'd63;
a_sign0 = 4'd4; a_sign1 = 4'd1; a_sign2 = 4'd6; a_sign3 = 4'd11;
b_sign0 = 4'd8; b_sign1 = 4'd9; b_sign2 = 4'd9; b_sign3 = 4'd7;
@(posedge clk_i);
a_mant0 = 8'd34; a_mant1 = 8'd114; a_mant2 = 8'd121; a_mant3 = 8'd184;
b_mant0 = 8'd213; b_mant1 = 8'd132; b_mant2 = 8'd50; b_mant3 = 8'd91;
a_exp0 = 10'd55; a_exp1 = 10'd699; a_exp2 = 10'd974; a_exp3 = 10'd289;
b_exp0 = 10'd738; b_exp1 = 10'd866; b_exp2 = 10'd466; b_exp3 = 10'd1;
a_sign0 = 4'd3; a_sign1 = 4'd9; a_sign2 = 4'd3; a_sign3 = 4'd4;
b_sign0 = 4'd15; b_sign1 = 4'd10; b_sign2 = 4'd16; b_sign3 = 4'd14;
@(posedge clk_i);
a_mant0 = 8'd162; a_mant1 = 8'd254; a_mant2 = 8'd62; a_mant3 = 8'd175;
b_mant0 = 8'd10; b_mant1 = 8'd148; b_mant2 = 8'd157; b_mant3 = 8'd45;
a_exp0 = 10'd729; a_exp1 = 10'd551; a_exp2 = 10'd683; a_exp3 = 10'd549;
b_exp0 = 10'd695; b_exp1 = 10'd40; b_exp2 = 10'd793; b_exp3 = 10'd832;
a_sign0 = 4'd14; a_sign1 = 4'd7; a_sign2 = 4'd14; a_sign3 = 4'd11;
b_sign0 = 4'd15; b_sign1 = 4'd13; b_sign2 = 4'd5; b_sign3 = 4'd4;
@(posedge clk_i);
shared_exps0 = 8'd135;
shared_exps1 = 8'd144;
a_mant0 = 8'd57; a_mant1 = 8'd164; a_mant2 = 8'd10; a_mant3 = 8'd206;
b_mant0 = 8'd247; b_mant1 = 8'd6; b_mant2 = 8'd175; b_mant3 = 8'd1;
a_exp0 = 10'd890; a_exp1 = 10'd725; a_exp2 = 10'd150; a_exp3 = 10'd368;
b_exp0 = 10'd731; b_exp1 = 10'd34; b_exp2 = 10'd713; b_exp3 = 10'd51;
a_sign0 = 4'd9; a_sign1 = 4'd3; a_sign2 = 4'd8; a_sign3 = 4'd12;
b_sign0 = 4'd15; b_sign1 = 4'd16; b_sign2 = 4'd3; b_sign3 = 4'd5;
@(posedge clk_i);
a_mant0 = 8'd10; a_mant1 = 8'd85; a_mant2 = 8'd104; a_mant3 = 8'd203;
b_mant0 = 8'd118; b_mant1 = 8'd1; b_mant2 = 8'd213; b_mant3 = 8'd61;
a_exp0 = 10'd406; a_exp1 = 10'd590; a_exp2 = 10'd323; a_exp3 = 10'd590;
b_exp0 = 10'd110; b_exp1 = 10'd180; b_exp2 = 10'd538; b_exp3 = 10'd117;
a_sign0 = 4'd12; a_sign1 = 4'd4; a_sign2 = 4'd14; a_sign3 = 4'd10;
b_sign0 = 4'd14; b_sign1 = 4'd5; b_sign2 = 4'd16; b_sign3 = 4'd15;
@(posedge clk_i);
a_mant0 = 8'd41; a_mant1 = 8'd91; a_mant2 = 8'd117; a_mant3 = 8'd5;
b_mant0 = 8'd135; b_mant1 = 8'd175; b_mant2 = 8'd11; b_mant3 = 8'd239;
a_exp0 = 10'd943; a_exp1 = 10'd553; a_exp2 = 10'd844; a_exp3 = 10'd652;
b_exp0 = 10'd923; b_exp1 = 10'd591; b_exp2 = 10'd403; b_exp3 = 10'd505;
a_sign0 = 4'd10; a_sign1 = 4'd6; a_sign2 = 4'd13; a_sign3 = 4'd0;
b_sign0 = 4'd6; b_sign1 = 4'd5; b_sign2 = 4'd0; b_sign3 = 4'd15;
@(posedge clk_i);
a_mant0 = 8'd25; a_mant1 = 8'd92; a_mant2 = 8'd17; a_mant3 = 8'd240;
b_mant0 = 8'd201; b_mant1 = 8'd143; b_mant2 = 8'd121; b_mant3 = 8'd128;
a_exp0 = 10'd325; a_exp1 = 10'd699; a_exp2 = 10'd377; a_exp3 = 10'd988;
b_exp0 = 10'd590; b_exp1 = 10'd989; b_exp2 = 10'd199; b_exp3 = 10'd190;
a_sign0 = 4'd16; a_sign1 = 4'd1; a_sign2 = 4'd8; a_sign3 = 4'd15;
b_sign0 = 4'd11; b_sign1 = 4'd4; b_sign2 = 4'd3; b_sign3 = 4'd1;
@(posedge clk_i);
a_mant0 = 8'd97; a_mant1 = 8'd107; a_mant2 = 8'd44; a_mant3 = 8'd178;
b_mant0 = 8'd69; b_mant1 = 8'd183; b_mant2 = 8'd51; b_mant3 = 8'd236;
a_exp0 = 10'd12; a_exp1 = 10'd131; a_exp2 = 10'd845; a_exp3 = 10'd728;
b_exp0 = 10'd580; b_exp1 = 10'd92; b_exp2 = 10'd166; b_exp3 = 10'd625;
a_sign0 = 4'd4; a_sign1 = 4'd12; a_sign2 = 4'd13; a_sign3 = 4'd11;
b_sign0 = 4'd14; b_sign1 = 4'd2; b_sign2 = 4'd0; b_sign3 = 4'd11;
@(posedge clk_i);
a_mant0 = 8'd198; a_mant1 = 8'd249; a_mant2 = 8'd189; a_mant3 = 8'd84;
b_mant0 = 8'd209; b_mant1 = 8'd197; b_mant2 = 8'd4; b_mant3 = 8'd48;
a_exp0 = 10'd167; a_exp1 = 10'd704; a_exp2 = 10'd519; a_exp3 = 10'd609;
b_exp0 = 10'd901; b_exp1 = 10'd674; b_exp2 = 10'd243; b_exp3 = 10'd206;
a_sign0 = 4'd5; a_sign1 = 4'd14; a_sign2 = 4'd5; a_sign3 = 4'd11;
b_sign0 = 4'd2; b_sign1 = 4'd7; b_sign2 = 4'd14; b_sign3 = 4'd13;
@(posedge clk_i);
a_mant0 = 8'd117; a_mant1 = 8'd223; a_mant2 = 8'd119; a_mant3 = 8'd218;
b_mant0 = 8'd78; b_mant1 = 8'd249; b_mant2 = 8'd253; b_mant3 = 8'd86;
a_exp0 = 10'd546; a_exp1 = 10'd925; a_exp2 = 10'd579; a_exp3 = 10'd486;
b_exp0 = 10'd221; b_exp1 = 10'd50; b_exp2 = 10'd961; b_exp3 = 10'd403;
a_sign0 = 4'd1; a_sign1 = 4'd8; a_sign2 = 4'd16; a_sign3 = 4'd3;
b_sign0 = 4'd11; b_sign1 = 4'd9; b_sign2 = 4'd0; b_sign3 = 4'd6;
@(posedge clk_i);
a_mant0 = 8'd115; a_mant1 = 8'd0; a_mant2 = 8'd3; a_mant3 = 8'd71;
b_mant0 = 8'd250; b_mant1 = 8'd229; b_mant2 = 8'd113; b_mant3 = 8'd159;
a_exp0 = 10'd33; a_exp1 = 10'd465; a_exp2 = 10'd714; a_exp3 = 10'd1007;
b_exp0 = 10'd592; b_exp1 = 10'd451; b_exp2 = 10'd654; b_exp3 = 10'd101;
a_sign0 = 4'd1; a_sign1 = 4'd16; a_sign2 = 4'd7; a_sign3 = 4'd12;
b_sign0 = 4'd12; b_sign1 = 4'd5; b_sign2 = 4'd3; b_sign3 = 4'd5;
@(posedge clk_i);
shared_exps0 = 8'd111;
shared_exps1 = 8'd129;
rstn = 0;
@(posedge clk_i);
rstn = 1;
a_mant0 = 8'd69; a_mant1 = 8'd226; a_mant2 = 8'd161; a_mant3 = 8'd188;
b_mant0 = 8'd183; b_mant1 = 8'd151; b_mant2 = 8'd94; b_mant3 = 8'd227;
a_exp0 = 10'd235; a_exp1 = 10'd467; a_exp2 = 10'd405; a_exp3 = 10'd744;
b_exp0 = 10'd262; b_exp1 = 10'd854; b_exp2 = 10'd9; b_exp3 = 10'd820;
a_sign0 = 4'd4; a_sign1 = 4'd8; a_sign2 = 4'd13; a_sign3 = 4'd6;
b_sign0 = 4'd11; b_sign1 = 4'd13; b_sign2 = 4'd3; b_sign3 = 4'd5;
@(posedge clk_i);
a_mant0 = 8'd222; a_mant1 = 8'd144; a_mant2 = 8'd206; a_mant3 = 8'd112;
b_mant0 = 8'd37; b_mant1 = 8'd55; b_mant2 = 8'd166; b_mant3 = 8'd120;
a_exp0 = 10'd952; a_exp1 = 10'd389; a_exp2 = 10'd412; a_exp3 = 10'd838;
b_exp0 = 10'd124; b_exp1 = 10'd853; b_exp2 = 10'd428; b_exp3 = 10'd125;
a_sign0 = 4'd11; a_sign1 = 4'd7; a_sign2 = 4'd6; a_sign3 = 4'd4;
b_sign0 = 4'd5; b_sign1 = 4'd15; b_sign2 = 4'd2; b_sign3 = 4'd2;
@(posedge clk_i);
a_mant0 = 8'd138; a_mant1 = 8'd13; a_mant2 = 8'd44; a_mant3 = 8'd80;
b_mant0 = 8'd135; b_mant1 = 8'd96; b_mant2 = 8'd132; b_mant3 = 8'd66;
a_exp0 = 10'd336; a_exp1 = 10'd782; a_exp2 = 10'd874; a_exp3 = 10'd17;
b_exp0 = 10'd303; b_exp1 = 10'd994; b_exp2 = 10'd112; b_exp3 = 10'd372;
a_sign0 = 4'd5; a_sign1 = 4'd2; a_sign2 = 4'd7; a_sign3 = 4'd14;
b_sign0 = 4'd5; b_sign1 = 4'd7; b_sign2 = 4'd5; b_sign3 = 4'd2;
@(posedge clk_i);
a_mant0 = 8'd20; a_mant1 = 8'd21; a_mant2 = 8'd192; a_mant3 = 8'd63;
b_mant0 = 8'd7; b_mant1 = 8'd129; b_mant2 = 8'd251; b_mant3 = 8'd194;
a_exp0 = 10'd737; a_exp1 = 10'd38; a_exp2 = 10'd620; a_exp3 = 10'd42;
b_exp0 = 10'd718; b_exp1 = 10'd302; b_exp2 = 10'd653; b_exp3 = 10'd719;
a_sign0 = 4'd14; a_sign1 = 4'd1; a_sign2 = 4'd12; a_sign3 = 4'd6;
b_sign0 = 4'd9; b_sign1 = 4'd12; b_sign2 = 4'd9; b_sign3 = 4'd7;
@(posedge clk_i);
a_mant0 = 8'd154; a_mant1 = 8'd61; a_mant2 = 8'd176; a_mant3 = 8'd165;
b_mant0 = 8'd162; b_mant1 = 8'd241; b_mant2 = 8'd85; b_mant3 = 8'd123;
a_exp0 = 10'd176; a_exp1 = 10'd90; a_exp2 = 10'd64; a_exp3 = 10'd204;
b_exp0 = 10'd676; b_exp1 = 10'd446; b_exp2 = 10'd94; b_exp3 = 10'd921;
a_sign0 = 4'd8; a_sign1 = 4'd7; a_sign2 = 4'd1; a_sign3 = 4'd13;
b_sign0 = 4'd2; b_sign1 = 4'd13; b_sign2 = 4'd9; b_sign3 = 4'd4;
@(posedge clk_i);
a_mant0 = 8'd177; a_mant1 = 8'd213; a_mant2 = 8'd189; a_mant3 = 8'd29;
b_mant0 = 8'd141; b_mant1 = 8'd177; b_mant2 = 8'd20; b_mant3 = 8'd185;
a_exp0 = 10'd773; a_exp1 = 10'd625; a_exp2 = 10'd116; a_exp3 = 10'd407;
b_exp0 = 10'd116; b_exp1 = 10'd377; b_exp2 = 10'd850; b_exp3 = 10'd349;
a_sign0 = 4'd14; a_sign1 = 4'd8; a_sign2 = 4'd14; a_sign3 = 4'd13;
b_sign0 = 4'd13; b_sign1 = 4'd14; b_sign2 = 4'd8; b_sign3 = 4'd4;
@(posedge clk_i);
a_mant0 = 8'd28; a_mant1 = 8'd81; a_mant2 = 8'd17; a_mant3 = 8'd83;
b_mant0 = 8'd221; b_mant1 = 8'd215; b_mant2 = 8'd2; b_mant3 = 8'd245;
a_exp0 = 10'd828; a_exp1 = 10'd322; a_exp2 = 10'd672; a_exp3 = 10'd416;
b_exp0 = 10'd968; b_exp1 = 10'd550; b_exp2 = 10'd504; b_exp3 = 10'd440;
a_sign0 = 4'd15; a_sign1 = 4'd8; a_sign2 = 4'd13; a_sign3 = 4'd15;
b_sign0 = 4'd16; b_sign1 = 4'd12; b_sign2 = 4'd15; b_sign3 = 4'd7;
@(posedge clk_i);
shared_exps0 = 8'd151;
shared_exps1 = 8'd99;
a_mant0 = 8'd81; a_mant1 = 8'd10; a_mant2 = 8'd123; a_mant3 = 8'd71;
b_mant0 = 8'd28; b_mant1 = 8'd2; b_mant2 = 8'd138; b_mant3 = 8'd92;
a_exp0 = 10'd304; a_exp1 = 10'd997; a_exp2 = 10'd488; a_exp3 = 10'd619;
b_exp0 = 10'd315; b_exp1 = 10'd175; b_exp2 = 10'd524; b_exp3 = 10'd817;
a_sign0 = 4'd13; a_sign1 = 4'd16; a_sign2 = 4'd9; a_sign3 = 4'd0;
b_sign0 = 4'd9; b_sign1 = 4'd15; b_sign2 = 4'd7; b_sign3 = 4'd15;
@(posedge clk_i);
a_mant0 = 8'd29; a_mant1 = 8'd123; a_mant2 = 8'd197; a_mant3 = 8'd117;
b_mant0 = 8'd243; b_mant1 = 8'd124; b_mant2 = 8'd249; b_mant3 = 8'd153;
a_exp0 = 10'd990; a_exp1 = 10'd367; a_exp2 = 10'd665; a_exp3 = 10'd426;
b_exp0 = 10'd97; b_exp1 = 10'd451; b_exp2 = 10'd795; b_exp3 = 10'd569;
a_sign0 = 4'd0; a_sign1 = 4'd15; a_sign2 = 4'd15; a_sign3 = 4'd3;
b_sign0 = 4'd8; b_sign1 = 4'd10; b_sign2 = 4'd10; b_sign3 = 4'd7;
@(posedge clk_i);
a_mant0 = 8'd180; a_mant1 = 8'd23; a_mant2 = 8'd48; a_mant3 = 8'd216;
b_mant0 = 8'd48; b_mant1 = 8'd66; b_mant2 = 8'd22; b_mant3 = 8'd81;
a_exp0 = 10'd312; a_exp1 = 10'd870; a_exp2 = 10'd44; a_exp3 = 10'd117;
b_exp0 = 10'd723; b_exp1 = 10'd812; b_exp2 = 10'd76; b_exp3 = 10'd690;
a_sign0 = 4'd12; a_sign1 = 4'd10; a_sign2 = 4'd6; a_sign3 = 4'd10;
b_sign0 = 4'd3; b_sign1 = 4'd0; b_sign2 = 4'd8; b_sign3 = 4'd10;
@(posedge clk_i);
a_mant0 = 8'd242; a_mant1 = 8'd123; a_mant2 = 8'd21; a_mant3 = 8'd45;
b_mant0 = 8'd31; b_mant1 = 8'd164; b_mant2 = 8'd196; b_mant3 = 8'd104;
a_exp0 = 10'd718; a_exp1 = 10'd719; a_exp2 = 10'd980; a_exp3 = 10'd86;
b_exp0 = 10'd147; b_exp1 = 10'd116; b_exp2 = 10'd432; b_exp3 = 10'd393;
a_sign0 = 4'd15; a_sign1 = 4'd11; a_sign2 = 4'd15; a_sign3 = 4'd2;
b_sign0 = 4'd9; b_sign1 = 4'd14; b_sign2 = 4'd1; b_sign3 = 4'd3;
@(posedge clk_i);
a_mant0 = 8'd193; a_mant1 = 8'd56; a_mant2 = 8'd90; a_mant3 = 8'd206;
b_mant0 = 8'd246; b_mant1 = 8'd112; b_mant2 = 8'd145; b_mant3 = 8'd160;
a_exp0 = 10'd276; a_exp1 = 10'd572; a_exp2 = 10'd242; a_exp3 = 10'd592;
b_exp0 = 10'd975; b_exp1 = 10'd56; b_exp2 = 10'd822; b_exp3 = 10'd780;
a_sign0 = 4'd15; a_sign1 = 4'd2; a_sign2 = 4'd16; a_sign3 = 4'd5;
b_sign0 = 4'd10; b_sign1 = 4'd10; b_sign2 = 4'd6; b_sign3 = 4'd15;
@(posedge clk_i);
a_mant0 = 8'd90; a_mant1 = 8'd3; a_mant2 = 8'd133; a_mant3 = 8'd3;
b_mant0 = 8'd95; b_mant1 = 8'd29; b_mant2 = 8'd87; b_mant3 = 8'd22;
a_exp0 = 10'd150; a_exp1 = 10'd632; a_exp2 = 10'd848; a_exp3 = 10'd584;
b_exp0 = 10'd760; b_exp1 = 10'd60; b_exp2 = 10'd963; b_exp3 = 10'd80;
a_sign0 = 4'd12; a_sign1 = 4'd1; a_sign2 = 4'd0; a_sign3 = 4'd6;
b_sign0 = 4'd3; b_sign1 = 4'd14; b_sign2 = 4'd3; b_sign3 = 4'd15;
@(posedge clk_i);
a_mant0 = 8'd147; a_mant1 = 8'd177; a_mant2 = 8'd45; a_mant3 = 8'd118;
b_mant0 = 8'd128; b_mant1 = 8'd254; b_mant2 = 8'd158; b_mant3 = 8'd128;
a_exp0 = 10'd950; a_exp1 = 10'd161; a_exp2 = 10'd378; a_exp3 = 10'd174;
b_exp0 = 10'd250; b_exp1 = 10'd513; b_exp2 = 10'd805; b_exp3 = 10'd509;
a_sign0 = 4'd3; a_sign1 = 4'd9; a_sign2 = 4'd13; a_sign3 = 4'd3;
b_sign0 = 4'd7; b_sign1 = 4'd5; b_sign2 = 4'd0; b_sign3 = 4'd2;
@(posedge clk_i);
a_mant0 = 8'd92; a_mant1 = 8'd226; a_mant2 = 8'd76; a_mant3 = 8'd43;
b_mant0 = 8'd106; b_mant1 = 8'd231; b_mant2 = 8'd217; b_mant3 = 8'd198;
a_exp0 = 10'd637; a_exp1 = 10'd690; a_exp2 = 10'd129; a_exp3 = 10'd640;
b_exp0 = 10'd550; b_exp1 = 10'd606; b_exp2 = 10'd351; b_exp3 = 10'd476;
a_sign0 = 4'd11; a_sign1 = 4'd3; a_sign2 = 4'd15; a_sign3 = 4'd2;
b_sign0 = 4'd6; b_sign1 = 4'd11; b_sign2 = 4'd1; b_sign3 = 4'd12;
@(posedge clk_i);
shared_exps0 = 8'd119;
shared_exps1 = 8'd137;
a_mant0 = 8'd130; a_mant1 = 8'd114; a_mant2 = 8'd211; a_mant3 = 8'd202;
b_mant0 = 8'd51; b_mant1 = 8'd88; b_mant2 = 8'd164; b_mant3 = 8'd255;
a_exp0 = 10'd118; a_exp1 = 10'd881; a_exp2 = 10'd411; a_exp3 = 10'd270;
b_exp0 = 10'd765; b_exp1 = 10'd465; b_exp2 = 10'd43; b_exp3 = 10'd13;
a_sign0 = 4'd7; a_sign1 = 4'd6; a_sign2 = 4'd13; a_sign3 = 4'd10;
b_sign0 = 4'd1; b_sign1 = 4'd2; b_sign2 = 4'd4; b_sign3 = 4'd3;
@(posedge clk_i);
a_mant0 = 8'd44; a_mant1 = 8'd52; a_mant2 = 8'd57; a_mant3 = 8'd19;
b_mant0 = 8'd42; b_mant1 = 8'd220; b_mant2 = 8'd47; b_mant3 = 8'd66;
a_exp0 = 10'd473; a_exp1 = 10'd609; a_exp2 = 10'd538; a_exp3 = 10'd302;
b_exp0 = 10'd767; b_exp1 = 10'd595; b_exp2 = 10'd327; b_exp3 = 10'd884;
a_sign0 = 4'd13; a_sign1 = 4'd10; a_sign2 = 4'd5; a_sign3 = 4'd0;
b_sign0 = 4'd15; b_sign1 = 4'd14; b_sign2 = 4'd15; b_sign3 = 4'd1;
@(posedge clk_i);
a_mant0 = 8'd128; a_mant1 = 8'd231; a_mant2 = 8'd195; a_mant3 = 8'd228;
b_mant0 = 8'd81; b_mant1 = 8'd191; b_mant2 = 8'd243; b_mant3 = 8'd125;
a_exp0 = 10'd441; a_exp1 = 10'd544; a_exp2 = 10'd141; a_exp3 = 10'd203;
b_exp0 = 10'd623; b_exp1 = 10'd453; b_exp2 = 10'd229; b_exp3 = 10'd931;
a_sign0 = 4'd16; a_sign1 = 4'd1; a_sign2 = 4'd5; a_sign3 = 4'd12;
b_sign0 = 4'd6; b_sign1 = 4'd5; b_sign2 = 4'd13; b_sign3 = 4'd5;
@(posedge clk_i);
a_mant0 = 8'd154; a_mant1 = 8'd130; a_mant2 = 8'd11; a_mant3 = 8'd141;
b_mant0 = 8'd72; b_mant1 = 8'd101; b_mant2 = 8'd54; b_mant3 = 8'd39;
a_exp0 = 10'd726; a_exp1 = 10'd849; a_exp2 = 10'd89; a_exp3 = 10'd152;
b_exp0 = 10'd505; b_exp1 = 10'd288; b_exp2 = 10'd190; b_exp3 = 10'd769;
a_sign0 = 4'd7; a_sign1 = 4'd10; a_sign2 = 4'd2; a_sign3 = 4'd13;
b_sign0 = 4'd2; b_sign1 = 4'd10; b_sign2 = 4'd16; b_sign3 = 4'd1;
@(posedge clk_i);
a_mant0 = 8'd147; a_mant1 = 8'd149; a_mant2 = 8'd211; a_mant3 = 8'd81;
b_mant0 = 8'd66; b_mant1 = 8'd113; b_mant2 = 8'd11; b_mant3 = 8'd182;
a_exp0 = 10'd502; a_exp1 = 10'd561; a_exp2 = 10'd747; a_exp3 = 10'd294;
b_exp0 = 10'd446; b_exp1 = 10'd860; b_exp2 = 10'd201; b_exp3 = 10'd519;
a_sign0 = 4'd9; a_sign1 = 4'd1; a_sign2 = 4'd11; a_sign3 = 4'd11;
b_sign0 = 4'd14; b_sign1 = 4'd2; b_sign2 = 4'd10; b_sign3 = 4'd3;
@(posedge clk_i);
a_mant0 = 8'd57; a_mant1 = 8'd214; a_mant2 = 8'd249; a_mant3 = 8'd162;
b_mant0 = 8'd221; b_mant1 = 8'd119; b_mant2 = 8'd63; b_mant3 = 8'd20;
a_exp0 = 10'd996; a_exp1 = 10'd160; a_exp2 = 10'd728; a_exp3 = 10'd1011;
b_exp0 = 10'd915; b_exp1 = 10'd64; b_exp2 = 10'd517; b_exp3 = 10'd908;
a_sign0 = 4'd0; a_sign1 = 4'd13; a_sign2 = 4'd4; a_sign3 = 4'd13;
b_sign0 = 4'd6; b_sign1 = 4'd1; b_sign2 = 4'd10; b_sign3 = 4'd11;
@(posedge clk_i);
a_mant0 = 8'd6; a_mant1 = 8'd126; a_mant2 = 8'd116; a_mant3 = 8'd30;
b_mant0 = 8'd227; b_mant1 = 8'd221; b_mant2 = 8'd112; b_mant3 = 8'd193;
a_exp0 = 10'd935; a_exp1 = 10'd550; a_exp2 = 10'd712; a_exp3 = 10'd22;
b_exp0 = 10'd269; b_exp1 = 10'd94; b_exp2 = 10'd396; b_exp3 = 10'd64;
a_sign0 = 4'd5; a_sign1 = 4'd13; a_sign2 = 4'd6; a_sign3 = 4'd5;
b_sign0 = 4'd16; b_sign1 = 4'd4; b_sign2 = 4'd0; b_sign3 = 4'd15;
@(posedge clk_i);
a_mant0 = 8'd56; a_mant1 = 8'd192; a_mant2 = 8'd95; a_mant3 = 8'd92;
b_mant0 = 8'd39; b_mant1 = 8'd96; b_mant2 = 8'd215; b_mant3 = 8'd245;
a_exp0 = 10'd853; a_exp1 = 10'd971; a_exp2 = 10'd253; a_exp3 = 10'd393;
b_exp0 = 10'd197; b_exp1 = 10'd411; b_exp2 = 10'd492; b_exp3 = 10'd663;
a_sign0 = 4'd0; a_sign1 = 4'd5; a_sign2 = 4'd12; a_sign3 = 4'd6;
b_sign0 = 4'd11; b_sign1 = 4'd0; b_sign2 = 4'd3; b_sign3 = 4'd13;
@(posedge clk_i);
shared_exps0 = 8'd107;
shared_exps1 = 8'd116;
a_mant0 = 8'd17; a_mant1 = 8'd169; a_mant2 = 8'd211; a_mant3 = 8'd27;
b_mant0 = 8'd12; b_mant1 = 8'd201; b_mant2 = 8'd138; b_mant3 = 8'd72;
a_exp0 = 10'd953; a_exp1 = 10'd110; a_exp2 = 10'd635; a_exp3 = 10'd195;
b_exp0 = 10'd961; b_exp1 = 10'd276; b_exp2 = 10'd847; b_exp3 = 10'd544;
a_sign0 = 4'd3; a_sign1 = 4'd4; a_sign2 = 4'd12; a_sign3 = 4'd0;
b_sign0 = 4'd5; b_sign1 = 4'd7; b_sign2 = 4'd9; b_sign3 = 4'd9;
@(posedge clk_i);
a_mant0 = 8'd46; a_mant1 = 8'd149; a_mant2 = 8'd36; a_mant3 = 8'd231;
b_mant0 = 8'd156; b_mant1 = 8'd208; b_mant2 = 8'd35; b_mant3 = 8'd202;
a_exp0 = 10'd775; a_exp1 = 10'd199; a_exp2 = 10'd496; a_exp3 = 10'd546;
b_exp0 = 10'd943; b_exp1 = 10'd968; b_exp2 = 10'd229; b_exp3 = 10'd808;
a_sign0 = 4'd15; a_sign1 = 4'd12; a_sign2 = 4'd9; a_sign3 = 4'd11;
b_sign0 = 4'd12; b_sign1 = 4'd4; b_sign2 = 4'd6; b_sign3 = 4'd12;
@(posedge clk_i);
a_mant0 = 8'd21; a_mant1 = 8'd0; a_mant2 = 8'd142; a_mant3 = 8'd204;
b_mant0 = 8'd85; b_mant1 = 8'd31; b_mant2 = 8'd212; b_mant3 = 8'd33;
a_exp0 = 10'd642; a_exp1 = 10'd704; a_exp2 = 10'd249; a_exp3 = 10'd395;
b_exp0 = 10'd510; b_exp1 = 10'd996; b_exp2 = 10'd480; b_exp3 = 10'd9;
a_sign0 = 4'd0; a_sign1 = 4'd10; a_sign2 = 4'd8; a_sign3 = 4'd15;
b_sign0 = 4'd8; b_sign1 = 4'd7; b_sign2 = 4'd11; b_sign3 = 4'd7;
@(posedge clk_i);
a_mant0 = 8'd1; a_mant1 = 8'd44; a_mant2 = 8'd71; a_mant3 = 8'd239;
b_mant0 = 8'd228; b_mant1 = 8'd73; b_mant2 = 8'd236; b_mant3 = 8'd212;
a_exp0 = 10'd1003; a_exp1 = 10'd355; a_exp2 = 10'd491; a_exp3 = 10'd883;
b_exp0 = 10'd50; b_exp1 = 10'd901; b_exp2 = 10'd758; b_exp3 = 10'd115;
a_sign0 = 4'd4; a_sign1 = 4'd7; a_sign2 = 4'd0; a_sign3 = 4'd7;
b_sign0 = 4'd12; b_sign1 = 4'd0; b_sign2 = 4'd9; b_sign3 = 4'd1;
@(posedge clk_i);
a_mant0 = 8'd44; a_mant1 = 8'd111; a_mant2 = 8'd165; a_mant3 = 8'd54;
b_mant0 = 8'd69; b_mant1 = 8'd173; b_mant2 = 8'd21; b_mant3 = 8'd58;
a_exp0 = 10'd113; a_exp1 = 10'd852; a_exp2 = 10'd475; a_exp3 = 10'd195;
b_exp0 = 10'd813; b_exp1 = 10'd669; b_exp2 = 10'd474; b_exp3 = 10'd717;
a_sign0 = 4'd7; a_sign1 = 4'd0; a_sign2 = 4'd3; a_sign3 = 4'd11;
b_sign0 = 4'd10; b_sign1 = 4'd10; b_sign2 = 4'd16; b_sign3 = 4'd5;
@(posedge clk_i);
a_mant0 = 8'd72; a_mant1 = 8'd65; a_mant2 = 8'd159; a_mant3 = 8'd155;
b_mant0 = 8'd132; b_mant1 = 8'd70; b_mant2 = 8'd185; b_mant3 = 8'd193;
a_exp0 = 10'd173; a_exp1 = 10'd356; a_exp2 = 10'd640; a_exp3 = 10'd676;
b_exp0 = 10'd406; b_exp1 = 10'd738; b_exp2 = 10'd394; b_exp3 = 10'd496;
a_sign0 = 4'd8; a_sign1 = 4'd5; a_sign2 = 4'd12; a_sign3 = 4'd7;
b_sign0 = 4'd1; b_sign1 = 4'd3; b_sign2 = 4'd11; b_sign3 = 4'd14;
@(posedge clk_i);
a_mant0 = 8'd105; a_mant1 = 8'd199; a_mant2 = 8'd133; a_mant3 = 8'd124;
b_mant0 = 8'd27; b_mant1 = 8'd142; b_mant2 = 8'd79; b_mant3 = 8'd231;
a_exp0 = 10'd540; a_exp1 = 10'd689; a_exp2 = 10'd507; a_exp3 = 10'd400;
b_exp0 = 10'd711; b_exp1 = 10'd395; b_exp2 = 10'd222; b_exp3 = 10'd842;
a_sign0 = 4'd2; a_sign1 = 4'd14; a_sign2 = 4'd1; a_sign3 = 4'd8;
b_sign0 = 4'd4; b_sign1 = 4'd4; b_sign2 = 4'd1; b_sign3 = 4'd15;
@(posedge clk_i);
a_mant0 = 8'd209; a_mant1 = 8'd86; a_mant2 = 8'd165; a_mant3 = 8'd137;
b_mant0 = 8'd232; b_mant1 = 8'd101; b_mant2 = 8'd105; b_mant3 = 8'd90;
a_exp0 = 10'd995; a_exp1 = 10'd781; a_exp2 = 10'd114; a_exp3 = 10'd999;
b_exp0 = 10'd882; b_exp1 = 10'd886; b_exp2 = 10'd249; b_exp3 = 10'd943;
a_sign0 = 4'd8; a_sign1 = 4'd1; a_sign2 = 4'd5; a_sign3 = 4'd6;
b_sign0 = 4'd4; b_sign1 = 4'd13; b_sign2 = 4'd0; b_sign3 = 4'd6;
@(posedge clk_i);
shared_exps0 = 8'd107;
shared_exps1 = 8'd128;
rstn = 0;
@(posedge clk_i);
rstn = 1;
a_mant0 = 8'd219; a_mant1 = 8'd13; a_mant2 = 8'd196; a_mant3 = 8'd218;
b_mant0 = 8'd75; b_mant1 = 8'd86; b_mant2 = 8'd136; b_mant3 = 8'd191;
a_exp0 = 10'd797; a_exp1 = 10'd734; a_exp2 = 10'd554; a_exp3 = 10'd882;
b_exp0 = 10'd370; b_exp1 = 10'd270; b_exp2 = 10'd190; b_exp3 = 10'd280;
a_sign0 = 4'd3; a_sign1 = 4'd9; a_sign2 = 4'd11; a_sign3 = 4'd14;
b_sign0 = 4'd15; b_sign1 = 4'd11; b_sign2 = 4'd15; b_sign3 = 4'd1;
@(posedge clk_i);
a_mant0 = 8'd103; a_mant1 = 8'd228; a_mant2 = 8'd199; a_mant3 = 8'd202;
b_mant0 = 8'd173; b_mant1 = 8'd18; b_mant2 = 8'd90; b_mant3 = 8'd136;
a_exp0 = 10'd890; a_exp1 = 10'd50; a_exp2 = 10'd864; a_exp3 = 10'd181;
b_exp0 = 10'd516; b_exp1 = 10'd414; b_exp2 = 10'd154; b_exp3 = 10'd641;
a_sign0 = 4'd3; a_sign1 = 4'd16; a_sign2 = 4'd9; a_sign3 = 4'd12;
b_sign0 = 4'd14; b_sign1 = 4'd2; b_sign2 = 4'd12; b_sign3 = 4'd6;
@(posedge clk_i);
a_mant0 = 8'd70; a_mant1 = 8'd129; a_mant2 = 8'd176; a_mant3 = 8'd21;
b_mant0 = 8'd42; b_mant1 = 8'd255; b_mant2 = 8'd80; b_mant3 = 8'd13;
a_exp0 = 10'd407; a_exp1 = 10'd97; a_exp2 = 10'd538; a_exp3 = 10'd631;
b_exp0 = 10'd538; b_exp1 = 10'd258; b_exp2 = 10'd531; b_exp3 = 10'd849;
a_sign0 = 4'd10; a_sign1 = 4'd8; a_sign2 = 4'd0; a_sign3 = 4'd1;
b_sign0 = 4'd5; b_sign1 = 4'd12; b_sign2 = 4'd15; b_sign3 = 4'd15;
@(posedge clk_i);
a_mant0 = 8'd18; a_mant1 = 8'd27; a_mant2 = 8'd83; a_mant3 = 8'd19;
b_mant0 = 8'd109; b_mant1 = 8'd56; b_mant2 = 8'd225; b_mant3 = 8'd39;
a_exp0 = 10'd289; a_exp1 = 10'd752; a_exp2 = 10'd806; a_exp3 = 10'd564;
b_exp0 = 10'd489; b_exp1 = 10'd414; b_exp2 = 10'd715; b_exp3 = 10'd108;
a_sign0 = 4'd10; a_sign1 = 4'd15; a_sign2 = 4'd16; a_sign3 = 4'd1;
b_sign0 = 4'd8; b_sign1 = 4'd16; b_sign2 = 4'd7; b_sign3 = 4'd5;
@(posedge clk_i);
a_mant0 = 8'd38; a_mant1 = 8'd115; a_mant2 = 8'd230; a_mant3 = 8'd58;
b_mant0 = 8'd193; b_mant1 = 8'd70; b_mant2 = 8'd67; b_mant3 = 8'd164;
a_exp0 = 10'd274; a_exp1 = 10'd835; a_exp2 = 10'd781; a_exp3 = 10'd742;
b_exp0 = 10'd871; b_exp1 = 10'd496; b_exp2 = 10'd871; b_exp3 = 10'd553;
a_sign0 = 4'd15; a_sign1 = 4'd8; a_sign2 = 4'd3; a_sign3 = 4'd7;
b_sign0 = 4'd3; b_sign1 = 4'd12; b_sign2 = 4'd6; b_sign3 = 4'd11;
@(posedge clk_i);
a_mant0 = 8'd71; a_mant1 = 8'd148; a_mant2 = 8'd180; a_mant3 = 8'd86;
b_mant0 = 8'd239; b_mant1 = 8'd24; b_mant2 = 8'd232; b_mant3 = 8'd84;
a_exp0 = 10'd956; a_exp1 = 10'd368; a_exp2 = 10'd158; a_exp3 = 10'd25;
b_exp0 = 10'd808; b_exp1 = 10'd803; b_exp2 = 10'd893; b_exp3 = 10'd894;
a_sign0 = 4'd3; a_sign1 = 4'd2; a_sign2 = 4'd15; a_sign3 = 4'd16;
b_sign0 = 4'd0; b_sign1 = 4'd15; b_sign2 = 4'd12; b_sign3 = 4'd0;
@(posedge clk_i);
a_mant0 = 8'd117; a_mant1 = 8'd17; a_mant2 = 8'd43; a_mant3 = 8'd4;
b_mant0 = 8'd62; b_mant1 = 8'd88; b_mant2 = 8'd132; b_mant3 = 8'd18;
a_exp0 = 10'd446; a_exp1 = 10'd164; a_exp2 = 10'd663; a_exp3 = 10'd913;
b_exp0 = 10'd941; b_exp1 = 10'd129; b_exp2 = 10'd173; b_exp3 = 10'd202;
a_sign0 = 4'd11; a_sign1 = 4'd5; a_sign2 = 4'd0; a_sign3 = 4'd13;
b_sign0 = 4'd6; b_sign1 = 4'd2; b_sign2 = 4'd12; b_sign3 = 4'd4;
@(posedge clk_i);
shared_exps0 = 8'd157;
shared_exps1 = 8'd128;
a_mant0 = 8'd176; a_mant1 = 8'd124; a_mant2 = 8'd81; a_mant3 = 8'd107;
b_mant0 = 8'd171; b_mant1 = 8'd212; b_mant2 = 8'd14; b_mant3 = 8'd209;
a_exp0 = 10'd251; a_exp1 = 10'd776; a_exp2 = 10'd527; a_exp3 = 10'd900;
b_exp0 = 10'd917; b_exp1 = 10'd722; b_exp2 = 10'd996; b_exp3 = 10'd80;
a_sign0 = 4'd16; a_sign1 = 4'd3; a_sign2 = 4'd6; a_sign3 = 4'd10;
b_sign0 = 4'd16; b_sign1 = 4'd6; b_sign2 = 4'd10; b_sign3 = 4'd3;
@(posedge clk_i);
a_mant0 = 8'd59; a_mant1 = 8'd100; a_mant2 = 8'd110; a_mant3 = 8'd247;
b_mant0 = 8'd201; b_mant1 = 8'd138; b_mant2 = 8'd109; b_mant3 = 8'd28;
a_exp0 = 10'd417; a_exp1 = 10'd946; a_exp2 = 10'd498; a_exp3 = 10'd524;
b_exp0 = 10'd558; b_exp1 = 10'd877; b_exp2 = 10'd94; b_exp3 = 10'd213;
a_sign0 = 4'd7; a_sign1 = 4'd15; a_sign2 = 4'd9; a_sign3 = 4'd8;
b_sign0 = 4'd15; b_sign1 = 4'd2; b_sign2 = 4'd12; b_sign3 = 4'd16;
@(posedge clk_i);
a_mant0 = 8'd227; a_mant1 = 8'd153; a_mant2 = 8'd195; a_mant3 = 8'd228;
b_mant0 = 8'd231; b_mant1 = 8'd220; b_mant2 = 8'd168; b_mant3 = 8'd114;
a_exp0 = 10'd760; a_exp1 = 10'd622; a_exp2 = 10'd249; a_exp3 = 10'd992;
b_exp0 = 10'd330; b_exp1 = 10'd509; b_exp2 = 10'd165; b_exp3 = 10'd656;
a_sign0 = 4'd5; a_sign1 = 4'd9; a_sign2 = 4'd0; a_sign3 = 4'd3;
b_sign0 = 4'd3; b_sign1 = 4'd1; b_sign2 = 4'd4; b_sign3 = 4'd0;
@(posedge clk_i);
a_mant0 = 8'd150; a_mant1 = 8'd41; a_mant2 = 8'd108; a_mant3 = 8'd181;
b_mant0 = 8'd130; b_mant1 = 8'd85; b_mant2 = 8'd181; b_mant3 = 8'd131;
a_exp0 = 10'd249; a_exp1 = 10'd463; a_exp2 = 10'd174; a_exp3 = 10'd676;
b_exp0 = 10'd840; b_exp1 = 10'd428; b_exp2 = 10'd725; b_exp3 = 10'd852;
a_sign0 = 4'd9; a_sign1 = 4'd9; a_sign2 = 4'd16; a_sign3 = 4'd9;
b_sign0 = 4'd9; b_sign1 = 4'd1; b_sign2 = 4'd11; b_sign3 = 4'd10;
@(posedge clk_i);
a_mant0 = 8'd22; a_mant1 = 8'd174; a_mant2 = 8'd90; a_mant3 = 8'd79;
b_mant0 = 8'd42; b_mant1 = 8'd3; b_mant2 = 8'd151; b_mant3 = 8'd133;
a_exp0 = 10'd140; a_exp1 = 10'd498; a_exp2 = 10'd156; a_exp3 = 10'd363;
b_exp0 = 10'd887; b_exp1 = 10'd666; b_exp2 = 10'd903; b_exp3 = 10'd513;
a_sign0 = 4'd2; a_sign1 = 4'd3; a_sign2 = 4'd3; a_sign3 = 4'd16;
b_sign0 = 4'd4; b_sign1 = 4'd7; b_sign2 = 4'd13; b_sign3 = 4'd7;
@(posedge clk_i);
a_mant0 = 8'd32; a_mant1 = 8'd159; a_mant2 = 8'd218; a_mant3 = 8'd163;
b_mant0 = 8'd141; b_mant1 = 8'd112; b_mant2 = 8'd84; b_mant3 = 8'd233;
a_exp0 = 10'd927; a_exp1 = 10'd498; a_exp2 = 10'd173; a_exp3 = 10'd427;
b_exp0 = 10'd181; b_exp1 = 10'd474; b_exp2 = 10'd936; b_exp3 = 10'd265;
a_sign0 = 4'd9; a_sign1 = 4'd0; a_sign2 = 4'd15; a_sign3 = 4'd16;
b_sign0 = 4'd3; b_sign1 = 4'd10; b_sign2 = 4'd7; b_sign3 = 4'd3;
@(posedge clk_i);
a_mant0 = 8'd22; a_mant1 = 8'd19; a_mant2 = 8'd167; a_mant3 = 8'd233;
b_mant0 = 8'd43; b_mant1 = 8'd9; b_mant2 = 8'd241; b_mant3 = 8'd180;
a_exp0 = 10'd220; a_exp1 = 10'd461; a_exp2 = 10'd950; a_exp3 = 10'd477;
b_exp0 = 10'd767; b_exp1 = 10'd48; b_exp2 = 10'd432; b_exp3 = 10'd413;
a_sign0 = 4'd2; a_sign1 = 4'd2; a_sign2 = 4'd15; a_sign3 = 4'd8;
b_sign0 = 4'd11; b_sign1 = 4'd9; b_sign2 = 4'd4; b_sign3 = 4'd11;
@(posedge clk_i);
a_mant0 = 8'd87; a_mant1 = 8'd27; a_mant2 = 8'd157; a_mant3 = 8'd6;
b_mant0 = 8'd79; b_mant1 = 8'd134; b_mant2 = 8'd120; b_mant3 = 8'd191;
a_exp0 = 10'd483; a_exp1 = 10'd906; a_exp2 = 10'd336; a_exp3 = 10'd923;
b_exp0 = 10'd414; b_exp1 = 10'd85; b_exp2 = 10'd402; b_exp3 = 10'd695;
a_sign0 = 4'd1; a_sign1 = 4'd10; a_sign2 = 4'd6; a_sign3 = 4'd14;
b_sign0 = 4'd13; b_sign1 = 4'd11; b_sign2 = 4'd9; b_sign3 = 4'd7;
@(posedge clk_i);
shared_exps0 = 8'd130;
shared_exps1 = 8'd114;
a_mant0 = 8'd65; a_mant1 = 8'd36; a_mant2 = 8'd247; a_mant3 = 8'd25;
b_mant0 = 8'd1; b_mant1 = 8'd242; b_mant2 = 8'd143; b_mant3 = 8'd129;
a_exp0 = 10'd573; a_exp1 = 10'd854; a_exp2 = 10'd290; a_exp3 = 10'd528;
b_exp0 = 10'd113; b_exp1 = 10'd141; b_exp2 = 10'd718; b_exp3 = 10'd764;
a_sign0 = 4'd15; a_sign1 = 4'd12; a_sign2 = 4'd11; a_sign3 = 4'd4;
b_sign0 = 4'd9; b_sign1 = 4'd8; b_sign2 = 4'd13; b_sign3 = 4'd12;
@(posedge clk_i);
a_mant0 = 8'd27; a_mant1 = 8'd165; a_mant2 = 8'd80; a_mant3 = 8'd5;
b_mant0 = 8'd155; b_mant1 = 8'd19; b_mant2 = 8'd200; b_mant3 = 8'd174;
a_exp0 = 10'd393; a_exp1 = 10'd123; a_exp2 = 10'd19; a_exp3 = 10'd836;
b_exp0 = 10'd322; b_exp1 = 10'd256; b_exp2 = 10'd367; b_exp3 = 10'd922;
a_sign0 = 4'd8; a_sign1 = 4'd9; a_sign2 = 4'd14; a_sign3 = 4'd0;
b_sign0 = 4'd10; b_sign1 = 4'd14; b_sign2 = 4'd3; b_sign3 = 4'd12;
@(posedge clk_i);
a_mant0 = 8'd50; a_mant1 = 8'd61; a_mant2 = 8'd59; a_mant3 = 8'd252;
b_mant0 = 8'd90; b_mant1 = 8'd191; b_mant2 = 8'd143; b_mant3 = 8'd18;
a_exp0 = 10'd225; a_exp1 = 10'd79; a_exp2 = 10'd583; a_exp3 = 10'd175;
b_exp0 = 10'd94; b_exp1 = 10'd496; b_exp2 = 10'd1008; b_exp3 = 10'd1005;
a_sign0 = 4'd16; a_sign1 = 4'd6; a_sign2 = 4'd1; a_sign3 = 4'd11;
b_sign0 = 4'd16; b_sign1 = 4'd14; b_sign2 = 4'd1; b_sign3 = 4'd15;
@(posedge clk_i);
a_mant0 = 8'd17; a_mant1 = 8'd163; a_mant2 = 8'd251; a_mant3 = 8'd39;
b_mant0 = 8'd178; b_mant1 = 8'd38; b_mant2 = 8'd213; b_mant3 = 8'd254;
a_exp0 = 10'd799; a_exp1 = 10'd959; a_exp2 = 10'd556; a_exp3 = 10'd402;
b_exp0 = 10'd93; b_exp1 = 10'd103; b_exp2 = 10'd132; b_exp3 = 10'd539;
a_sign0 = 4'd1; a_sign1 = 4'd10; a_sign2 = 4'd8; a_sign3 = 4'd2;
b_sign0 = 4'd9; b_sign1 = 4'd9; b_sign2 = 4'd3; b_sign3 = 4'd2;
@(posedge clk_i);
a_mant0 = 8'd168; a_mant1 = 8'd43; a_mant2 = 8'd80; a_mant3 = 8'd224;
b_mant0 = 8'd25; b_mant1 = 8'd92; b_mant2 = 8'd114; b_mant3 = 8'd27;
a_exp0 = 10'd809; a_exp1 = 10'd697; a_exp2 = 10'd91; a_exp3 = 10'd167;
b_exp0 = 10'd859; b_exp1 = 10'd192; b_exp2 = 10'd15; b_exp3 = 10'd257;
a_sign0 = 4'd9; a_sign1 = 4'd5; a_sign2 = 4'd7; a_sign3 = 4'd7;
b_sign0 = 4'd11; b_sign1 = 4'd9; b_sign2 = 4'd6; b_sign3 = 4'd4;
@(posedge clk_i);
a_mant0 = 8'd73; a_mant1 = 8'd3; a_mant2 = 8'd214; a_mant3 = 8'd68;
b_mant0 = 8'd52; b_mant1 = 8'd176; b_mant2 = 8'd94; b_mant3 = 8'd12;
a_exp0 = 10'd935; a_exp1 = 10'd400; a_exp2 = 10'd768; a_exp3 = 10'd892;
b_exp0 = 10'd971; b_exp1 = 10'd297; b_exp2 = 10'd819; b_exp3 = 10'd416;
a_sign0 = 4'd7; a_sign1 = 4'd16; a_sign2 = 4'd13; a_sign3 = 4'd3;
b_sign0 = 4'd1; b_sign1 = 4'd10; b_sign2 = 4'd1; b_sign3 = 4'd16;
@(posedge clk_i);
a_mant0 = 8'd243; a_mant1 = 8'd218; a_mant2 = 8'd143; a_mant3 = 8'd14;
b_mant0 = 8'd116; b_mant1 = 8'd117; b_mant2 = 8'd123; b_mant3 = 8'd158;
a_exp0 = 10'd671; a_exp1 = 10'd754; a_exp2 = 10'd298; a_exp3 = 10'd752;
b_exp0 = 10'd27; b_exp1 = 10'd493; b_exp2 = 10'd238; b_exp3 = 10'd147;
a_sign0 = 4'd15; a_sign1 = 4'd0; a_sign2 = 4'd7; a_sign3 = 4'd8;
b_sign0 = 4'd10; b_sign1 = 4'd9; b_sign2 = 4'd1; b_sign3 = 4'd2;
@(posedge clk_i);
a_mant0 = 8'd218; a_mant1 = 8'd26; a_mant2 = 8'd76; a_mant3 = 8'd195;
b_mant0 = 8'd43; b_mant1 = 8'd70; b_mant2 = 8'd235; b_mant3 = 8'd208;
a_exp0 = 10'd336; a_exp1 = 10'd199; a_exp2 = 10'd1014; a_exp3 = 10'd902;
b_exp0 = 10'd396; b_exp1 = 10'd162; b_exp2 = 10'd248; b_exp3 = 10'd484;
a_sign0 = 4'd13; a_sign1 = 4'd7; a_sign2 = 4'd14; a_sign3 = 4'd14;
b_sign0 = 4'd1; b_sign1 = 4'd7; b_sign2 = 4'd4; b_sign3 = 4'd15;
@(posedge clk_i);
shared_exps0 = 8'd146;
shared_exps1 = 8'd125;
a_mant0 = 8'd102; a_mant1 = 8'd253; a_mant2 = 8'd237; a_mant3 = 8'd69;
b_mant0 = 8'd85; b_mant1 = 8'd148; b_mant2 = 8'd84; b_mant3 = 8'd181;
a_exp0 = 10'd323; a_exp1 = 10'd345; a_exp2 = 10'd611; a_exp3 = 10'd905;
b_exp0 = 10'd29; b_exp1 = 10'd986; b_exp2 = 10'd282; b_exp3 = 10'd294;
a_sign0 = 4'd6; a_sign1 = 4'd7; a_sign2 = 4'd16; a_sign3 = 4'd11;
b_sign0 = 4'd6; b_sign1 = 4'd1; b_sign2 = 4'd9; b_sign3 = 4'd5;
@(posedge clk_i);
a_mant0 = 8'd153; a_mant1 = 8'd97; a_mant2 = 8'd220; a_mant3 = 8'd62;
b_mant0 = 8'd65; b_mant1 = 8'd59; b_mant2 = 8'd147; b_mant3 = 8'd97;
a_exp0 = 10'd946; a_exp1 = 10'd568; a_exp2 = 10'd385; a_exp3 = 10'd636;
b_exp0 = 10'd345; b_exp1 = 10'd475; b_exp2 = 10'd248; b_exp3 = 10'd724;
a_sign0 = 4'd11; a_sign1 = 4'd7; a_sign2 = 4'd8; a_sign3 = 4'd6;
b_sign0 = 4'd6; b_sign1 = 4'd6; b_sign2 = 4'd10; b_sign3 = 4'd5;
@(posedge clk_i);
a_mant0 = 8'd164; a_mant1 = 8'd12; a_mant2 = 8'd181; a_mant3 = 8'd65;
b_mant0 = 8'd47; b_mant1 = 8'd93; b_mant2 = 8'd120; b_mant3 = 8'd90;
a_exp0 = 10'd787; a_exp1 = 10'd497; a_exp2 = 10'd275; a_exp3 = 10'd146;
b_exp0 = 10'd330; b_exp1 = 10'd955; b_exp2 = 10'd268; b_exp3 = 10'd402;
a_sign0 = 4'd11; a_sign1 = 4'd14; a_sign2 = 4'd12; a_sign3 = 4'd7;
b_sign0 = 4'd2; b_sign1 = 4'd4; b_sign2 = 4'd16; b_sign3 = 4'd13;
@(posedge clk_i);
a_mant0 = 8'd67; a_mant1 = 8'd239; a_mant2 = 8'd246; a_mant3 = 8'd0;
b_mant0 = 8'd163; b_mant1 = 8'd106; b_mant2 = 8'd236; b_mant3 = 8'd149;
a_exp0 = 10'd644; a_exp1 = 10'd210; a_exp2 = 10'd794; a_exp3 = 10'd871;
b_exp0 = 10'd12; b_exp1 = 10'd651; b_exp2 = 10'd583; b_exp3 = 10'd692;
a_sign0 = 4'd5; a_sign1 = 4'd1; a_sign2 = 4'd12; a_sign3 = 4'd12;
b_sign0 = 4'd7; b_sign1 = 4'd0; b_sign2 = 4'd5; b_sign3 = 4'd6;
@(posedge clk_i);
a_mant0 = 8'd30; a_mant1 = 8'd137; a_mant2 = 8'd69; a_mant3 = 8'd89;
b_mant0 = 8'd200; b_mant1 = 8'd52; b_mant2 = 8'd87; b_mant3 = 8'd148;
a_exp0 = 10'd338; a_exp1 = 10'd412; a_exp2 = 10'd898; a_exp3 = 10'd1016;
b_exp0 = 10'd827; b_exp1 = 10'd593; b_exp2 = 10'd624; b_exp3 = 10'd913;
a_sign0 = 4'd14; a_sign1 = 4'd15; a_sign2 = 4'd9; a_sign3 = 4'd1;
b_sign0 = 4'd12; b_sign1 = 4'd12; b_sign2 = 4'd1; b_sign3 = 4'd1;
@(posedge clk_i);
a_mant0 = 8'd87; a_mant1 = 8'd77; a_mant2 = 8'd157; a_mant3 = 8'd197;
b_mant0 = 8'd218; b_mant1 = 8'd55; b_mant2 = 8'd117; b_mant3 = 8'd20;
a_exp0 = 10'd99; a_exp1 = 10'd477; a_exp2 = 10'd982; a_exp3 = 10'd91;
b_exp0 = 10'd740; b_exp1 = 10'd552; b_exp2 = 10'd473; b_exp3 = 10'd669;
a_sign0 = 4'd0; a_sign1 = 4'd4; a_sign2 = 4'd3; a_sign3 = 4'd5;
b_sign0 = 4'd1; b_sign1 = 4'd13; b_sign2 = 4'd15; b_sign3 = 4'd0;
@(posedge clk_i);
a_mant0 = 8'd230; a_mant1 = 8'd45; a_mant2 = 8'd165; a_mant3 = 8'd58;
b_mant0 = 8'd22; b_mant1 = 8'd73; b_mant2 = 8'd10; b_mant3 = 8'd17;
a_exp0 = 10'd939; a_exp1 = 10'd458; a_exp2 = 10'd63; a_exp3 = 10'd255;
b_exp0 = 10'd430; b_exp1 = 10'd56; b_exp2 = 10'd902; b_exp3 = 10'd670;
a_sign0 = 4'd7; a_sign1 = 4'd9; a_sign2 = 4'd9; a_sign3 = 4'd12;
b_sign0 = 4'd10; b_sign1 = 4'd16; b_sign2 = 4'd12; b_sign3 = 4'd13;
@(posedge clk_i);
a_mant0 = 8'd227; a_mant1 = 8'd11; a_mant2 = 8'd192; a_mant3 = 8'd187;
b_mant0 = 8'd81; b_mant1 = 8'd154; b_mant2 = 8'd231; b_mant3 = 8'd28;
a_exp0 = 10'd759; a_exp1 = 10'd203; a_exp2 = 10'd337; a_exp3 = 10'd937;
b_exp0 = 10'd199; b_exp1 = 10'd157; b_exp2 = 10'd1020; b_exp3 = 10'd507;
a_sign0 = 4'd0; a_sign1 = 4'd12; a_sign2 = 4'd16; a_sign3 = 4'd2;
b_sign0 = 4'd5; b_sign1 = 4'd3; b_sign2 = 4'd7; b_sign3 = 4'd2;
@(posedge clk_i);
shared_exps0 = 8'd120;
shared_exps1 = 8'd153;
rstn = 0;
@(posedge clk_i);
rstn = 1;
a_mant0 = 8'd197; a_mant1 = 8'd130; a_mant2 = 8'd209; a_mant3 = 8'd56;
b_mant0 = 8'd80; b_mant1 = 8'd79; b_mant2 = 8'd81; b_mant3 = 8'd112;
a_exp0 = 10'd1021; a_exp1 = 10'd909; a_exp2 = 10'd39; a_exp3 = 10'd392;
b_exp0 = 10'd838; b_exp1 = 10'd41; b_exp2 = 10'd230; b_exp3 = 10'd444;
a_sign0 = 4'd13; a_sign1 = 4'd6; a_sign2 = 4'd15; a_sign3 = 4'd9;
b_sign0 = 4'd5; b_sign1 = 4'd0; b_sign2 = 4'd6; b_sign3 = 4'd12;
@(posedge clk_i);
a_mant0 = 8'd11; a_mant1 = 8'd158; a_mant2 = 8'd196; a_mant3 = 8'd237;
b_mant0 = 8'd30; b_mant1 = 8'd155; b_mant2 = 8'd28; b_mant3 = 8'd170;
a_exp0 = 10'd96; a_exp1 = 10'd56; a_exp2 = 10'd958; a_exp3 = 10'd503;
b_exp0 = 10'd257; b_exp1 = 10'd214; b_exp2 = 10'd103; b_exp3 = 10'd891;
a_sign0 = 4'd4; a_sign1 = 4'd14; a_sign2 = 4'd6; a_sign3 = 4'd8;
b_sign0 = 4'd6; b_sign1 = 4'd11; b_sign2 = 4'd10; b_sign3 = 4'd4;
@(posedge clk_i);
a_mant0 = 8'd237; a_mant1 = 8'd39; a_mant2 = 8'd19; a_mant3 = 8'd67;
b_mant0 = 8'd38; b_mant1 = 8'd85; b_mant2 = 8'd53; b_mant3 = 8'd33;
a_exp0 = 10'd922; a_exp1 = 10'd147; a_exp2 = 10'd1001; a_exp3 = 10'd761;
b_exp0 = 10'd679; b_exp1 = 10'd90; b_exp2 = 10'd344; b_exp3 = 10'd89;
a_sign0 = 4'd0; a_sign1 = 4'd1; a_sign2 = 4'd10; a_sign3 = 4'd0;
b_sign0 = 4'd1; b_sign1 = 4'd3; b_sign2 = 4'd12; b_sign3 = 4'd0;
@(posedge clk_i);
a_mant0 = 8'd144; a_mant1 = 8'd147; a_mant2 = 8'd175; a_mant3 = 8'd212;
b_mant0 = 8'd91; b_mant1 = 8'd22; b_mant2 = 8'd108; b_mant3 = 8'd83;
a_exp0 = 10'd314; a_exp1 = 10'd296; a_exp2 = 10'd665; a_exp3 = 10'd828;
b_exp0 = 10'd776; b_exp1 = 10'd561; b_exp2 = 10'd925; b_exp3 = 10'd319;
a_sign0 = 4'd15; a_sign1 = 4'd1; a_sign2 = 4'd11; a_sign3 = 4'd12;
b_sign0 = 4'd12; b_sign1 = 4'd10; b_sign2 = 4'd2; b_sign3 = 4'd0;
@(posedge clk_i);
a_mant0 = 8'd9; a_mant1 = 8'd210; a_mant2 = 8'd155; a_mant3 = 8'd157;
b_mant0 = 8'd69; b_mant1 = 8'd251; b_mant2 = 8'd243; b_mant3 = 8'd171;
a_exp0 = 10'd754; a_exp1 = 10'd990; a_exp2 = 10'd855; a_exp3 = 10'd559;
b_exp0 = 10'd534; b_exp1 = 10'd32; b_exp2 = 10'd803; b_exp3 = 10'd778;
a_sign0 = 4'd1; a_sign1 = 4'd13; a_sign2 = 4'd1; a_sign3 = 4'd15;
b_sign0 = 4'd7; b_sign1 = 4'd0; b_sign2 = 4'd6; b_sign3 = 4'd3;
@(posedge clk_i);
a_mant0 = 8'd234; a_mant1 = 8'd22; a_mant2 = 8'd52; a_mant3 = 8'd165;
b_mant0 = 8'd151; b_mant1 = 8'd205; b_mant2 = 8'd205; b_mant3 = 8'd28;
a_exp0 = 10'd941; a_exp1 = 10'd719; a_exp2 = 10'd272; a_exp3 = 10'd50;
b_exp0 = 10'd441; b_exp1 = 10'd207; b_exp2 = 10'd476; b_exp3 = 10'd752;
a_sign0 = 4'd0; a_sign1 = 4'd10; a_sign2 = 4'd4; a_sign3 = 4'd15;
b_sign0 = 4'd11; b_sign1 = 4'd1; b_sign2 = 4'd2; b_sign3 = 4'd4;
@(posedge clk_i);
a_mant0 = 8'd132; a_mant1 = 8'd109; a_mant2 = 8'd100; a_mant3 = 8'd23;
b_mant0 = 8'd224; b_mant1 = 8'd29; b_mant2 = 8'd57; b_mant3 = 8'd137;
a_exp0 = 10'd592; a_exp1 = 10'd892; a_exp2 = 10'd429; a_exp3 = 10'd977;
b_exp0 = 10'd543; b_exp1 = 10'd292; b_exp2 = 10'd123; b_exp3 = 10'd867;
a_sign0 = 4'd12; a_sign1 = 4'd16; a_sign2 = 4'd1; a_sign3 = 4'd4;
b_sign0 = 4'd5; b_sign1 = 4'd12; b_sign2 = 4'd4; b_sign3 = 4'd7;
@(posedge clk_i);
shared_exps0 = 8'd124;
shared_exps1 = 8'd123;
a_mant0 = 8'd148; a_mant1 = 8'd10; a_mant2 = 8'd146; a_mant3 = 8'd9;
b_mant0 = 8'd199; b_mant1 = 8'd193; b_mant2 = 8'd47; b_mant3 = 8'd221;
a_exp0 = 10'd24; a_exp1 = 10'd122; a_exp2 = 10'd145; a_exp3 = 10'd979;
b_exp0 = 10'd145; b_exp1 = 10'd579; b_exp2 = 10'd43; b_exp3 = 10'd198;
a_sign0 = 4'd10; a_sign1 = 4'd13; a_sign2 = 4'd16; a_sign3 = 4'd16;
b_sign0 = 4'd0; b_sign1 = 4'd1; b_sign2 = 4'd7; b_sign3 = 4'd5;
@(posedge clk_i);
a_mant0 = 8'd1; a_mant1 = 8'd67; a_mant2 = 8'd189; a_mant3 = 8'd47;
b_mant0 = 8'd60; b_mant1 = 8'd127; b_mant2 = 8'd104; b_mant3 = 8'd241;
a_exp0 = 10'd770; a_exp1 = 10'd318; a_exp2 = 10'd402; a_exp3 = 10'd92;
b_exp0 = 10'd10; b_exp1 = 10'd412; b_exp2 = 10'd227; b_exp3 = 10'd663;
a_sign0 = 4'd8; a_sign1 = 4'd2; a_sign2 = 4'd14; a_sign3 = 4'd3;
b_sign0 = 4'd10; b_sign1 = 4'd12; b_sign2 = 4'd16; b_sign3 = 4'd10;
@(posedge clk_i);
a_mant0 = 8'd125; a_mant1 = 8'd150; a_mant2 = 8'd27; a_mant3 = 8'd134;
b_mant0 = 8'd221; b_mant1 = 8'd198; b_mant2 = 8'd183; b_mant3 = 8'd124;
a_exp0 = 10'd394; a_exp1 = 10'd530; a_exp2 = 10'd921; a_exp3 = 10'd166;
b_exp0 = 10'd82; b_exp1 = 10'd635; b_exp2 = 10'd857; b_exp3 = 10'd993;
a_sign0 = 4'd2; a_sign1 = 4'd10; a_sign2 = 4'd2; a_sign3 = 4'd4;
b_sign0 = 4'd4; b_sign1 = 4'd16; b_sign2 = 4'd8; b_sign3 = 4'd13;
@(posedge clk_i);
a_mant0 = 8'd129; a_mant1 = 8'd100; a_mant2 = 8'd69; a_mant3 = 8'd139;
b_mant0 = 8'd206; b_mant1 = 8'd112; b_mant2 = 8'd94; b_mant3 = 8'd30;
a_exp0 = 10'd69; a_exp1 = 10'd949; a_exp2 = 10'd811; a_exp3 = 10'd402;
b_exp0 = 10'd456; b_exp1 = 10'd597; b_exp2 = 10'd708; b_exp3 = 10'd114;
a_sign0 = 4'd8; a_sign1 = 4'd6; a_sign2 = 4'd1; a_sign3 = 4'd11;
b_sign0 = 4'd1; b_sign1 = 4'd4; b_sign2 = 4'd13; b_sign3 = 4'd15;
@(posedge clk_i);
a_mant0 = 8'd59; a_mant1 = 8'd127; a_mant2 = 8'd57; a_mant3 = 8'd235;
b_mant0 = 8'd127; b_mant1 = 8'd208; b_mant2 = 8'd237; b_mant3 = 8'd15;
a_exp0 = 10'd554; a_exp1 = 10'd145; a_exp2 = 10'd624; a_exp3 = 10'd848;
b_exp0 = 10'd84; b_exp1 = 10'd395; b_exp2 = 10'd206; b_exp3 = 10'd253;
a_sign0 = 4'd1; a_sign1 = 4'd5; a_sign2 = 4'd1; a_sign3 = 4'd11;
b_sign0 = 4'd9; b_sign1 = 4'd16; b_sign2 = 4'd5; b_sign3 = 4'd2;
@(posedge clk_i);
a_mant0 = 8'd173; a_mant1 = 8'd124; a_mant2 = 8'd137; a_mant3 = 8'd179;
b_mant0 = 8'd84; b_mant1 = 8'd228; b_mant2 = 8'd157; b_mant3 = 8'd83;
a_exp0 = 10'd276; a_exp1 = 10'd465; a_exp2 = 10'd107; a_exp3 = 10'd896;
b_exp0 = 10'd125; b_exp1 = 10'd666; b_exp2 = 10'd477; b_exp3 = 10'd746;
a_sign0 = 4'd2; a_sign1 = 4'd12; a_sign2 = 4'd7; a_sign3 = 4'd14;
b_sign0 = 4'd7; b_sign1 = 4'd3; b_sign2 = 4'd16; b_sign3 = 4'd0;
@(posedge clk_i);
a_mant0 = 8'd245; a_mant1 = 8'd231; a_mant2 = 8'd169; a_mant3 = 8'd64;
b_mant0 = 8'd175; b_mant1 = 8'd116; b_mant2 = 8'd2; b_mant3 = 8'd205;
a_exp0 = 10'd636; a_exp1 = 10'd701; a_exp2 = 10'd979; a_exp3 = 10'd344;
b_exp0 = 10'd277; b_exp1 = 10'd472; b_exp2 = 10'd279; b_exp3 = 10'd860;
a_sign0 = 4'd6; a_sign1 = 4'd7; a_sign2 = 4'd6; a_sign3 = 4'd2;
b_sign0 = 4'd9; b_sign1 = 4'd4; b_sign2 = 4'd0; b_sign3 = 4'd12;
@(posedge clk_i);
a_mant0 = 8'd228; a_mant1 = 8'd74; a_mant2 = 8'd47; a_mant3 = 8'd203;
b_mant0 = 8'd218; b_mant1 = 8'd188; b_mant2 = 8'd181; b_mant3 = 8'd254;
a_exp0 = 10'd100; a_exp1 = 10'd414; a_exp2 = 10'd812; a_exp3 = 10'd922;
b_exp0 = 10'd914; b_exp1 = 10'd695; b_exp2 = 10'd481; b_exp3 = 10'd320;
a_sign0 = 4'd3; a_sign1 = 4'd8; a_sign2 = 4'd7; a_sign3 = 4'd10;
b_sign0 = 4'd14; b_sign1 = 4'd12; b_sign2 = 4'd13; b_sign3 = 4'd8;
@(posedge clk_i);
shared_exps0 = 8'd115;
shared_exps1 = 8'd126;
a_mant0 = 8'd133; a_mant1 = 8'd93; a_mant2 = 8'd110; a_mant3 = 8'd108;
b_mant0 = 8'd166; b_mant1 = 8'd141; b_mant2 = 8'd154; b_mant3 = 8'd9;
a_exp0 = 10'd522; a_exp1 = 10'd667; a_exp2 = 10'd615; a_exp3 = 10'd736;
b_exp0 = 10'd316; b_exp1 = 10'd462; b_exp2 = 10'd20; b_exp3 = 10'd729;
a_sign0 = 4'd6; a_sign1 = 4'd15; a_sign2 = 4'd1; a_sign3 = 4'd10;
b_sign0 = 4'd13; b_sign1 = 4'd15; b_sign2 = 4'd4; b_sign3 = 4'd14;
@(posedge clk_i);
a_mant0 = 8'd114; a_mant1 = 8'd1; a_mant2 = 8'd40; a_mant3 = 8'd177;
b_mant0 = 8'd238; b_mant1 = 8'd212; b_mant2 = 8'd157; b_mant3 = 8'd104;
a_exp0 = 10'd907; a_exp1 = 10'd9; a_exp2 = 10'd65; a_exp3 = 10'd794;
b_exp0 = 10'd39; b_exp1 = 10'd6; b_exp2 = 10'd546; b_exp3 = 10'd665;
a_sign0 = 4'd2; a_sign1 = 4'd6; a_sign2 = 4'd15; a_sign3 = 4'd1;
b_sign0 = 4'd5; b_sign1 = 4'd15; b_sign2 = 4'd3; b_sign3 = 4'd0;
@(posedge clk_i);
a_mant0 = 8'd247; a_mant1 = 8'd16; a_mant2 = 8'd116; a_mant3 = 8'd147;
b_mant0 = 8'd82; b_mant1 = 8'd232; b_mant2 = 8'd48; b_mant3 = 8'd101;
a_exp0 = 10'd412; a_exp1 = 10'd868; a_exp2 = 10'd402; a_exp3 = 10'd305;
b_exp0 = 10'd370; b_exp1 = 10'd461; b_exp2 = 10'd367; b_exp3 = 10'd421;
a_sign0 = 4'd4; a_sign1 = 4'd5; a_sign2 = 4'd5; a_sign3 = 4'd13;
b_sign0 = 4'd8; b_sign1 = 4'd14; b_sign2 = 4'd12; b_sign3 = 4'd5;
@(posedge clk_i);
a_mant0 = 8'd109; a_mant1 = 8'd206; a_mant2 = 8'd42; a_mant3 = 8'd219;
b_mant0 = 8'd65; b_mant1 = 8'd83; b_mant2 = 8'd100; b_mant3 = 8'd85;
a_exp0 = 10'd355; a_exp1 = 10'd584; a_exp2 = 10'd652; a_exp3 = 10'd935;
b_exp0 = 10'd1020; b_exp1 = 10'd447; b_exp2 = 10'd841; b_exp3 = 10'd363;
a_sign0 = 4'd6; a_sign1 = 4'd8; a_sign2 = 4'd16; a_sign3 = 4'd16;
b_sign0 = 4'd16; b_sign1 = 4'd4; b_sign2 = 4'd3; b_sign3 = 4'd5;
@(posedge clk_i);
a_mant0 = 8'd115; a_mant1 = 8'd52; a_mant2 = 8'd147; a_mant3 = 8'd129;
b_mant0 = 8'd237; b_mant1 = 8'd152; b_mant2 = 8'd66; b_mant3 = 8'd155;
a_exp0 = 10'd294; a_exp1 = 10'd920; a_exp2 = 10'd445; a_exp3 = 10'd935;
b_exp0 = 10'd251; b_exp1 = 10'd171; b_exp2 = 10'd161; b_exp3 = 10'd200;
a_sign0 = 4'd11; a_sign1 = 4'd8; a_sign2 = 4'd8; a_sign3 = 4'd8;
b_sign0 = 4'd13; b_sign1 = 4'd12; b_sign2 = 4'd15; b_sign3 = 4'd16;
@(posedge clk_i);
a_mant0 = 8'd13; a_mant1 = 8'd42; a_mant2 = 8'd238; a_mant3 = 8'd96;
b_mant0 = 8'd245; b_mant1 = 8'd132; b_mant2 = 8'd181; b_mant3 = 8'd30;
a_exp0 = 10'd120; a_exp1 = 10'd682; a_exp2 = 10'd908; a_exp3 = 10'd20;
b_exp0 = 10'd897; b_exp1 = 10'd334; b_exp2 = 10'd395; b_exp3 = 10'd413;
a_sign0 = 4'd5; a_sign1 = 4'd6; a_sign2 = 4'd12; a_sign3 = 4'd4;
b_sign0 = 4'd11; b_sign1 = 4'd8; b_sign2 = 4'd7; b_sign3 = 4'd6;
@(posedge clk_i);
a_mant0 = 8'd123; a_mant1 = 8'd150; a_mant2 = 8'd149; a_mant3 = 8'd22;
b_mant0 = 8'd13; b_mant1 = 8'd245; b_mant2 = 8'd73; b_mant3 = 8'd41;
a_exp0 = 10'd562; a_exp1 = 10'd928; a_exp2 = 10'd198; a_exp3 = 10'd266;
b_exp0 = 10'd826; b_exp1 = 10'd479; b_exp2 = 10'd812; b_exp3 = 10'd784;
a_sign0 = 4'd9; a_sign1 = 4'd4; a_sign2 = 4'd6; a_sign3 = 4'd11;
b_sign0 = 4'd3; b_sign1 = 4'd13; b_sign2 = 4'd4; b_sign3 = 4'd16;
@(posedge clk_i);
a_mant0 = 8'd150; a_mant1 = 8'd178; a_mant2 = 8'd139; a_mant3 = 8'd118;
b_mant0 = 8'd20; b_mant1 = 8'd194; b_mant2 = 8'd69; b_mant3 = 8'd16;
a_exp0 = 10'd912; a_exp1 = 10'd844; a_exp2 = 10'd58; a_exp3 = 10'd109;
b_exp0 = 10'd538; b_exp1 = 10'd565; b_exp2 = 10'd221; b_exp3 = 10'd628;
a_sign0 = 4'd14; a_sign1 = 4'd12; a_sign2 = 4'd14; a_sign3 = 4'd16;
b_sign0 = 4'd0; b_sign1 = 4'd16; b_sign2 = 4'd3; b_sign3 = 4'd0;
@(posedge clk_i);
shared_exps0 = 8'd122;
shared_exps1 = 8'd137;
a_mant0 = 8'd205; a_mant1 = 8'd127; a_mant2 = 8'd41; a_mant3 = 8'd18;
b_mant0 = 8'd137; b_mant1 = 8'd84; b_mant2 = 8'd137; b_mant3 = 8'd222;
a_exp0 = 10'd958; a_exp1 = 10'd100; a_exp2 = 10'd757; a_exp3 = 10'd487;
b_exp0 = 10'd992; b_exp1 = 10'd1011; b_exp2 = 10'd258; b_exp3 = 10'd533;
a_sign0 = 4'd3; a_sign1 = 4'd4; a_sign2 = 4'd15; a_sign3 = 4'd0;
b_sign0 = 4'd8; b_sign1 = 4'd14; b_sign2 = 4'd6; b_sign3 = 4'd3;
@(posedge clk_i);
a_mant0 = 8'd93; a_mant1 = 8'd226; a_mant2 = 8'd1; a_mant3 = 8'd250;
b_mant0 = 8'd132; b_mant1 = 8'd159; b_mant2 = 8'd183; b_mant3 = 8'd211;
a_exp0 = 10'd403; a_exp1 = 10'd248; a_exp2 = 10'd614; a_exp3 = 10'd251;
b_exp0 = 10'd296; b_exp1 = 10'd274; b_exp2 = 10'd855; b_exp3 = 10'd853;
a_sign0 = 4'd11; a_sign1 = 4'd4; a_sign2 = 4'd15; a_sign3 = 4'd12;
b_sign0 = 4'd16; b_sign1 = 4'd1; b_sign2 = 4'd15; b_sign3 = 4'd16;
@(posedge clk_i);
a_mant0 = 8'd215; a_mant1 = 8'd150; a_mant2 = 8'd249; a_mant3 = 8'd72;
b_mant0 = 8'd16; b_mant1 = 8'd51; b_mant2 = 8'd68; b_mant3 = 8'd136;
a_exp0 = 10'd753; a_exp1 = 10'd705; a_exp2 = 10'd410; a_exp3 = 10'd900;
b_exp0 = 10'd817; b_exp1 = 10'd736; b_exp2 = 10'd620; b_exp3 = 10'd818;
a_sign0 = 4'd14; a_sign1 = 4'd13; a_sign2 = 4'd6; a_sign3 = 4'd15;
b_sign0 = 4'd8; b_sign1 = 4'd6; b_sign2 = 4'd12; b_sign3 = 4'd13;
@(posedge clk_i);
a_mant0 = 8'd192; a_mant1 = 8'd142; a_mant2 = 8'd181; a_mant3 = 8'd98;
b_mant0 = 8'd21; b_mant1 = 8'd111; b_mant2 = 8'd19; b_mant3 = 8'd122;
a_exp0 = 10'd965; a_exp1 = 10'd938; a_exp2 = 10'd814; a_exp3 = 10'd249;
b_exp0 = 10'd752; b_exp1 = 10'd581; b_exp2 = 10'd172; b_exp3 = 10'd908;
a_sign0 = 4'd12; a_sign1 = 4'd7; a_sign2 = 4'd8; a_sign3 = 4'd2;
b_sign0 = 4'd4; b_sign1 = 4'd4; b_sign2 = 4'd13; b_sign3 = 4'd4;
@(posedge clk_i);
a_mant0 = 8'd111; a_mant1 = 8'd252; a_mant2 = 8'd141; a_mant3 = 8'd170;
b_mant0 = 8'd50; b_mant1 = 8'd68; b_mant2 = 8'd219; b_mant3 = 8'd111;
a_exp0 = 10'd636; a_exp1 = 10'd575; a_exp2 = 10'd950; a_exp3 = 10'd94;
b_exp0 = 10'd920; b_exp1 = 10'd257; b_exp2 = 10'd1; b_exp3 = 10'd589;
a_sign0 = 4'd13; a_sign1 = 4'd3; a_sign2 = 4'd3; a_sign3 = 4'd15;
b_sign0 = 4'd15; b_sign1 = 4'd3; b_sign2 = 4'd1; b_sign3 = 4'd4;
@(posedge clk_i);
a_mant0 = 8'd206; a_mant1 = 8'd225; a_mant2 = 8'd81; a_mant3 = 8'd134;
b_mant0 = 8'd68; b_mant1 = 8'd252; b_mant2 = 8'd222; b_mant3 = 8'd46;
a_exp0 = 10'd672; a_exp1 = 10'd587; a_exp2 = 10'd953; a_exp3 = 10'd339;
b_exp0 = 10'd31; b_exp1 = 10'd717; b_exp2 = 10'd784; b_exp3 = 10'd532;
a_sign0 = 4'd9; a_sign1 = 4'd2; a_sign2 = 4'd10; a_sign3 = 4'd8;
b_sign0 = 4'd0; b_sign1 = 4'd3; b_sign2 = 4'd8; b_sign3 = 4'd7;
@(posedge clk_i);
a_mant0 = 8'd118; a_mant1 = 8'd45; a_mant2 = 8'd15; a_mant3 = 8'd110;
b_mant0 = 8'd222; b_mant1 = 8'd60; b_mant2 = 8'd10; b_mant3 = 8'd173;
a_exp0 = 10'd352; a_exp1 = 10'd414; a_exp2 = 10'd382; a_exp3 = 10'd125;
b_exp0 = 10'd735; b_exp1 = 10'd277; b_exp2 = 10'd1003; b_exp3 = 10'd643;
a_sign0 = 4'd16; a_sign1 = 4'd16; a_sign2 = 4'd2; a_sign3 = 4'd5;
b_sign0 = 4'd5; b_sign1 = 4'd11; b_sign2 = 4'd5; b_sign3 = 4'd6;
@(posedge clk_i);
a_mant0 = 8'd94; a_mant1 = 8'd181; a_mant2 = 8'd222; a_mant3 = 8'd133;
b_mant0 = 8'd131; b_mant1 = 8'd215; b_mant2 = 8'd197; b_mant3 = 8'd142;
a_exp0 = 10'd745; a_exp1 = 10'd1008; a_exp2 = 10'd634; a_exp3 = 10'd414;
b_exp0 = 10'd353; b_exp1 = 10'd402; b_exp2 = 10'd218; b_exp3 = 10'd808;
a_sign0 = 4'd10; a_sign1 = 4'd6; a_sign2 = 4'd16; a_sign3 = 4'd3;
b_sign0 = 4'd11; b_sign1 = 4'd2; b_sign2 = 4'd5; b_sign3 = 4'd0;
@(posedge clk_i);
shared_exps0 = 8'd100;
shared_exps1 = 8'd126;
rstn = 0;
@(posedge clk_i);
rstn = 1;
a_mant0 = 8'd220; a_mant1 = 8'd88; a_mant2 = 8'd105; a_mant3 = 8'd224;
b_mant0 = 8'd4; b_mant1 = 8'd120; b_mant2 = 8'd238; b_mant3 = 8'd7;
a_exp0 = 10'd271; a_exp1 = 10'd444; a_exp2 = 10'd682; a_exp3 = 10'd636;
b_exp0 = 10'd814; b_exp1 = 10'd659; b_exp2 = 10'd819; b_exp3 = 10'd798;
a_sign0 = 4'd7; a_sign1 = 4'd7; a_sign2 = 4'd5; a_sign3 = 4'd7;
b_sign0 = 4'd3; b_sign1 = 4'd7; b_sign2 = 4'd15; b_sign3 = 4'd12;
@(posedge clk_i);
a_mant0 = 8'd207; a_mant1 = 8'd69; a_mant2 = 8'd252; a_mant3 = 8'd126;
b_mant0 = 8'd242; b_mant1 = 8'd6; b_mant2 = 8'd92; b_mant3 = 8'd247;
a_exp0 = 10'd310; a_exp1 = 10'd986; a_exp2 = 10'd232; a_exp3 = 10'd433;
b_exp0 = 10'd94; b_exp1 = 10'd409; b_exp2 = 10'd847; b_exp3 = 10'd525;
a_sign0 = 4'd2; a_sign1 = 4'd3; a_sign2 = 4'd16; a_sign3 = 4'd16;
b_sign0 = 4'd15; b_sign1 = 4'd7; b_sign2 = 4'd14; b_sign3 = 4'd10;
@(posedge clk_i);
a_mant0 = 8'd188; a_mant1 = 8'd55; a_mant2 = 8'd225; a_mant3 = 8'd140;
b_mant0 = 8'd240; b_mant1 = 8'd213; b_mant2 = 8'd115; b_mant3 = 8'd37;
a_exp0 = 10'd798; a_exp1 = 10'd818; a_exp2 = 10'd299; a_exp3 = 10'd532;
b_exp0 = 10'd402; b_exp1 = 10'd993; b_exp2 = 10'd329; b_exp3 = 10'd884;
a_sign0 = 4'd16; a_sign1 = 4'd11; a_sign2 = 4'd7; a_sign3 = 4'd14;
b_sign0 = 4'd5; b_sign1 = 4'd14; b_sign2 = 4'd10; b_sign3 = 4'd10;
@(posedge clk_i);
a_mant0 = 8'd3; a_mant1 = 8'd116; a_mant2 = 8'd123; a_mant3 = 8'd149;
b_mant0 = 8'd75; b_mant1 = 8'd44; b_mant2 = 8'd63; b_mant3 = 8'd139;
a_exp0 = 10'd856; a_exp1 = 10'd500; a_exp2 = 10'd553; a_exp3 = 10'd553;
b_exp0 = 10'd392; b_exp1 = 10'd252; b_exp2 = 10'd154; b_exp3 = 10'd815;
a_sign0 = 4'd13; a_sign1 = 4'd5; a_sign2 = 4'd8; a_sign3 = 4'd3;
b_sign0 = 4'd8; b_sign1 = 4'd15; b_sign2 = 4'd13; b_sign3 = 4'd3;
@(posedge clk_i);
a_mant0 = 8'd41; a_mant1 = 8'd28; a_mant2 = 8'd1; a_mant3 = 8'd99;
b_mant0 = 8'd199; b_mant1 = 8'd230; b_mant2 = 8'd201; b_mant3 = 8'd85;
a_exp0 = 10'd434; a_exp1 = 10'd84; a_exp2 = 10'd561; a_exp3 = 10'd590;
b_exp0 = 10'd41; b_exp1 = 10'd793; b_exp2 = 10'd23; b_exp3 = 10'd856;
a_sign0 = 4'd0; a_sign1 = 4'd13; a_sign2 = 4'd1; a_sign3 = 4'd15;
b_sign0 = 4'd16; b_sign1 = 4'd6; b_sign2 = 4'd8; b_sign3 = 4'd12;
@(posedge clk_i);
a_mant0 = 8'd240; a_mant1 = 8'd249; a_mant2 = 8'd201; a_mant3 = 8'd87;
b_mant0 = 8'd197; b_mant1 = 8'd206; b_mant2 = 8'd146; b_mant3 = 8'd78;
a_exp0 = 10'd447; a_exp1 = 10'd821; a_exp2 = 10'd931; a_exp3 = 10'd834;
b_exp0 = 10'd726; b_exp1 = 10'd773; b_exp2 = 10'd235; b_exp3 = 10'd135;
a_sign0 = 4'd16; a_sign1 = 4'd6; a_sign2 = 4'd3; a_sign3 = 4'd14;
b_sign0 = 4'd9; b_sign1 = 4'd2; b_sign2 = 4'd0; b_sign3 = 4'd15;
@(posedge clk_i);
a_mant0 = 8'd50; a_mant1 = 8'd249; a_mant2 = 8'd247; a_mant3 = 8'd149;
b_mant0 = 8'd61; b_mant1 = 8'd54; b_mant2 = 8'd176; b_mant3 = 8'd152;
a_exp0 = 10'd997; a_exp1 = 10'd203; a_exp2 = 10'd8; a_exp3 = 10'd358;
b_exp0 = 10'd533; b_exp1 = 10'd868; b_exp2 = 10'd106; b_exp3 = 10'd656;
a_sign0 = 4'd5; a_sign1 = 4'd13; a_sign2 = 4'd3; a_sign3 = 4'd3;
b_sign0 = 4'd3; b_sign1 = 4'd14; b_sign2 = 4'd6; b_sign3 = 4'd13;
@(posedge clk_i);
shared_exps0 = 8'd114;
shared_exps1 = 8'd141;
a_mant0 = 8'd213; a_mant1 = 8'd215; a_mant2 = 8'd128; a_mant3 = 8'd129;
b_mant0 = 8'd240; b_mant1 = 8'd33; b_mant2 = 8'd138; b_mant3 = 8'd1;
a_exp0 = 10'd795; a_exp1 = 10'd238; a_exp2 = 10'd784; a_exp3 = 10'd393;
b_exp0 = 10'd108; b_exp1 = 10'd179; b_exp2 = 10'd963; b_exp3 = 10'd922;
a_sign0 = 4'd3; a_sign1 = 4'd8; a_sign2 = 4'd2; a_sign3 = 4'd11;
b_sign0 = 4'd13; b_sign1 = 4'd0; b_sign2 = 4'd8; b_sign3 = 4'd6;
@(posedge clk_i);
a_mant0 = 8'd196; a_mant1 = 8'd54; a_mant2 = 8'd190; a_mant3 = 8'd215;
b_mant0 = 8'd95; b_mant1 = 8'd241; b_mant2 = 8'd156; b_mant3 = 8'd221;
a_exp0 = 10'd277; a_exp1 = 10'd814; a_exp2 = 10'd58; a_exp3 = 10'd433;
b_exp0 = 10'd927; b_exp1 = 10'd673; b_exp2 = 10'd998; b_exp3 = 10'd223;
a_sign0 = 4'd14; a_sign1 = 4'd12; a_sign2 = 4'd8; a_sign3 = 4'd1;
b_sign0 = 4'd15; b_sign1 = 4'd14; b_sign2 = 4'd15; b_sign3 = 4'd11;
@(posedge clk_i);
a_mant0 = 8'd59; a_mant1 = 8'd160; a_mant2 = 8'd6; a_mant3 = 8'd1;
b_mant0 = 8'd207; b_mant1 = 8'd252; b_mant2 = 8'd190; b_mant3 = 8'd219;
a_exp0 = 10'd791; a_exp1 = 10'd744; a_exp2 = 10'd418; a_exp3 = 10'd966;
b_exp0 = 10'd128; b_exp1 = 10'd243; b_exp2 = 10'd944; b_exp3 = 10'd574;
a_sign0 = 4'd12; a_sign1 = 4'd6; a_sign2 = 4'd5; a_sign3 = 4'd6;
b_sign0 = 4'd9; b_sign1 = 4'd2; b_sign2 = 4'd12; b_sign3 = 4'd0;
@(posedge clk_i);
a_mant0 = 8'd65; a_mant1 = 8'd27; a_mant2 = 8'd51; a_mant3 = 8'd67;
b_mant0 = 8'd192; b_mant1 = 8'd170; b_mant2 = 8'd3; b_mant3 = 8'd47;
a_exp0 = 10'd303; a_exp1 = 10'd695; a_exp2 = 10'd53; a_exp3 = 10'd936;
b_exp0 = 10'd298; b_exp1 = 10'd554; b_exp2 = 10'd146; b_exp3 = 10'd717;
a_sign0 = 4'd16; a_sign1 = 4'd4; a_sign2 = 4'd2; a_sign3 = 4'd2;
b_sign0 = 4'd13; b_sign1 = 4'd5; b_sign2 = 4'd2; b_sign3 = 4'd11;
@(posedge clk_i);
a_mant0 = 8'd1; a_mant1 = 8'd186; a_mant2 = 8'd191; a_mant3 = 8'd107;
b_mant0 = 8'd2; b_mant1 = 8'd250; b_mant2 = 8'd19; b_mant3 = 8'd8;
a_exp0 = 10'd670; a_exp1 = 10'd475; a_exp2 = 10'd53; a_exp3 = 10'd836;
b_exp0 = 10'd650; b_exp1 = 10'd314; b_exp2 = 10'd374; b_exp3 = 10'd997;
a_sign0 = 4'd11; a_sign1 = 4'd14; a_sign2 = 4'd16; a_sign3 = 4'd15;
b_sign0 = 4'd5; b_sign1 = 4'd14; b_sign2 = 4'd2; b_sign3 = 4'd9;
@(posedge clk_i);
a_mant0 = 8'd254; a_mant1 = 8'd50; a_mant2 = 8'd116; a_mant3 = 8'd141;
b_mant0 = 8'd57; b_mant1 = 8'd134; b_mant2 = 8'd89; b_mant3 = 8'd103;
a_exp0 = 10'd238; a_exp1 = 10'd816; a_exp2 = 10'd414; a_exp3 = 10'd161;
b_exp0 = 10'd470; b_exp1 = 10'd701; b_exp2 = 10'd785; b_exp3 = 10'd238;
a_sign0 = 4'd11; a_sign1 = 4'd10; a_sign2 = 4'd6; a_sign3 = 4'd10;
b_sign0 = 4'd8; b_sign1 = 4'd12; b_sign2 = 4'd8; b_sign3 = 4'd1;
@(posedge clk_i);
a_mant0 = 8'd45; a_mant1 = 8'd76; a_mant2 = 8'd51; a_mant3 = 8'd208;
b_mant0 = 8'd216; b_mant1 = 8'd30; b_mant2 = 8'd15; b_mant3 = 8'd117;
a_exp0 = 10'd247; a_exp1 = 10'd775; a_exp2 = 10'd917; a_exp3 = 10'd875;
b_exp0 = 10'd169; b_exp1 = 10'd162; b_exp2 = 10'd204; b_exp3 = 10'd1023;
a_sign0 = 4'd8; a_sign1 = 4'd12; a_sign2 = 4'd1; a_sign3 = 4'd12;
b_sign0 = 4'd7; b_sign1 = 4'd15; b_sign2 = 4'd13; b_sign3 = 4'd10;
@(posedge clk_i);
a_mant0 = 8'd243; a_mant1 = 8'd207; a_mant2 = 8'd105; a_mant3 = 8'd141;
b_mant0 = 8'd0; b_mant1 = 8'd142; b_mant2 = 8'd98; b_mant3 = 8'd21;
a_exp0 = 10'd941; a_exp1 = 10'd585; a_exp2 = 10'd818; a_exp3 = 10'd319;
b_exp0 = 10'd914; b_exp1 = 10'd926; b_exp2 = 10'd600; b_exp3 = 10'd134;
a_sign0 = 4'd10; a_sign1 = 4'd2; a_sign2 = 4'd4; a_sign3 = 4'd14;
b_sign0 = 4'd2; b_sign1 = 4'd10; b_sign2 = 4'd1; b_sign3 = 4'd9;
@(posedge clk_i);
shared_exps0 = 8'd107;
shared_exps1 = 8'd131;
a_mant0 = 8'd150; a_mant1 = 8'd183; a_mant2 = 8'd186; a_mant3 = 8'd178;
b_mant0 = 8'd188; b_mant1 = 8'd80; b_mant2 = 8'd124; b_mant3 = 8'd34;
a_exp0 = 10'd351; a_exp1 = 10'd543; a_exp2 = 10'd494; a_exp3 = 10'd308;
b_exp0 = 10'd819; b_exp1 = 10'd719; b_exp2 = 10'd732; b_exp3 = 10'd896;
a_sign0 = 4'd2; a_sign1 = 4'd15; a_sign2 = 4'd11; a_sign3 = 4'd5;
b_sign0 = 4'd0; b_sign1 = 4'd6; b_sign2 = 4'd10; b_sign3 = 4'd3;
@(posedge clk_i);
a_mant0 = 8'd2; a_mant1 = 8'd96; a_mant2 = 8'd216; a_mant3 = 8'd133;
b_mant0 = 8'd254; b_mant1 = 8'd17; b_mant2 = 8'd145; b_mant3 = 8'd222;
a_exp0 = 10'd513; a_exp1 = 10'd330; a_exp2 = 10'd623; a_exp3 = 10'd794;
b_exp0 = 10'd909; b_exp1 = 10'd293; b_exp2 = 10'd273; b_exp3 = 10'd598;
a_sign0 = 4'd2; a_sign1 = 4'd4; a_sign2 = 4'd4; a_sign3 = 4'd8;
b_sign0 = 4'd10; b_sign1 = 4'd5; b_sign2 = 4'd10; b_sign3 = 4'd9;
@(posedge clk_i);
a_mant0 = 8'd54; a_mant1 = 8'd85; a_mant2 = 8'd88; a_mant3 = 8'd112;
b_mant0 = 8'd102; b_mant1 = 8'd128; b_mant2 = 8'd207; b_mant3 = 8'd219;
a_exp0 = 10'd354; a_exp1 = 10'd846; a_exp2 = 10'd425; a_exp3 = 10'd897;
b_exp0 = 10'd228; b_exp1 = 10'd616; b_exp2 = 10'd83; b_exp3 = 10'd649;
a_sign0 = 4'd13; a_sign1 = 4'd4; a_sign2 = 4'd0; a_sign3 = 4'd11;
b_sign0 = 4'd8; b_sign1 = 4'd15; b_sign2 = 4'd11; b_sign3 = 4'd8;
@(posedge clk_i);
a_mant0 = 8'd66; a_mant1 = 8'd51; a_mant2 = 8'd102; a_mant3 = 8'd184;
b_mant0 = 8'd110; b_mant1 = 8'd26; b_mant2 = 8'd201; b_mant3 = 8'd167;
a_exp0 = 10'd805; a_exp1 = 10'd775; a_exp2 = 10'd671; a_exp3 = 10'd864;
b_exp0 = 10'd73; b_exp1 = 10'd466; b_exp2 = 10'd597; b_exp3 = 10'd62;
a_sign0 = 4'd12; a_sign1 = 4'd16; a_sign2 = 4'd10; a_sign3 = 4'd1;
b_sign0 = 4'd15; b_sign1 = 4'd15; b_sign2 = 4'd13; b_sign3 = 4'd9;
@(posedge clk_i);
a_mant0 = 8'd111; a_mant1 = 8'd138; a_mant2 = 8'd135; a_mant3 = 8'd213;
b_mant0 = 8'd252; b_mant1 = 8'd200; b_mant2 = 8'd226; b_mant3 = 8'd230;
a_exp0 = 10'd923; a_exp1 = 10'd570; a_exp2 = 10'd133; a_exp3 = 10'd237;
b_exp0 = 10'd463; b_exp1 = 10'd745; b_exp2 = 10'd758; b_exp3 = 10'd686;
a_sign0 = 4'd2; a_sign1 = 4'd4; a_sign2 = 4'd11; a_sign3 = 4'd6;
b_sign0 = 4'd15; b_sign1 = 4'd5; b_sign2 = 4'd15; b_sign3 = 4'd4;
@(posedge clk_i);
a_mant0 = 8'd187; a_mant1 = 8'd50; a_mant2 = 8'd61; a_mant3 = 8'd13;
b_mant0 = 8'd227; b_mant1 = 8'd51; b_mant2 = 8'd0; b_mant3 = 8'd108;
a_exp0 = 10'd518; a_exp1 = 10'd311; a_exp2 = 10'd508; a_exp3 = 10'd792;
b_exp0 = 10'd196; b_exp1 = 10'd734; b_exp2 = 10'd552; b_exp3 = 10'd732;
a_sign0 = 4'd10; a_sign1 = 4'd7; a_sign2 = 4'd7; a_sign3 = 4'd16;
b_sign0 = 4'd12; b_sign1 = 4'd8; b_sign2 = 4'd15; b_sign3 = 4'd6;
@(posedge clk_i);
a_mant0 = 8'd222; a_mant1 = 8'd249; a_mant2 = 8'd81; a_mant3 = 8'd86;
b_mant0 = 8'd255; b_mant1 = 8'd124; b_mant2 = 8'd137; b_mant3 = 8'd192;
a_exp0 = 10'd416; a_exp1 = 10'd1015; a_exp2 = 10'd320; a_exp3 = 10'd760;
b_exp0 = 10'd344; b_exp1 = 10'd267; b_exp2 = 10'd482; b_exp3 = 10'd762;
a_sign0 = 4'd7; a_sign1 = 4'd5; a_sign2 = 4'd4; a_sign3 = 4'd12;
b_sign0 = 4'd0; b_sign1 = 4'd14; b_sign2 = 4'd11; b_sign3 = 4'd9;
@(posedge clk_i);
a_mant0 = 8'd78; a_mant1 = 8'd240; a_mant2 = 8'd152; a_mant3 = 8'd182;
b_mant0 = 8'd83; b_mant1 = 8'd18; b_mant2 = 8'd130; b_mant3 = 8'd2;
a_exp0 = 10'd324; a_exp1 = 10'd208; a_exp2 = 10'd344; a_exp3 = 10'd438;
b_exp0 = 10'd350; b_exp1 = 10'd325; b_exp2 = 10'd613; b_exp3 = 10'd921;
a_sign0 = 4'd6; a_sign1 = 4'd7; a_sign2 = 4'd4; a_sign3 = 4'd16;
b_sign0 = 4'd8; b_sign1 = 4'd7; b_sign2 = 4'd11; b_sign3 = 4'd4;
@(posedge clk_i);
shared_exps0 = 8'd142;
shared_exps1 = 8'd108;
a_mant0 = 8'd88; a_mant1 = 8'd36; a_mant2 = 8'd251; a_mant3 = 8'd60;
b_mant0 = 8'd231; b_mant1 = 8'd185; b_mant2 = 8'd224; b_mant3 = 8'd152;
a_exp0 = 10'd393; a_exp1 = 10'd26; a_exp2 = 10'd307; a_exp3 = 10'd724;
b_exp0 = 10'd672; b_exp1 = 10'd583; b_exp2 = 10'd335; b_exp3 = 10'd492;
a_sign0 = 4'd12; a_sign1 = 4'd1; a_sign2 = 4'd3; a_sign3 = 4'd1;
b_sign0 = 4'd1; b_sign1 = 4'd5; b_sign2 = 4'd10; b_sign3 = 4'd1;
@(posedge clk_i);
a_mant0 = 8'd113; a_mant1 = 8'd163; a_mant2 = 8'd172; a_mant3 = 8'd193;
b_mant0 = 8'd178; b_mant1 = 8'd205; b_mant2 = 8'd4; b_mant3 = 8'd215;
a_exp0 = 10'd494; a_exp1 = 10'd372; a_exp2 = 10'd273; a_exp3 = 10'd873;
b_exp0 = 10'd357; b_exp1 = 10'd1013; b_exp2 = 10'd800; b_exp3 = 10'd610;
a_sign0 = 4'd0; a_sign1 = 4'd11; a_sign2 = 4'd12; a_sign3 = 4'd6;
b_sign0 = 4'd12; b_sign1 = 4'd1; b_sign2 = 4'd12; b_sign3 = 4'd6;
@(posedge clk_i);
a_mant0 = 8'd45; a_mant1 = 8'd168; a_mant2 = 8'd58; a_mant3 = 8'd106;
b_mant0 = 8'd251; b_mant1 = 8'd195; b_mant2 = 8'd114; b_mant3 = 8'd111;
a_exp0 = 10'd250; a_exp1 = 10'd217; a_exp2 = 10'd216; a_exp3 = 10'd616;
b_exp0 = 10'd661; b_exp1 = 10'd1006; b_exp2 = 10'd387; b_exp3 = 10'd752;
a_sign0 = 4'd9; a_sign1 = 4'd7; a_sign2 = 4'd5; a_sign3 = 4'd5;
b_sign0 = 4'd10; b_sign1 = 4'd14; b_sign2 = 4'd0; b_sign3 = 4'd0;
@(posedge clk_i);
a_mant0 = 8'd40; a_mant1 = 8'd116; a_mant2 = 8'd56; a_mant3 = 8'd57;
b_mant0 = 8'd234; b_mant1 = 8'd129; b_mant2 = 8'd85; b_mant3 = 8'd31;
a_exp0 = 10'd310; a_exp1 = 10'd120; a_exp2 = 10'd16; a_exp3 = 10'd803;
b_exp0 = 10'd340; b_exp1 = 10'd230; b_exp2 = 10'd930; b_exp3 = 10'd183;
a_sign0 = 4'd8; a_sign1 = 4'd1; a_sign2 = 4'd7; a_sign3 = 4'd13;
b_sign0 = 4'd4; b_sign1 = 4'd7; b_sign2 = 4'd1; b_sign3 = 4'd13;
@(posedge clk_i);
a_mant0 = 8'd194; a_mant1 = 8'd51; a_mant2 = 8'd49; a_mant3 = 8'd121;
b_mant0 = 8'd27; b_mant1 = 8'd186; b_mant2 = 8'd34; b_mant3 = 8'd67;
a_exp0 = 10'd399; a_exp1 = 10'd954; a_exp2 = 10'd345; a_exp3 = 10'd189;
b_exp0 = 10'd385; b_exp1 = 10'd900; b_exp2 = 10'd684; b_exp3 = 10'd837;
a_sign0 = 4'd14; a_sign1 = 4'd14; a_sign2 = 4'd6; a_sign3 = 4'd14;
b_sign0 = 4'd13; b_sign1 = 4'd15; b_sign2 = 4'd0; b_sign3 = 4'd11;
@(posedge clk_i);
a_mant0 = 8'd32; a_mant1 = 8'd107; a_mant2 = 8'd44; a_mant3 = 8'd121;
b_mant0 = 8'd168; b_mant1 = 8'd55; b_mant2 = 8'd160; b_mant3 = 8'd85;
a_exp0 = 10'd362; a_exp1 = 10'd37; a_exp2 = 10'd619; a_exp3 = 10'd248;
b_exp0 = 10'd515; b_exp1 = 10'd490; b_exp2 = 10'd578; b_exp3 = 10'd305;
a_sign0 = 4'd15; a_sign1 = 4'd6; a_sign2 = 4'd3; a_sign3 = 4'd5;
b_sign0 = 4'd2; b_sign1 = 4'd16; b_sign2 = 4'd12; b_sign3 = 4'd9;
@(posedge clk_i);
a_mant0 = 8'd90; a_mant1 = 8'd89; a_mant2 = 8'd151; a_mant3 = 8'd58;
b_mant0 = 8'd135; b_mant1 = 8'd145; b_mant2 = 8'd113; b_mant3 = 8'd168;
a_exp0 = 10'd756; a_exp1 = 10'd678; a_exp2 = 10'd528; a_exp3 = 10'd469;
b_exp0 = 10'd38; b_exp1 = 10'd383; b_exp2 = 10'd795; b_exp3 = 10'd791;
a_sign0 = 4'd14; a_sign1 = 4'd4; a_sign2 = 4'd13; a_sign3 = 4'd3;
b_sign0 = 4'd4; b_sign1 = 4'd0; b_sign2 = 4'd12; b_sign3 = 4'd13;
@(posedge clk_i);
a_mant0 = 8'd64; a_mant1 = 8'd28; a_mant2 = 8'd54; a_mant3 = 8'd137;
b_mant0 = 8'd59; b_mant1 = 8'd135; b_mant2 = 8'd66; b_mant3 = 8'd76;
a_exp0 = 10'd847; a_exp1 = 10'd184; a_exp2 = 10'd257; a_exp3 = 10'd484;
b_exp0 = 10'd115; b_exp1 = 10'd169; b_exp2 = 10'd128; b_exp3 = 10'd301;
a_sign0 = 4'd13; a_sign1 = 4'd8; a_sign2 = 4'd7; a_sign3 = 4'd6;
b_sign0 = 4'd9; b_sign1 = 4'd15; b_sign2 = 4'd10; b_sign3 = 4'd12;
@(posedge clk_i);
shared_exps0 = 8'd156;
shared_exps1 = 8'd140;
rstn = 0;
@(posedge clk_i);
rstn = 1;
a_mant0 = 8'd163; a_mant1 = 8'd65; a_mant2 = 8'd35; a_mant3 = 8'd105;
b_mant0 = 8'd248; b_mant1 = 8'd196; b_mant2 = 8'd31; b_mant3 = 8'd252;
a_exp0 = 10'd583; a_exp1 = 10'd126; a_exp2 = 10'd268; a_exp3 = 10'd646;
b_exp0 = 10'd924; b_exp1 = 10'd321; b_exp2 = 10'd1004; b_exp3 = 10'd104;
a_sign0 = 4'd7; a_sign1 = 4'd16; a_sign2 = 4'd11; a_sign3 = 4'd9;
b_sign0 = 4'd3; b_sign1 = 4'd16; b_sign2 = 4'd4; b_sign3 = 4'd12;
@(posedge clk_i);
a_mant0 = 8'd82; a_mant1 = 8'd61; a_mant2 = 8'd222; a_mant3 = 8'd228;
b_mant0 = 8'd235; b_mant1 = 8'd103; b_mant2 = 8'd142; b_mant3 = 8'd61;
a_exp0 = 10'd614; a_exp1 = 10'd307; a_exp2 = 10'd306; a_exp3 = 10'd329;
b_exp0 = 10'd143; b_exp1 = 10'd741; b_exp2 = 10'd35; b_exp3 = 10'd667;
a_sign0 = 4'd1; a_sign1 = 4'd7; a_sign2 = 4'd1; a_sign3 = 4'd11;
b_sign0 = 4'd2; b_sign1 = 4'd15; b_sign2 = 4'd14; b_sign3 = 4'd16;
@(posedge clk_i);
a_mant0 = 8'd163; a_mant1 = 8'd62; a_mant2 = 8'd71; a_mant3 = 8'd194;
b_mant0 = 8'd46; b_mant1 = 8'd158; b_mant2 = 8'd175; b_mant3 = 8'd12;
a_exp0 = 10'd424; a_exp1 = 10'd715; a_exp2 = 10'd212; a_exp3 = 10'd138;
b_exp0 = 10'd389; b_exp1 = 10'd889; b_exp2 = 10'd584; b_exp3 = 10'd222;
a_sign0 = 4'd12; a_sign1 = 4'd9; a_sign2 = 4'd8; a_sign3 = 4'd15;
b_sign0 = 4'd8; b_sign1 = 4'd7; b_sign2 = 4'd13; b_sign3 = 4'd4;
@(posedge clk_i);
a_mant0 = 8'd117; a_mant1 = 8'd170; a_mant2 = 8'd207; a_mant3 = 8'd109;
b_mant0 = 8'd45; b_mant1 = 8'd2; b_mant2 = 8'd120; b_mant3 = 8'd76;
a_exp0 = 10'd930; a_exp1 = 10'd581; a_exp2 = 10'd855; a_exp3 = 10'd606;
b_exp0 = 10'd898; b_exp1 = 10'd254; b_exp2 = 10'd729; b_exp3 = 10'd781;
a_sign0 = 4'd8; a_sign1 = 4'd13; a_sign2 = 4'd9; a_sign3 = 4'd5;
b_sign0 = 4'd10; b_sign1 = 4'd4; b_sign2 = 4'd0; b_sign3 = 4'd11;
@(posedge clk_i);
a_mant0 = 8'd2; a_mant1 = 8'd136; a_mant2 = 8'd128; a_mant3 = 8'd210;
b_mant0 = 8'd90; b_mant1 = 8'd79; b_mant2 = 8'd165; b_mant3 = 8'd62;
a_exp0 = 10'd323; a_exp1 = 10'd848; a_exp2 = 10'd173; a_exp3 = 10'd271;
b_exp0 = 10'd663; b_exp1 = 10'd878; b_exp2 = 10'd28; b_exp3 = 10'd976;
a_sign0 = 4'd10; a_sign1 = 4'd13; a_sign2 = 4'd9; a_sign3 = 4'd5;
b_sign0 = 4'd7; b_sign1 = 4'd11; b_sign2 = 4'd3; b_sign3 = 4'd11;
@(posedge clk_i);
a_mant0 = 8'd144; a_mant1 = 8'd209; a_mant2 = 8'd66; a_mant3 = 8'd169;
b_mant0 = 8'd123; b_mant1 = 8'd222; b_mant2 = 8'd189; b_mant3 = 8'd98;
a_exp0 = 10'd903; a_exp1 = 10'd182; a_exp2 = 10'd511; a_exp3 = 10'd50;
b_exp0 = 10'd23; b_exp1 = 10'd258; b_exp2 = 10'd418; b_exp3 = 10'd402;
a_sign0 = 4'd11; a_sign1 = 4'd13; a_sign2 = 4'd8; a_sign3 = 4'd16;
b_sign0 = 4'd15; b_sign1 = 4'd11; b_sign2 = 4'd10; b_sign3 = 4'd3;
@(posedge clk_i);
a_mant0 = 8'd100; a_mant1 = 8'd108; a_mant2 = 8'd18; a_mant3 = 8'd5;
b_mant0 = 8'd177; b_mant1 = 8'd99; b_mant2 = 8'd174; b_mant3 = 8'd74;
a_exp0 = 10'd76; a_exp1 = 10'd572; a_exp2 = 10'd523; a_exp3 = 10'd319;
b_exp0 = 10'd487; b_exp1 = 10'd656; b_exp2 = 10'd172; b_exp3 = 10'd1021;
a_sign0 = 4'd2; a_sign1 = 4'd2; a_sign2 = 4'd6; a_sign3 = 4'd6;
b_sign0 = 4'd11; b_sign1 = 4'd8; b_sign2 = 4'd6; b_sign3 = 4'd6;
@(posedge clk_i);
shared_exps0 = 8'd145;
shared_exps1 = 8'd125;
a_mant0 = 8'd54; a_mant1 = 8'd151; a_mant2 = 8'd236; a_mant3 = 8'd248;
b_mant0 = 8'd68; b_mant1 = 8'd73; b_mant2 = 8'd200; b_mant3 = 8'd43;
a_exp0 = 10'd179; a_exp1 = 10'd356; a_exp2 = 10'd271; a_exp3 = 10'd377;
b_exp0 = 10'd88; b_exp1 = 10'd433; b_exp2 = 10'd264; b_exp3 = 10'd847;
a_sign0 = 4'd8; a_sign1 = 4'd14; a_sign2 = 4'd10; a_sign3 = 4'd13;
b_sign0 = 4'd15; b_sign1 = 4'd16; b_sign2 = 4'd11; b_sign3 = 4'd4;
@(posedge clk_i);
a_mant0 = 8'd58; a_mant1 = 8'd152; a_mant2 = 8'd181; a_mant3 = 8'd209;
b_mant0 = 8'd254; b_mant1 = 8'd149; b_mant2 = 8'd215; b_mant3 = 8'd33;
a_exp0 = 10'd249; a_exp1 = 10'd333; a_exp2 = 10'd146; a_exp3 = 10'd410;
b_exp0 = 10'd422; b_exp1 = 10'd538; b_exp2 = 10'd113; b_exp3 = 10'd181;
a_sign0 = 4'd12; a_sign1 = 4'd16; a_sign2 = 4'd11; a_sign3 = 4'd6;
b_sign0 = 4'd12; b_sign1 = 4'd0; b_sign2 = 4'd1; b_sign3 = 4'd1;
@(posedge clk_i);
a_mant0 = 8'd189; a_mant1 = 8'd177; a_mant2 = 8'd214; a_mant3 = 8'd92;
b_mant0 = 8'd111; b_mant1 = 8'd55; b_mant2 = 8'd2; b_mant3 = 8'd78;
a_exp0 = 10'd321; a_exp1 = 10'd612; a_exp2 = 10'd380; a_exp3 = 10'd764;
b_exp0 = 10'd618; b_exp1 = 10'd171; b_exp2 = 10'd333; b_exp3 = 10'd194;
a_sign0 = 4'd7; a_sign1 = 4'd12; a_sign2 = 4'd4; a_sign3 = 4'd14;
b_sign0 = 4'd10; b_sign1 = 4'd15; b_sign2 = 4'd0; b_sign3 = 4'd4;
@(posedge clk_i);
a_mant0 = 8'd61; a_mant1 = 8'd144; a_mant2 = 8'd195; a_mant3 = 8'd223;
b_mant0 = 8'd152; b_mant1 = 8'd225; b_mant2 = 8'd174; b_mant3 = 8'd211;
a_exp0 = 10'd687; a_exp1 = 10'd1021; a_exp2 = 10'd816; a_exp3 = 10'd234;
b_exp0 = 10'd710; b_exp1 = 10'd514; b_exp2 = 10'd186; b_exp3 = 10'd181;
a_sign0 = 4'd15; a_sign1 = 4'd1; a_sign2 = 4'd15; a_sign3 = 4'd5;
b_sign0 = 4'd8; b_sign1 = 4'd1; b_sign2 = 4'd16; b_sign3 = 4'd6;
@(posedge clk_i);
a_mant0 = 8'd92; a_mant1 = 8'd11; a_mant2 = 8'd95; a_mant3 = 8'd158;
b_mant0 = 8'd78; b_mant1 = 8'd204; b_mant2 = 8'd221; b_mant3 = 8'd158;
a_exp0 = 10'd831; a_exp1 = 10'd298; a_exp2 = 10'd1015; a_exp3 = 10'd381;
b_exp0 = 10'd170; b_exp1 = 10'd707; b_exp2 = 10'd337; b_exp3 = 10'd633;
a_sign0 = 4'd13; a_sign1 = 4'd10; a_sign2 = 4'd10; a_sign3 = 4'd9;
b_sign0 = 4'd10; b_sign1 = 4'd15; b_sign2 = 4'd11; b_sign3 = 4'd7;
@(posedge clk_i);
a_mant0 = 8'd19; a_mant1 = 8'd132; a_mant2 = 8'd55; a_mant3 = 8'd26;
b_mant0 = 8'd164; b_mant1 = 8'd206; b_mant2 = 8'd177; b_mant3 = 8'd210;
a_exp0 = 10'd783; a_exp1 = 10'd44; a_exp2 = 10'd795; a_exp3 = 10'd334;
b_exp0 = 10'd185; b_exp1 = 10'd56; b_exp2 = 10'd76; b_exp3 = 10'd112;
a_sign0 = 4'd6; a_sign1 = 4'd10; a_sign2 = 4'd1; a_sign3 = 4'd6;
b_sign0 = 4'd14; b_sign1 = 4'd1; b_sign2 = 4'd6; b_sign3 = 4'd8;
@(posedge clk_i);
a_mant0 = 8'd182; a_mant1 = 8'd36; a_mant2 = 8'd14; a_mant3 = 8'd23;
b_mant0 = 8'd170; b_mant1 = 8'd74; b_mant2 = 8'd28; b_mant3 = 8'd143;
a_exp0 = 10'd914; a_exp1 = 10'd22; a_exp2 = 10'd657; a_exp3 = 10'd178;
b_exp0 = 10'd277; b_exp1 = 10'd445; b_exp2 = 10'd1017; b_exp3 = 10'd642;
a_sign0 = 4'd1; a_sign1 = 4'd15; a_sign2 = 4'd4; a_sign3 = 4'd8;
b_sign0 = 4'd3; b_sign1 = 4'd15; b_sign2 = 4'd2; b_sign3 = 4'd14;
@(posedge clk_i);
a_mant0 = 8'd138; a_mant1 = 8'd15; a_mant2 = 8'd255; a_mant3 = 8'd121;
b_mant0 = 8'd102; b_mant1 = 8'd230; b_mant2 = 8'd206; b_mant3 = 8'd75;
a_exp0 = 10'd520; a_exp1 = 10'd461; a_exp2 = 10'd151; a_exp3 = 10'd676;
b_exp0 = 10'd185; b_exp1 = 10'd288; b_exp2 = 10'd471; b_exp3 = 10'd627;
a_sign0 = 4'd1; a_sign1 = 4'd8; a_sign2 = 4'd1; a_sign3 = 4'd7;
b_sign0 = 4'd13; b_sign1 = 4'd0; b_sign2 = 4'd1; b_sign3 = 4'd4;
@(posedge clk_i);
shared_exps0 = 8'd136;
shared_exps1 = 8'd111;
a_mant0 = 8'd188; a_mant1 = 8'd61; a_mant2 = 8'd193; a_mant3 = 8'd207;
b_mant0 = 8'd227; b_mant1 = 8'd21; b_mant2 = 8'd43; b_mant3 = 8'd55;
a_exp0 = 10'd896; a_exp1 = 10'd199; a_exp2 = 10'd549; a_exp3 = 10'd251;
b_exp0 = 10'd735; b_exp1 = 10'd709; b_exp2 = 10'd343; b_exp3 = 10'd146;
a_sign0 = 4'd11; a_sign1 = 4'd2; a_sign2 = 4'd10; a_sign3 = 4'd8;
b_sign0 = 4'd4; b_sign1 = 4'd8; b_sign2 = 4'd12; b_sign3 = 4'd8;
@(posedge clk_i);
a_mant0 = 8'd81; a_mant1 = 8'd70; a_mant2 = 8'd118; a_mant3 = 8'd56;
b_mant0 = 8'd203; b_mant1 = 8'd63; b_mant2 = 8'd152; b_mant3 = 8'd10;
a_exp0 = 10'd462; a_exp1 = 10'd470; a_exp2 = 10'd531; a_exp3 = 10'd277;
b_exp0 = 10'd921; b_exp1 = 10'd111; b_exp2 = 10'd370; b_exp3 = 10'd558;
a_sign0 = 4'd10; a_sign1 = 4'd1; a_sign2 = 4'd1; a_sign3 = 4'd12;
b_sign0 = 4'd9; b_sign1 = 4'd14; b_sign2 = 4'd9; b_sign3 = 4'd4;
@(posedge clk_i);
a_mant0 = 8'd97; a_mant1 = 8'd156; a_mant2 = 8'd27; a_mant3 = 8'd254;
b_mant0 = 8'd199; b_mant1 = 8'd151; b_mant2 = 8'd252; b_mant3 = 8'd153;
a_exp0 = 10'd168; a_exp1 = 10'd214; a_exp2 = 10'd528; a_exp3 = 10'd1015;
b_exp0 = 10'd936; b_exp1 = 10'd214; b_exp2 = 10'd935; b_exp3 = 10'd520;
a_sign0 = 4'd5; a_sign1 = 4'd6; a_sign2 = 4'd15; a_sign3 = 4'd15;
b_sign0 = 4'd14; b_sign1 = 4'd8; b_sign2 = 4'd11; b_sign3 = 4'd16;
@(posedge clk_i);
a_mant0 = 8'd79; a_mant1 = 8'd139; a_mant2 = 8'd30; a_mant3 = 8'd153;
b_mant0 = 8'd78; b_mant1 = 8'd222; b_mant2 = 8'd65; b_mant3 = 8'd170;
a_exp0 = 10'd940; a_exp1 = 10'd225; a_exp2 = 10'd650; a_exp3 = 10'd612;
b_exp0 = 10'd913; b_exp1 = 10'd592; b_exp2 = 10'd571; b_exp3 = 10'd518;
a_sign0 = 4'd16; a_sign1 = 4'd6; a_sign2 = 4'd14; a_sign3 = 4'd15;
b_sign0 = 4'd0; b_sign1 = 4'd16; b_sign2 = 4'd14; b_sign3 = 4'd16;
@(posedge clk_i);
a_mant0 = 8'd100; a_mant1 = 8'd98; a_mant2 = 8'd94; a_mant3 = 8'd36;
b_mant0 = 8'd144; b_mant1 = 8'd41; b_mant2 = 8'd161; b_mant3 = 8'd82;
a_exp0 = 10'd746; a_exp1 = 10'd801; a_exp2 = 10'd357; a_exp3 = 10'd263;
b_exp0 = 10'd661; b_exp1 = 10'd220; b_exp2 = 10'd788; b_exp3 = 10'd295;
a_sign0 = 4'd1; a_sign1 = 4'd16; a_sign2 = 4'd8; a_sign3 = 4'd12;
b_sign0 = 4'd9; b_sign1 = 4'd16; b_sign2 = 4'd12; b_sign3 = 4'd14;
@(posedge clk_i);
a_mant0 = 8'd85; a_mant1 = 8'd29; a_mant2 = 8'd138; a_mant3 = 8'd25;
b_mant0 = 8'd169; b_mant1 = 8'd66; b_mant2 = 8'd221; b_mant3 = 8'd239;
a_exp0 = 10'd462; a_exp1 = 10'd859; a_exp2 = 10'd775; a_exp3 = 10'd235;
b_exp0 = 10'd881; b_exp1 = 10'd611; b_exp2 = 10'd103; b_exp3 = 10'd554;
a_sign0 = 4'd4; a_sign1 = 4'd10; a_sign2 = 4'd12; a_sign3 = 4'd10;
b_sign0 = 4'd0; b_sign1 = 4'd5; b_sign2 = 4'd16; b_sign3 = 4'd7;
@(posedge clk_i);
a_mant0 = 8'd150; a_mant1 = 8'd227; a_mant2 = 8'd205; a_mant3 = 8'd246;
b_mant0 = 8'd10; b_mant1 = 8'd3; b_mant2 = 8'd221; b_mant3 = 8'd51;
a_exp0 = 10'd478; a_exp1 = 10'd858; a_exp2 = 10'd949; a_exp3 = 10'd33;
b_exp0 = 10'd859; b_exp1 = 10'd251; b_exp2 = 10'd993; b_exp3 = 10'd440;
a_sign0 = 4'd6; a_sign1 = 4'd1; a_sign2 = 4'd13; a_sign3 = 4'd2;
b_sign0 = 4'd7; b_sign1 = 4'd13; b_sign2 = 4'd6; b_sign3 = 4'd3;
@(posedge clk_i);
a_mant0 = 8'd203; a_mant1 = 8'd65; a_mant2 = 8'd140; a_mant3 = 8'd239;
b_mant0 = 8'd15; b_mant1 = 8'd245; b_mant2 = 8'd23; b_mant3 = 8'd2;
a_exp0 = 10'd90; a_exp1 = 10'd3; a_exp2 = 10'd514; a_exp3 = 10'd822;
b_exp0 = 10'd795; b_exp1 = 10'd914; b_exp2 = 10'd802; b_exp3 = 10'd931;
a_sign0 = 4'd10; a_sign1 = 4'd16; a_sign2 = 4'd8; a_sign3 = 4'd0;
b_sign0 = 4'd10; b_sign1 = 4'd0; b_sign2 = 4'd1; b_sign3 = 4'd15;
@(posedge clk_i);
shared_exps0 = 8'd123;
shared_exps1 = 8'd98;
a_mant0 = 8'd95; a_mant1 = 8'd159; a_mant2 = 8'd148; a_mant3 = 8'd31;
b_mant0 = 8'd120; b_mant1 = 8'd168; b_mant2 = 8'd194; b_mant3 = 8'd25;
a_exp0 = 10'd298; a_exp1 = 10'd14; a_exp2 = 10'd6; a_exp3 = 10'd906;
b_exp0 = 10'd258; b_exp1 = 10'd348; b_exp2 = 10'd997; b_exp3 = 10'd818;
a_sign0 = 4'd10; a_sign1 = 4'd12; a_sign2 = 4'd5; a_sign3 = 4'd1;
b_sign0 = 4'd6; b_sign1 = 4'd8; b_sign2 = 4'd8; b_sign3 = 4'd15;
@(posedge clk_i);
a_mant0 = 8'd222; a_mant1 = 8'd121; a_mant2 = 8'd85; a_mant3 = 8'd167;
b_mant0 = 8'd146; b_mant1 = 8'd116; b_mant2 = 8'd238; b_mant3 = 8'd162;
a_exp0 = 10'd949; a_exp1 = 10'd963; a_exp2 = 10'd145; a_exp3 = 10'd467;
b_exp0 = 10'd547; b_exp1 = 10'd335; b_exp2 = 10'd200; b_exp3 = 10'd962;
a_sign0 = 4'd11; a_sign1 = 4'd4; a_sign2 = 4'd8; a_sign3 = 4'd10;
b_sign0 = 4'd12; b_sign1 = 4'd11; b_sign2 = 4'd15; b_sign3 = 4'd7;
@(posedge clk_i);
a_mant0 = 8'd147; a_mant1 = 8'd60; a_mant2 = 8'd77; a_mant3 = 8'd89;
b_mant0 = 8'd85; b_mant1 = 8'd50; b_mant2 = 8'd51; b_mant3 = 8'd57;
a_exp0 = 10'd24; a_exp1 = 10'd199; a_exp2 = 10'd352; a_exp3 = 10'd49;
b_exp0 = 10'd932; b_exp1 = 10'd143; b_exp2 = 10'd882; b_exp3 = 10'd226;
a_sign0 = 4'd11; a_sign1 = 4'd10; a_sign2 = 4'd6; a_sign3 = 4'd15;
b_sign0 = 4'd10; b_sign1 = 4'd8; b_sign2 = 4'd9; b_sign3 = 4'd11;
@(posedge clk_i);
a_mant0 = 8'd135; a_mant1 = 8'd230; a_mant2 = 8'd148; a_mant3 = 8'd194;
b_mant0 = 8'd213; b_mant1 = 8'd30; b_mant2 = 8'd136; b_mant3 = 8'd195;
a_exp0 = 10'd316; a_exp1 = 10'd195; a_exp2 = 10'd308; a_exp3 = 10'd271;
b_exp0 = 10'd233; b_exp1 = 10'd898; b_exp2 = 10'd933; b_exp3 = 10'd362;
a_sign0 = 4'd1; a_sign1 = 4'd16; a_sign2 = 4'd6; a_sign3 = 4'd4;
b_sign0 = 4'd14; b_sign1 = 4'd9; b_sign2 = 4'd5; b_sign3 = 4'd12;
@(posedge clk_i);
a_mant0 = 8'd67; a_mant1 = 8'd89; a_mant2 = 8'd49; a_mant3 = 8'd186;
b_mant0 = 8'd77; b_mant1 = 8'd70; b_mant2 = 8'd65; b_mant3 = 8'd188;
a_exp0 = 10'd925; a_exp1 = 10'd750; a_exp2 = 10'd103; a_exp3 = 10'd902;
b_exp0 = 10'd158; b_exp1 = 10'd686; b_exp2 = 10'd858; b_exp3 = 10'd695;
a_sign0 = 4'd6; a_sign1 = 4'd11; a_sign2 = 4'd2; a_sign3 = 4'd12;
b_sign0 = 4'd1; b_sign1 = 4'd16; b_sign2 = 4'd14; b_sign3 = 4'd12;
@(posedge clk_i);
a_mant0 = 8'd161; a_mant1 = 8'd41; a_mant2 = 8'd134; a_mant3 = 8'd200;
b_mant0 = 8'd122; b_mant1 = 8'd127; b_mant2 = 8'd69; b_mant3 = 8'd140;
a_exp0 = 10'd764; a_exp1 = 10'd1020; a_exp2 = 10'd11; a_exp3 = 10'd73;
b_exp0 = 10'd652; b_exp1 = 10'd893; b_exp2 = 10'd248; b_exp3 = 10'd579;
a_sign0 = 4'd0; a_sign1 = 4'd3; a_sign2 = 4'd16; a_sign3 = 4'd16;
b_sign0 = 4'd12; b_sign1 = 4'd2; b_sign2 = 4'd8; b_sign3 = 4'd9;
@(posedge clk_i);
a_mant0 = 8'd218; a_mant1 = 8'd65; a_mant2 = 8'd185; a_mant3 = 8'd20;
b_mant0 = 8'd54; b_mant1 = 8'd223; b_mant2 = 8'd107; b_mant3 = 8'd38;
a_exp0 = 10'd694; a_exp1 = 10'd716; a_exp2 = 10'd601; a_exp3 = 10'd413;
b_exp0 = 10'd923; b_exp1 = 10'd85; b_exp2 = 10'd329; b_exp3 = 10'd280;
a_sign0 = 4'd4; a_sign1 = 4'd11; a_sign2 = 4'd12; a_sign3 = 4'd13;
b_sign0 = 4'd3; b_sign1 = 4'd15; b_sign2 = 4'd3; b_sign3 = 4'd7;
@(posedge clk_i);
a_mant0 = 8'd171; a_mant1 = 8'd0; a_mant2 = 8'd182; a_mant3 = 8'd105;
b_mant0 = 8'd215; b_mant1 = 8'd94; b_mant2 = 8'd69; b_mant3 = 8'd63;
a_exp0 = 10'd1016; a_exp1 = 10'd625; a_exp2 = 10'd151; a_exp3 = 10'd795;
b_exp0 = 10'd605; b_exp1 = 10'd144; b_exp2 = 10'd626; b_exp3 = 10'd809;
a_sign0 = 4'd5; a_sign1 = 4'd4; a_sign2 = 4'd1; a_sign3 = 4'd11;
b_sign0 = 4'd2; b_sign1 = 4'd8; b_sign2 = 4'd10; b_sign3 = 4'd8;
@(posedge clk_i);
shared_exps0 = 8'd128;
shared_exps1 = 8'd120;
rstn = 0;
@(posedge clk_i);
rstn = 1;
a_mant0 = 8'd9; a_mant1 = 8'd254; a_mant2 = 8'd102; a_mant3 = 8'd114;
b_mant0 = 8'd196; b_mant1 = 8'd172; b_mant2 = 8'd142; b_mant3 = 8'd57;
a_exp0 = 10'd985; a_exp1 = 10'd575; a_exp2 = 10'd236; a_exp3 = 10'd407;
b_exp0 = 10'd847; b_exp1 = 10'd895; b_exp2 = 10'd918; b_exp3 = 10'd579;
a_sign0 = 4'd11; a_sign1 = 4'd7; a_sign2 = 4'd10; a_sign3 = 4'd12;
b_sign0 = 4'd14; b_sign1 = 4'd7; b_sign2 = 4'd8; b_sign3 = 4'd7;
@(posedge clk_i);
a_mant0 = 8'd247; a_mant1 = 8'd80; a_mant2 = 8'd26; a_mant3 = 8'd113;
b_mant0 = 8'd203; b_mant1 = 8'd13; b_mant2 = 8'd215; b_mant3 = 8'd65;
a_exp0 = 10'd151; a_exp1 = 10'd118; a_exp2 = 10'd26; a_exp3 = 10'd235;
b_exp0 = 10'd932; b_exp1 = 10'd412; b_exp2 = 10'd52; b_exp3 = 10'd701;
a_sign0 = 4'd7; a_sign1 = 4'd13; a_sign2 = 4'd3; a_sign3 = 4'd10;
b_sign0 = 4'd12; b_sign1 = 4'd3; b_sign2 = 4'd10; b_sign3 = 4'd10;
@(posedge clk_i);
a_mant0 = 8'd9; a_mant1 = 8'd106; a_mant2 = 8'd11; a_mant3 = 8'd37;
b_mant0 = 8'd226; b_mant1 = 8'd97; b_mant2 = 8'd24; b_mant3 = 8'd193;
a_exp0 = 10'd94; a_exp1 = 10'd104; a_exp2 = 10'd276; a_exp3 = 10'd658;
b_exp0 = 10'd244; b_exp1 = 10'd919; b_exp2 = 10'd61; b_exp3 = 10'd313;
a_sign0 = 4'd15; a_sign1 = 4'd16; a_sign2 = 4'd7; a_sign3 = 4'd4;
b_sign0 = 4'd10; b_sign1 = 4'd10; b_sign2 = 4'd1; b_sign3 = 4'd1;
@(posedge clk_i);
a_mant0 = 8'd125; a_mant1 = 8'd44; a_mant2 = 8'd214; a_mant3 = 8'd124;
b_mant0 = 8'd236; b_mant1 = 8'd88; b_mant2 = 8'd250; b_mant3 = 8'd151;
a_exp0 = 10'd169; a_exp1 = 10'd990; a_exp2 = 10'd852; a_exp3 = 10'd327;
b_exp0 = 10'd821; b_exp1 = 10'd307; b_exp2 = 10'd385; b_exp3 = 10'd1008;
a_sign0 = 4'd9; a_sign1 = 4'd12; a_sign2 = 4'd0; a_sign3 = 4'd12;
b_sign0 = 4'd9; b_sign1 = 4'd12; b_sign2 = 4'd8; b_sign3 = 4'd12;
@(posedge clk_i);
a_mant0 = 8'd157; a_mant1 = 8'd36; a_mant2 = 8'd102; a_mant3 = 8'd234;
b_mant0 = 8'd155; b_mant1 = 8'd75; b_mant2 = 8'd30; b_mant3 = 8'd156;
a_exp0 = 10'd487; a_exp1 = 10'd466; a_exp2 = 10'd646; a_exp3 = 10'd400;
b_exp0 = 10'd678; b_exp1 = 10'd481; b_exp2 = 10'd240; b_exp3 = 10'd636;
a_sign0 = 4'd14; a_sign1 = 4'd12; a_sign2 = 4'd2; a_sign3 = 4'd2;
b_sign0 = 4'd14; b_sign1 = 4'd5; b_sign2 = 4'd16; b_sign3 = 4'd0;
@(posedge clk_i);
a_mant0 = 8'd82; a_mant1 = 8'd212; a_mant2 = 8'd189; a_mant3 = 8'd28;
b_mant0 = 8'd111; b_mant1 = 8'd244; b_mant2 = 8'd29; b_mant3 = 8'd40;
a_exp0 = 10'd950; a_exp1 = 10'd457; a_exp2 = 10'd723; a_exp3 = 10'd692;
b_exp0 = 10'd582; b_exp1 = 10'd671; b_exp2 = 10'd400; b_exp3 = 10'd1010;
a_sign0 = 4'd15; a_sign1 = 4'd5; a_sign2 = 4'd9; a_sign3 = 4'd3;
b_sign0 = 4'd14; b_sign1 = 4'd5; b_sign2 = 4'd0; b_sign3 = 4'd13;
@(posedge clk_i);
a_mant0 = 8'd12; a_mant1 = 8'd189; a_mant2 = 8'd3; a_mant3 = 8'd241;
b_mant0 = 8'd70; b_mant1 = 8'd40; b_mant2 = 8'd239; b_mant3 = 8'd228;
a_exp0 = 10'd257; a_exp1 = 10'd512; a_exp2 = 10'd195; a_exp3 = 10'd249;
b_exp0 = 10'd909; b_exp1 = 10'd434; b_exp2 = 10'd372; b_exp3 = 10'd887;
a_sign0 = 4'd15; a_sign1 = 4'd0; a_sign2 = 4'd14; a_sign3 = 4'd15;
b_sign0 = 4'd8; b_sign1 = 4'd11; b_sign2 = 4'd13; b_sign3 = 4'd15;
@(posedge clk_i);
shared_exps0 = 8'd132;
shared_exps1 = 8'd137;
a_mant0 = 8'd63; a_mant1 = 8'd131; a_mant2 = 8'd44; a_mant3 = 8'd178;
b_mant0 = 8'd175; b_mant1 = 8'd94; b_mant2 = 8'd169; b_mant3 = 8'd219;
a_exp0 = 10'd429; a_exp1 = 10'd932; a_exp2 = 10'd536; a_exp3 = 10'd257;
b_exp0 = 10'd616; b_exp1 = 10'd425; b_exp2 = 10'd33; b_exp3 = 10'd532;
a_sign0 = 4'd7; a_sign1 = 4'd8; a_sign2 = 4'd11; a_sign3 = 4'd10;
b_sign0 = 4'd9; b_sign1 = 4'd13; b_sign2 = 4'd6; b_sign3 = 4'd13;
@(posedge clk_i);
a_mant0 = 8'd77; a_mant1 = 8'd166; a_mant2 = 8'd158; a_mant3 = 8'd244;
b_mant0 = 8'd209; b_mant1 = 8'd148; b_mant2 = 8'd221; b_mant3 = 8'd173;
a_exp0 = 10'd431; a_exp1 = 10'd317; a_exp2 = 10'd62; a_exp3 = 10'd17;
b_exp0 = 10'd509; b_exp1 = 10'd425; b_exp2 = 10'd184; b_exp3 = 10'd482;
a_sign0 = 4'd5; a_sign1 = 4'd16; a_sign2 = 4'd7; a_sign3 = 4'd14;
b_sign0 = 4'd1; b_sign1 = 4'd2; b_sign2 = 4'd9; b_sign3 = 4'd8;
@(posedge clk_i);
a_mant0 = 8'd83; a_mant1 = 8'd77; a_mant2 = 8'd145; a_mant3 = 8'd45;
b_mant0 = 8'd185; b_mant1 = 8'd179; b_mant2 = 8'd14; b_mant3 = 8'd168;
a_exp0 = 10'd575; a_exp1 = 10'd817; a_exp2 = 10'd548; a_exp3 = 10'd429;
b_exp0 = 10'd246; b_exp1 = 10'd1008; b_exp2 = 10'd447; b_exp3 = 10'd252;
a_sign0 = 4'd6; a_sign1 = 4'd6; a_sign2 = 4'd1; a_sign3 = 4'd3;
b_sign0 = 4'd5; b_sign1 = 4'd10; b_sign2 = 4'd10; b_sign3 = 4'd13;
@(posedge clk_i);
a_mant0 = 8'd86; a_mant1 = 8'd245; a_mant2 = 8'd243; a_mant3 = 8'd61;
b_mant0 = 8'd29; b_mant1 = 8'd31; b_mant2 = 8'd45; b_mant3 = 8'd28;
a_exp0 = 10'd580; a_exp1 = 10'd286; a_exp2 = 10'd781; a_exp3 = 10'd565;
b_exp0 = 10'd817; b_exp1 = 10'd993; b_exp2 = 10'd582; b_exp3 = 10'd886;
a_sign0 = 4'd8; a_sign1 = 4'd9; a_sign2 = 4'd16; a_sign3 = 4'd2;
b_sign0 = 4'd5; b_sign1 = 4'd11; b_sign2 = 4'd12; b_sign3 = 4'd10;
@(posedge clk_i);
a_mant0 = 8'd201; a_mant1 = 8'd166; a_mant2 = 8'd98; a_mant3 = 8'd226;
b_mant0 = 8'd221; b_mant1 = 8'd184; b_mant2 = 8'd140; b_mant3 = 8'd151;
a_exp0 = 10'd547; a_exp1 = 10'd688; a_exp2 = 10'd703; a_exp3 = 10'd78;
b_exp0 = 10'd293; b_exp1 = 10'd347; b_exp2 = 10'd30; b_exp3 = 10'd106;
a_sign0 = 4'd7; a_sign1 = 4'd8; a_sign2 = 4'd9; a_sign3 = 4'd9;
b_sign0 = 4'd1; b_sign1 = 4'd0; b_sign2 = 4'd9; b_sign3 = 4'd6;
@(posedge clk_i);
a_mant0 = 8'd65; a_mant1 = 8'd148; a_mant2 = 8'd77; a_mant3 = 8'd109;
b_mant0 = 8'd179; b_mant1 = 8'd186; b_mant2 = 8'd187; b_mant3 = 8'd240;
a_exp0 = 10'd357; a_exp1 = 10'd841; a_exp2 = 10'd832; a_exp3 = 10'd705;
b_exp0 = 10'd699; b_exp1 = 10'd734; b_exp2 = 10'd13; b_exp3 = 10'd445;
a_sign0 = 4'd11; a_sign1 = 4'd3; a_sign2 = 4'd12; a_sign3 = 4'd7;
b_sign0 = 4'd7; b_sign1 = 4'd3; b_sign2 = 4'd8; b_sign3 = 4'd8;
@(posedge clk_i);
a_mant0 = 8'd71; a_mant1 = 8'd125; a_mant2 = 8'd61; a_mant3 = 8'd33;
b_mant0 = 8'd194; b_mant1 = 8'd100; b_mant2 = 8'd98; b_mant3 = 8'd170;
a_exp0 = 10'd442; a_exp1 = 10'd687; a_exp2 = 10'd632; a_exp3 = 10'd732;
b_exp0 = 10'd1000; b_exp1 = 10'd281; b_exp2 = 10'd999; b_exp3 = 10'd606;
a_sign0 = 4'd7; a_sign1 = 4'd13; a_sign2 = 4'd3; a_sign3 = 4'd0;
b_sign0 = 4'd11; b_sign1 = 4'd3; b_sign2 = 4'd12; b_sign3 = 4'd6;
@(posedge clk_i);
a_mant0 = 8'd225; a_mant1 = 8'd29; a_mant2 = 8'd193; a_mant3 = 8'd192;
b_mant0 = 8'd136; b_mant1 = 8'd234; b_mant2 = 8'd153; b_mant3 = 8'd23;
a_exp0 = 10'd649; a_exp1 = 10'd556; a_exp2 = 10'd279; a_exp3 = 10'd601;
b_exp0 = 10'd601; b_exp1 = 10'd398; b_exp2 = 10'd576; b_exp3 = 10'd235;
a_sign0 = 4'd5; a_sign1 = 4'd9; a_sign2 = 4'd0; a_sign3 = 4'd5;
b_sign0 = 4'd7; b_sign1 = 4'd15; b_sign2 = 4'd6; b_sign3 = 4'd1;
@(posedge clk_i);
shared_exps0 = 8'd129;
shared_exps1 = 8'd132;
a_mant0 = 8'd189; a_mant1 = 8'd69; a_mant2 = 8'd25; a_mant3 = 8'd62;
b_mant0 = 8'd42; b_mant1 = 8'd1; b_mant2 = 8'd183; b_mant3 = 8'd161;
a_exp0 = 10'd948; a_exp1 = 10'd388; a_exp2 = 10'd1015; a_exp3 = 10'd993;
b_exp0 = 10'd343; b_exp1 = 10'd699; b_exp2 = 10'd258; b_exp3 = 10'd372;
a_sign0 = 4'd3; a_sign1 = 4'd2; a_sign2 = 4'd15; a_sign3 = 4'd3;
b_sign0 = 4'd7; b_sign1 = 4'd14; b_sign2 = 4'd5; b_sign3 = 4'd15;
@(posedge clk_i);
a_mant0 = 8'd3; a_mant1 = 8'd115; a_mant2 = 8'd185; a_mant3 = 8'd170;
b_mant0 = 8'd29; b_mant1 = 8'd198; b_mant2 = 8'd152; b_mant3 = 8'd67;
a_exp0 = 10'd789; a_exp1 = 10'd318; a_exp2 = 10'd668; a_exp3 = 10'd506;
b_exp0 = 10'd807; b_exp1 = 10'd590; b_exp2 = 10'd595; b_exp3 = 10'd452;
a_sign0 = 4'd15; a_sign1 = 4'd5; a_sign2 = 4'd15; a_sign3 = 4'd6;
b_sign0 = 4'd8; b_sign1 = 4'd7; b_sign2 = 4'd9; b_sign3 = 4'd4;
@(posedge clk_i);
a_mant0 = 8'd168; a_mant1 = 8'd198; a_mant2 = 8'd33; a_mant3 = 8'd246;
b_mant0 = 8'd1; b_mant1 = 8'd101; b_mant2 = 8'd59; b_mant3 = 8'd250;
a_exp0 = 10'd754; a_exp1 = 10'd923; a_exp2 = 10'd228; a_exp3 = 10'd485;
b_exp0 = 10'd453; b_exp1 = 10'd593; b_exp2 = 10'd560; b_exp3 = 10'd327;
a_sign0 = 4'd7; a_sign1 = 4'd2; a_sign2 = 4'd14; a_sign3 = 4'd7;
b_sign0 = 4'd4; b_sign1 = 4'd1; b_sign2 = 4'd10; b_sign3 = 4'd14;
@(posedge clk_i);
a_mant0 = 8'd162; a_mant1 = 8'd145; a_mant2 = 8'd242; a_mant3 = 8'd212;
b_mant0 = 8'd228; b_mant1 = 8'd130; b_mant2 = 8'd43; b_mant3 = 8'd202;
a_exp0 = 10'd844; a_exp1 = 10'd475; a_exp2 = 10'd386; a_exp3 = 10'd441;
b_exp0 = 10'd990; b_exp1 = 10'd574; b_exp2 = 10'd243; b_exp3 = 10'd408;
a_sign0 = 4'd2; a_sign1 = 4'd4; a_sign2 = 4'd6; a_sign3 = 4'd4;
b_sign0 = 4'd6; b_sign1 = 4'd8; b_sign2 = 4'd7; b_sign3 = 4'd9;
@(posedge clk_i);
a_mant0 = 8'd37; a_mant1 = 8'd21; a_mant2 = 8'd45; a_mant3 = 8'd55;
b_mant0 = 8'd41; b_mant1 = 8'd232; b_mant2 = 8'd150; b_mant3 = 8'd241;
a_exp0 = 10'd83; a_exp1 = 10'd90; a_exp2 = 10'd633; a_exp3 = 10'd178;
b_exp0 = 10'd590; b_exp1 = 10'd657; b_exp2 = 10'd161; b_exp3 = 10'd80;
a_sign0 = 4'd15; a_sign1 = 4'd7; a_sign2 = 4'd11; a_sign3 = 4'd13;
b_sign0 = 4'd3; b_sign1 = 4'd8; b_sign2 = 4'd4; b_sign3 = 4'd6;
@(posedge clk_i);
a_mant0 = 8'd14; a_mant1 = 8'd184; a_mant2 = 8'd149; a_mant3 = 8'd175;
b_mant0 = 8'd41; b_mant1 = 8'd98; b_mant2 = 8'd25; b_mant3 = 8'd101;
a_exp0 = 10'd1002; a_exp1 = 10'd879; a_exp2 = 10'd1000; a_exp3 = 10'd1006;
b_exp0 = 10'd340; b_exp1 = 10'd521; b_exp2 = 10'd879; b_exp3 = 10'd362;
a_sign0 = 4'd9; a_sign1 = 4'd11; a_sign2 = 4'd16; a_sign3 = 4'd4;
b_sign0 = 4'd2; b_sign1 = 4'd14; b_sign2 = 4'd11; b_sign3 = 4'd10;
@(posedge clk_i);
a_mant0 = 8'd96; a_mant1 = 8'd60; a_mant2 = 8'd126; a_mant3 = 8'd208;
b_mant0 = 8'd63; b_mant1 = 8'd185; b_mant2 = 8'd115; b_mant3 = 8'd229;
a_exp0 = 10'd226; a_exp1 = 10'd576; a_exp2 = 10'd287; a_exp3 = 10'd913;
b_exp0 = 10'd419; b_exp1 = 10'd269; b_exp2 = 10'd832; b_exp3 = 10'd91;
a_sign0 = 4'd7; a_sign1 = 4'd11; a_sign2 = 4'd6; a_sign3 = 4'd1;
b_sign0 = 4'd12; b_sign1 = 4'd5; b_sign2 = 4'd12; b_sign3 = 4'd15;
@(posedge clk_i);
a_mant0 = 8'd153; a_mant1 = 8'd225; a_mant2 = 8'd233; a_mant3 = 8'd245;
b_mant0 = 8'd138; b_mant1 = 8'd155; b_mant2 = 8'd239; b_mant3 = 8'd4;
a_exp0 = 10'd341; a_exp1 = 10'd178; a_exp2 = 10'd992; a_exp3 = 10'd751;
b_exp0 = 10'd315; b_exp1 = 10'd80; b_exp2 = 10'd716; b_exp3 = 10'd847;
a_sign0 = 4'd10; a_sign1 = 4'd12; a_sign2 = 4'd5; a_sign3 = 4'd3;
b_sign0 = 4'd7; b_sign1 = 4'd11; b_sign2 = 4'd6; b_sign3 = 4'd5;
@(posedge clk_i);
shared_exps0 = 8'd155;
shared_exps1 = 8'd134;
a_mant0 = 8'd139; a_mant1 = 8'd113; a_mant2 = 8'd152; a_mant3 = 8'd54;
b_mant0 = 8'd105; b_mant1 = 8'd145; b_mant2 = 8'd249; b_mant3 = 8'd12;
a_exp0 = 10'd260; a_exp1 = 10'd564; a_exp2 = 10'd986; a_exp3 = 10'd69;
b_exp0 = 10'd290; b_exp1 = 10'd241; b_exp2 = 10'd991; b_exp3 = 10'd999;
a_sign0 = 4'd11; a_sign1 = 4'd10; a_sign2 = 4'd1; a_sign3 = 4'd6;
b_sign0 = 4'd3; b_sign1 = 4'd13; b_sign2 = 4'd7; b_sign3 = 4'd5;
@(posedge clk_i);
a_mant0 = 8'd86; a_mant1 = 8'd181; a_mant2 = 8'd106; a_mant3 = 8'd169;
b_mant0 = 8'd48; b_mant1 = 8'd248; b_mant2 = 8'd86; b_mant3 = 8'd123;
a_exp0 = 10'd405; a_exp1 = 10'd79; a_exp2 = 10'd563; a_exp3 = 10'd385;
b_exp0 = 10'd817; b_exp1 = 10'd749; b_exp2 = 10'd361; b_exp3 = 10'd932;
a_sign0 = 4'd1; a_sign1 = 4'd16; a_sign2 = 4'd1; a_sign3 = 4'd5;
b_sign0 = 4'd8; b_sign1 = 4'd9; b_sign2 = 4'd4; b_sign3 = 4'd0;
@(posedge clk_i);
a_mant0 = 8'd190; a_mant1 = 8'd0; a_mant2 = 8'd51; a_mant3 = 8'd14;
b_mant0 = 8'd181; b_mant1 = 8'd112; b_mant2 = 8'd212; b_mant3 = 8'd132;
a_exp0 = 10'd921; a_exp1 = 10'd857; a_exp2 = 10'd439; a_exp3 = 10'd297;
b_exp0 = 10'd841; b_exp1 = 10'd1011; b_exp2 = 10'd379; b_exp3 = 10'd762;
a_sign0 = 4'd3; a_sign1 = 4'd8; a_sign2 = 4'd10; a_sign3 = 4'd3;
b_sign0 = 4'd10; b_sign1 = 4'd1; b_sign2 = 4'd16; b_sign3 = 4'd12;
@(posedge clk_i);
a_mant0 = 8'd116; a_mant1 = 8'd118; a_mant2 = 8'd237; a_mant3 = 8'd56;
b_mant0 = 8'd27; b_mant1 = 8'd129; b_mant2 = 8'd228; b_mant3 = 8'd162;
a_exp0 = 10'd142; a_exp1 = 10'd630; a_exp2 = 10'd995; a_exp3 = 10'd487;
b_exp0 = 10'd579; b_exp1 = 10'd1015; b_exp2 = 10'd507; b_exp3 = 10'd293;
a_sign0 = 4'd13; a_sign1 = 4'd14; a_sign2 = 4'd14; a_sign3 = 4'd6;
b_sign0 = 4'd15; b_sign1 = 4'd1; b_sign2 = 4'd5; b_sign3 = 4'd14;
@(posedge clk_i);
a_mant0 = 8'd10; a_mant1 = 8'd162; a_mant2 = 8'd208; a_mant3 = 8'd71;
b_mant0 = 8'd65; b_mant1 = 8'd211; b_mant2 = 8'd128; b_mant3 = 8'd159;
a_exp0 = 10'd802; a_exp1 = 10'd143; a_exp2 = 10'd243; a_exp3 = 10'd731;
b_exp0 = 10'd355; b_exp1 = 10'd973; b_exp2 = 10'd603; b_exp3 = 10'd848;
a_sign0 = 4'd16; a_sign1 = 4'd0; a_sign2 = 4'd1; a_sign3 = 4'd11;
b_sign0 = 4'd10; b_sign1 = 4'd7; b_sign2 = 4'd2; b_sign3 = 4'd10;
@(posedge clk_i);
a_mant0 = 8'd28; a_mant1 = 8'd77; a_mant2 = 8'd83; a_mant3 = 8'd98;
b_mant0 = 8'd65; b_mant1 = 8'd48; b_mant2 = 8'd152; b_mant3 = 8'd75;
a_exp0 = 10'd372; a_exp1 = 10'd389; a_exp2 = 10'd405; a_exp3 = 10'd538;
b_exp0 = 10'd663; b_exp1 = 10'd510; b_exp2 = 10'd844; b_exp3 = 10'd387;
a_sign0 = 4'd0; a_sign1 = 4'd10; a_sign2 = 4'd4; a_sign3 = 4'd5;
b_sign0 = 4'd1; b_sign1 = 4'd7; b_sign2 = 4'd0; b_sign3 = 4'd0;
@(posedge clk_i);
a_mant0 = 8'd122; a_mant1 = 8'd150; a_mant2 = 8'd33; a_mant3 = 8'd42;
b_mant0 = 8'd156; b_mant1 = 8'd212; b_mant2 = 8'd222; b_mant3 = 8'd59;
a_exp0 = 10'd1018; a_exp1 = 10'd995; a_exp2 = 10'd467; a_exp3 = 10'd711;
b_exp0 = 10'd143; b_exp1 = 10'd852; b_exp2 = 10'd45; b_exp3 = 10'd115;
a_sign0 = 4'd2; a_sign1 = 4'd12; a_sign2 = 4'd0; a_sign3 = 4'd1;
b_sign0 = 4'd12; b_sign1 = 4'd5; b_sign2 = 4'd3; b_sign3 = 4'd7;
@(posedge clk_i);
a_mant0 = 8'd155; a_mant1 = 8'd128; a_mant2 = 8'd240; a_mant3 = 8'd34;
b_mant0 = 8'd137; b_mant1 = 8'd232; b_mant2 = 8'd238; b_mant3 = 8'd50;
a_exp0 = 10'd268; a_exp1 = 10'd741; a_exp2 = 10'd734; a_exp3 = 10'd297;
b_exp0 = 10'd814; b_exp1 = 10'd729; b_exp2 = 10'd998; b_exp3 = 10'd535;
a_sign0 = 4'd11; a_sign1 = 4'd4; a_sign2 = 4'd13; a_sign3 = 4'd6;
b_sign0 = 4'd14; b_sign1 = 4'd14; b_sign2 = 4'd1; b_sign3 = 4'd16;
@(posedge clk_i);
shared_exps0 = 8'd153;
shared_exps1 = 8'd122;
rstn = 0;
@(posedge clk_i);
rstn = 1;
a_mant0 = 8'd7; a_mant1 = 8'd213; a_mant2 = 8'd17; a_mant3 = 8'd140;
b_mant0 = 8'd223; b_mant1 = 8'd106; b_mant2 = 8'd91; b_mant3 = 8'd238;
a_exp0 = 10'd476; a_exp1 = 10'd596; a_exp2 = 10'd587; a_exp3 = 10'd164;
b_exp0 = 10'd473; b_exp1 = 10'd116; b_exp2 = 10'd861; b_exp3 = 10'd309;
a_sign0 = 4'd8; a_sign1 = 4'd5; a_sign2 = 4'd6; a_sign3 = 4'd10;
b_sign0 = 4'd12; b_sign1 = 4'd0; b_sign2 = 4'd2; b_sign3 = 4'd15;
@(posedge clk_i);
a_mant0 = 8'd29; a_mant1 = 8'd237; a_mant2 = 8'd149; a_mant3 = 8'd136;
b_mant0 = 8'd38; b_mant1 = 8'd209; b_mant2 = 8'd66; b_mant3 = 8'd153;
a_exp0 = 10'd740; a_exp1 = 10'd109; a_exp2 = 10'd766; a_exp3 = 10'd998;
b_exp0 = 10'd750; b_exp1 = 10'd616; b_exp2 = 10'd182; b_exp3 = 10'd568;
a_sign0 = 4'd11; a_sign1 = 4'd0; a_sign2 = 4'd10; a_sign3 = 4'd13;
b_sign0 = 4'd16; b_sign1 = 4'd13; b_sign2 = 4'd8; b_sign3 = 4'd13;
@(posedge clk_i);
a_mant0 = 8'd8; a_mant1 = 8'd13; a_mant2 = 8'd198; a_mant3 = 8'd230;
b_mant0 = 8'd149; b_mant1 = 8'd83; b_mant2 = 8'd48; b_mant3 = 8'd10;
a_exp0 = 10'd601; a_exp1 = 10'd798; a_exp2 = 10'd855; a_exp3 = 10'd817;
b_exp0 = 10'd560; b_exp1 = 10'd847; b_exp2 = 10'd898; b_exp3 = 10'd346;
a_sign0 = 4'd2; a_sign1 = 4'd16; a_sign2 = 4'd3; a_sign3 = 4'd12;
b_sign0 = 4'd16; b_sign1 = 4'd4; b_sign2 = 4'd14; b_sign3 = 4'd16;
@(posedge clk_i);
a_mant0 = 8'd246; a_mant1 = 8'd65; a_mant2 = 8'd49; a_mant3 = 8'd201;
b_mant0 = 8'd207; b_mant1 = 8'd79; b_mant2 = 8'd8; b_mant3 = 8'd232;
a_exp0 = 10'd841; a_exp1 = 10'd270; a_exp2 = 10'd783; a_exp3 = 10'd478;
b_exp0 = 10'd503; b_exp1 = 10'd30; b_exp2 = 10'd143; b_exp3 = 10'd878;
a_sign0 = 4'd9; a_sign1 = 4'd14; a_sign2 = 4'd7; a_sign3 = 4'd5;
b_sign0 = 4'd14; b_sign1 = 4'd10; b_sign2 = 4'd9; b_sign3 = 4'd7;
@(posedge clk_i);
a_mant0 = 8'd54; a_mant1 = 8'd171; a_mant2 = 8'd247; a_mant3 = 8'd217;
b_mant0 = 8'd205; b_mant1 = 8'd208; b_mant2 = 8'd236; b_mant3 = 8'd35;
a_exp0 = 10'd236; a_exp1 = 10'd935; a_exp2 = 10'd702; a_exp3 = 10'd46;
b_exp0 = 10'd527; b_exp1 = 10'd863; b_exp2 = 10'd951; b_exp3 = 10'd336;
a_sign0 = 4'd16; a_sign1 = 4'd8; a_sign2 = 4'd16; a_sign3 = 4'd8;
b_sign0 = 4'd8; b_sign1 = 4'd15; b_sign2 = 4'd13; b_sign3 = 4'd15;
@(posedge clk_i);
a_mant0 = 8'd173; a_mant1 = 8'd135; a_mant2 = 8'd210; a_mant3 = 8'd197;
b_mant0 = 8'd204; b_mant1 = 8'd199; b_mant2 = 8'd219; b_mant3 = 8'd168;
a_exp0 = 10'd274; a_exp1 = 10'd185; a_exp2 = 10'd599; a_exp3 = 10'd424;
b_exp0 = 10'd370; b_exp1 = 10'd373; b_exp2 = 10'd38; b_exp3 = 10'd983;
a_sign0 = 4'd12; a_sign1 = 4'd11; a_sign2 = 4'd12; a_sign3 = 4'd2;
b_sign0 = 4'd12; b_sign1 = 4'd13; b_sign2 = 4'd15; b_sign3 = 4'd1;
@(posedge clk_i);
a_mant0 = 8'd127; a_mant1 = 8'd88; a_mant2 = 8'd216; a_mant3 = 8'd79;
b_mant0 = 8'd172; b_mant1 = 8'd189; b_mant2 = 8'd246; b_mant3 = 8'd145;
a_exp0 = 10'd652; a_exp1 = 10'd442; a_exp2 = 10'd998; a_exp3 = 10'd73;
b_exp0 = 10'd759; b_exp1 = 10'd399; b_exp2 = 10'd777; b_exp3 = 10'd649;
a_sign0 = 4'd8; a_sign1 = 4'd3; a_sign2 = 4'd8; a_sign3 = 4'd16;
b_sign0 = 4'd2; b_sign1 = 4'd1; b_sign2 = 4'd6; b_sign3 = 4'd13;
@(posedge clk_i);
shared_exps0 = 8'd93;
shared_exps1 = 8'd142;
a_mant0 = 8'd126; a_mant1 = 8'd167; a_mant2 = 8'd104; a_mant3 = 8'd228;
b_mant0 = 8'd114; b_mant1 = 8'd76; b_mant2 = 8'd157; b_mant3 = 8'd245;
a_exp0 = 10'd418; a_exp1 = 10'd167; a_exp2 = 10'd1000; a_exp3 = 10'd390;
b_exp0 = 10'd1023; b_exp1 = 10'd81; b_exp2 = 10'd9; b_exp3 = 10'd533;
a_sign0 = 4'd12; a_sign1 = 4'd1; a_sign2 = 4'd6; a_sign3 = 4'd2;
b_sign0 = 4'd15; b_sign1 = 4'd6; b_sign2 = 4'd0; b_sign3 = 4'd14;
@(posedge clk_i);
a_mant0 = 8'd50; a_mant1 = 8'd25; a_mant2 = 8'd113; a_mant3 = 8'd240;
b_mant0 = 8'd64; b_mant1 = 8'd143; b_mant2 = 8'd197; b_mant3 = 8'd78;
a_exp0 = 10'd699; a_exp1 = 10'd475; a_exp2 = 10'd17; a_exp3 = 10'd200;
b_exp0 = 10'd261; b_exp1 = 10'd939; b_exp2 = 10'd307; b_exp3 = 10'd885;
a_sign0 = 4'd8; a_sign1 = 4'd13; a_sign2 = 4'd10; a_sign3 = 4'd12;
b_sign0 = 4'd1; b_sign1 = 4'd5; b_sign2 = 4'd3; b_sign3 = 4'd1;
@(posedge clk_i);
a_mant0 = 8'd203; a_mant1 = 8'd83; a_mant2 = 8'd11; a_mant3 = 8'd28;
b_mant0 = 8'd85; b_mant1 = 8'd248; b_mant2 = 8'd238; b_mant3 = 8'd152;
a_exp0 = 10'd119; a_exp1 = 10'd617; a_exp2 = 10'd637; a_exp3 = 10'd202;
b_exp0 = 10'd251; b_exp1 = 10'd683; b_exp2 = 10'd441; b_exp3 = 10'd989;
a_sign0 = 4'd16; a_sign1 = 4'd2; a_sign2 = 4'd8; a_sign3 = 4'd2;
b_sign0 = 4'd6; b_sign1 = 4'd3; b_sign2 = 4'd15; b_sign3 = 4'd8;
@(posedge clk_i);
a_mant0 = 8'd139; a_mant1 = 8'd118; a_mant2 = 8'd125; a_mant3 = 8'd142;
b_mant0 = 8'd168; b_mant1 = 8'd214; b_mant2 = 8'd18; b_mant3 = 8'd217;
a_exp0 = 10'd19; a_exp1 = 10'd839; a_exp2 = 10'd1021; a_exp3 = 10'd499;
b_exp0 = 10'd564; b_exp1 = 10'd857; b_exp2 = 10'd168; b_exp3 = 10'd901;
a_sign0 = 4'd5; a_sign1 = 4'd5; a_sign2 = 4'd7; a_sign3 = 4'd16;
b_sign0 = 4'd8; b_sign1 = 4'd6; b_sign2 = 4'd5; b_sign3 = 4'd14;
@(posedge clk_i);
a_mant0 = 8'd152; a_mant1 = 8'd134; a_mant2 = 8'd16; a_mant3 = 8'd23;
b_mant0 = 8'd102; b_mant1 = 8'd112; b_mant2 = 8'd17; b_mant3 = 8'd23;
a_exp0 = 10'd860; a_exp1 = 10'd713; a_exp2 = 10'd640; a_exp3 = 10'd521;
b_exp0 = 10'd871; b_exp1 = 10'd502; b_exp2 = 10'd547; b_exp3 = 10'd233;
a_sign0 = 4'd8; a_sign1 = 4'd4; a_sign2 = 4'd2; a_sign3 = 4'd1;
b_sign0 = 4'd6; b_sign1 = 4'd6; b_sign2 = 4'd16; b_sign3 = 4'd8;
@(posedge clk_i);
a_mant0 = 8'd218; a_mant1 = 8'd54; a_mant2 = 8'd177; a_mant3 = 8'd219;
b_mant0 = 8'd25; b_mant1 = 8'd250; b_mant2 = 8'd227; b_mant3 = 8'd144;
a_exp0 = 10'd324; a_exp1 = 10'd677; a_exp2 = 10'd70; a_exp3 = 10'd609;
b_exp0 = 10'd164; b_exp1 = 10'd70; b_exp2 = 10'd82; b_exp3 = 10'd146;
a_sign0 = 4'd13; a_sign1 = 4'd13; a_sign2 = 4'd6; a_sign3 = 4'd0;
b_sign0 = 4'd11; b_sign1 = 4'd7; b_sign2 = 4'd11; b_sign3 = 4'd3;
@(posedge clk_i);
a_mant0 = 8'd108; a_mant1 = 8'd86; a_mant2 = 8'd143; a_mant3 = 8'd189;
b_mant0 = 8'd94; b_mant1 = 8'd253; b_mant2 = 8'd180; b_mant3 = 8'd97;
a_exp0 = 10'd660; a_exp1 = 10'd413; a_exp2 = 10'd902; a_exp3 = 10'd734;
b_exp0 = 10'd707; b_exp1 = 10'd373; b_exp2 = 10'd131; b_exp3 = 10'd107;
a_sign0 = 4'd15; a_sign1 = 4'd12; a_sign2 = 4'd10; a_sign3 = 4'd8;
b_sign0 = 4'd8; b_sign1 = 4'd9; b_sign2 = 4'd12; b_sign3 = 4'd15;
@(posedge clk_i);
a_mant0 = 8'd5; a_mant1 = 8'd23; a_mant2 = 8'd187; a_mant3 = 8'd189;
b_mant0 = 8'd197; b_mant1 = 8'd41; b_mant2 = 8'd207; b_mant3 = 8'd35;
a_exp0 = 10'd347; a_exp1 = 10'd732; a_exp2 = 10'd96; a_exp3 = 10'd318;
b_exp0 = 10'd630; b_exp1 = 10'd801; b_exp2 = 10'd516; b_exp3 = 10'd780;
a_sign0 = 4'd8; a_sign1 = 4'd8; a_sign2 = 4'd1; a_sign3 = 4'd13;
b_sign0 = 4'd12; b_sign1 = 4'd11; b_sign2 = 4'd16; b_sign3 = 4'd14;
@(posedge clk_i);
shared_exps0 = 8'd108;
shared_exps1 = 8'd122;
a_mant0 = 8'd228; a_mant1 = 8'd223; a_mant2 = 8'd215; a_mant3 = 8'd61;
b_mant0 = 8'd131; b_mant1 = 8'd151; b_mant2 = 8'd19; b_mant3 = 8'd107;
a_exp0 = 10'd758; a_exp1 = 10'd709; a_exp2 = 10'd770; a_exp3 = 10'd1007;
b_exp0 = 10'd128; b_exp1 = 10'd393; b_exp2 = 10'd157; b_exp3 = 10'd756;
a_sign0 = 4'd11; a_sign1 = 4'd11; a_sign2 = 4'd8; a_sign3 = 4'd15;
b_sign0 = 4'd14; b_sign1 = 4'd4; b_sign2 = 4'd10; b_sign3 = 4'd13;
@(posedge clk_i);
a_mant0 = 8'd140; a_mant1 = 8'd33; a_mant2 = 8'd236; a_mant3 = 8'd152;
b_mant0 = 8'd232; b_mant1 = 8'd230; b_mant2 = 8'd123; b_mant3 = 8'd223;
a_exp0 = 10'd71; a_exp1 = 10'd656; a_exp2 = 10'd68; a_exp3 = 10'd909;
b_exp0 = 10'd656; b_exp1 = 10'd543; b_exp2 = 10'd1015; b_exp3 = 10'd500;
a_sign0 = 4'd0; a_sign1 = 4'd13; a_sign2 = 4'd2; a_sign3 = 4'd12;
b_sign0 = 4'd7; b_sign1 = 4'd13; b_sign2 = 4'd13; b_sign3 = 4'd3;
@(posedge clk_i);
a_mant0 = 8'd90; a_mant1 = 8'd195; a_mant2 = 8'd189; a_mant3 = 8'd139;
b_mant0 = 8'd34; b_mant1 = 8'd79; b_mant2 = 8'd244; b_mant3 = 8'd4;
a_exp0 = 10'd722; a_exp1 = 10'd373; a_exp2 = 10'd250; a_exp3 = 10'd305;
b_exp0 = 10'd887; b_exp1 = 10'd516; b_exp2 = 10'd838; b_exp3 = 10'd346;
a_sign0 = 4'd7; a_sign1 = 4'd13; a_sign2 = 4'd8; a_sign3 = 4'd0;
b_sign0 = 4'd2; b_sign1 = 4'd3; b_sign2 = 4'd7; b_sign3 = 4'd10;
@(posedge clk_i);
a_mant0 = 8'd110; a_mant1 = 8'd225; a_mant2 = 8'd54; a_mant3 = 8'd140;
b_mant0 = 8'd147; b_mant1 = 8'd49; b_mant2 = 8'd218; b_mant3 = 8'd131;
a_exp0 = 10'd912; a_exp1 = 10'd991; a_exp2 = 10'd642; a_exp3 = 10'd409;
b_exp0 = 10'd257; b_exp1 = 10'd859; b_exp2 = 10'd163; b_exp3 = 10'd707;
a_sign0 = 4'd3; a_sign1 = 4'd5; a_sign2 = 4'd9; a_sign3 = 4'd6;
b_sign0 = 4'd5; b_sign1 = 4'd12; b_sign2 = 4'd13; b_sign3 = 4'd5;
@(posedge clk_i);
a_mant0 = 8'd104; a_mant1 = 8'd150; a_mant2 = 8'd0; a_mant3 = 8'd201;
b_mant0 = 8'd48; b_mant1 = 8'd184; b_mant2 = 8'd250; b_mant3 = 8'd203;
a_exp0 = 10'd284; a_exp1 = 10'd296; a_exp2 = 10'd563; a_exp3 = 10'd422;
b_exp0 = 10'd84; b_exp1 = 10'd450; b_exp2 = 10'd694; b_exp3 = 10'd828;
a_sign0 = 4'd16; a_sign1 = 4'd5; a_sign2 = 4'd4; a_sign3 = 4'd4;
b_sign0 = 4'd8; b_sign1 = 4'd0; b_sign2 = 4'd10; b_sign3 = 4'd0;
@(posedge clk_i);
a_mant0 = 8'd234; a_mant1 = 8'd57; a_mant2 = 8'd147; a_mant3 = 8'd17;
b_mant0 = 8'd205; b_mant1 = 8'd175; b_mant2 = 8'd13; b_mant3 = 8'd207;
a_exp0 = 10'd699; a_exp1 = 10'd939; a_exp2 = 10'd315; a_exp3 = 10'd716;
b_exp0 = 10'd1015; b_exp1 = 10'd623; b_exp2 = 10'd124; b_exp3 = 10'd524;
a_sign0 = 4'd15; a_sign1 = 4'd4; a_sign2 = 4'd4; a_sign3 = 4'd8;
b_sign0 = 4'd5; b_sign1 = 4'd12; b_sign2 = 4'd10; b_sign3 = 4'd5;
@(posedge clk_i);
a_mant0 = 8'd43; a_mant1 = 8'd108; a_mant2 = 8'd163; a_mant3 = 8'd153;
b_mant0 = 8'd126; b_mant1 = 8'd73; b_mant2 = 8'd174; b_mant3 = 8'd74;
a_exp0 = 10'd653; a_exp1 = 10'd69; a_exp2 = 10'd167; a_exp3 = 10'd978;
b_exp0 = 10'd713; b_exp1 = 10'd819; b_exp2 = 10'd293; b_exp3 = 10'd703;
a_sign0 = 4'd0; a_sign1 = 4'd0; a_sign2 = 4'd12; a_sign3 = 4'd5;
b_sign0 = 4'd10; b_sign1 = 4'd6; b_sign2 = 4'd1; b_sign3 = 4'd0;
@(posedge clk_i);
a_mant0 = 8'd34; a_mant1 = 8'd198; a_mant2 = 8'd237; a_mant3 = 8'd49;
b_mant0 = 8'd43; b_mant1 = 8'd248; b_mant2 = 8'd43; b_mant3 = 8'd10;
a_exp0 = 10'd786; a_exp1 = 10'd726; a_exp2 = 10'd3; a_exp3 = 10'd638;
b_exp0 = 10'd70; b_exp1 = 10'd966; b_exp2 = 10'd110; b_exp3 = 10'd479;
a_sign0 = 4'd14; a_sign1 = 4'd13; a_sign2 = 4'd5; a_sign3 = 4'd11;
b_sign0 = 4'd3; b_sign1 = 4'd10; b_sign2 = 4'd1; b_sign3 = 4'd11;
@(posedge clk_i);
shared_exps0 = 8'd127;
shared_exps1 = 8'd129;
a_mant0 = 8'd84; a_mant1 = 8'd232; a_mant2 = 8'd213; a_mant3 = 8'd170;
b_mant0 = 8'd16; b_mant1 = 8'd232; b_mant2 = 8'd248; b_mant3 = 8'd241;
a_exp0 = 10'd173; a_exp1 = 10'd913; a_exp2 = 10'd65; a_exp3 = 10'd250;
b_exp0 = 10'd87; b_exp1 = 10'd81; b_exp2 = 10'd671; b_exp3 = 10'd34;
a_sign0 = 4'd13; a_sign1 = 4'd2; a_sign2 = 4'd7; a_sign3 = 4'd11;
b_sign0 = 4'd11; b_sign1 = 4'd6; b_sign2 = 4'd9; b_sign3 = 4'd16;
@(posedge clk_i);
a_mant0 = 8'd8; a_mant1 = 8'd76; a_mant2 = 8'd175; a_mant3 = 8'd43;
b_mant0 = 8'd42; b_mant1 = 8'd30; b_mant2 = 8'd143; b_mant3 = 8'd37;
a_exp0 = 10'd235; a_exp1 = 10'd544; a_exp2 = 10'd554; a_exp3 = 10'd814;
b_exp0 = 10'd104; b_exp1 = 10'd338; b_exp2 = 10'd323; b_exp3 = 10'd765;
a_sign0 = 4'd13; a_sign1 = 4'd12; a_sign2 = 4'd6; a_sign3 = 4'd8;
b_sign0 = 4'd4; b_sign1 = 4'd5; b_sign2 = 4'd5; b_sign3 = 4'd6;
@(posedge clk_i);
a_mant0 = 8'd133; a_mant1 = 8'd251; a_mant2 = 8'd139; a_mant3 = 8'd28;
b_mant0 = 8'd85; b_mant1 = 8'd103; b_mant2 = 8'd244; b_mant3 = 8'd225;
a_exp0 = 10'd940; a_exp1 = 10'd1; a_exp2 = 10'd545; a_exp3 = 10'd568;
b_exp0 = 10'd311; b_exp1 = 10'd938; b_exp2 = 10'd677; b_exp3 = 10'd42;
a_sign0 = 4'd8; a_sign1 = 4'd2; a_sign2 = 4'd10; a_sign3 = 4'd1;
b_sign0 = 4'd9; b_sign1 = 4'd1; b_sign2 = 4'd15; b_sign3 = 4'd13;
@(posedge clk_i);
a_mant0 = 8'd147; a_mant1 = 8'd216; a_mant2 = 8'd15; a_mant3 = 8'd196;
b_mant0 = 8'd122; b_mant1 = 8'd88; b_mant2 = 8'd170; b_mant3 = 8'd80;
a_exp0 = 10'd47; a_exp1 = 10'd261; a_exp2 = 10'd963; a_exp3 = 10'd553;
b_exp0 = 10'd437; b_exp1 = 10'd781; b_exp2 = 10'd517; b_exp3 = 10'd673;
a_sign0 = 4'd9; a_sign1 = 4'd12; a_sign2 = 4'd0; a_sign3 = 4'd0;
b_sign0 = 4'd8; b_sign1 = 4'd15; b_sign2 = 4'd2; b_sign3 = 4'd8;
@(posedge clk_i);
a_mant0 = 8'd152; a_mant1 = 8'd108; a_mant2 = 8'd202; a_mant3 = 8'd187;
b_mant0 = 8'd3; b_mant1 = 8'd190; b_mant2 = 8'd65; b_mant3 = 8'd99;
a_exp0 = 10'd690; a_exp1 = 10'd945; a_exp2 = 10'd529; a_exp3 = 10'd82;
b_exp0 = 10'd479; b_exp1 = 10'd182; b_exp2 = 10'd749; b_exp3 = 10'd129;
a_sign0 = 4'd8; a_sign1 = 4'd14; a_sign2 = 4'd7; a_sign3 = 4'd6;
b_sign0 = 4'd6; b_sign1 = 4'd3; b_sign2 = 4'd9; b_sign3 = 4'd10;
@(posedge clk_i);
a_mant0 = 8'd175; a_mant1 = 8'd69; a_mant2 = 8'd224; a_mant3 = 8'd153;
b_mant0 = 8'd80; b_mant1 = 8'd43; b_mant2 = 8'd20; b_mant3 = 8'd159;
a_exp0 = 10'd93; a_exp1 = 10'd706; a_exp2 = 10'd218; a_exp3 = 10'd1016;
b_exp0 = 10'd981; b_exp1 = 10'd641; b_exp2 = 10'd735; b_exp3 = 10'd927;
a_sign0 = 4'd13; a_sign1 = 4'd12; a_sign2 = 4'd11; a_sign3 = 4'd3;
b_sign0 = 4'd11; b_sign1 = 4'd5; b_sign2 = 4'd12; b_sign3 = 4'd2;
@(posedge clk_i);
a_mant0 = 8'd157; a_mant1 = 8'd147; a_mant2 = 8'd145; a_mant3 = 8'd57;
b_mant0 = 8'd245; b_mant1 = 8'd81; b_mant2 = 8'd58; b_mant3 = 8'd219;
a_exp0 = 10'd598; a_exp1 = 10'd179; a_exp2 = 10'd775; a_exp3 = 10'd423;
b_exp0 = 10'd933; b_exp1 = 10'd812; b_exp2 = 10'd979; b_exp3 = 10'd711;
a_sign0 = 4'd5; a_sign1 = 4'd4; a_sign2 = 4'd10; a_sign3 = 4'd15;
b_sign0 = 4'd2; b_sign1 = 4'd10; b_sign2 = 4'd11; b_sign3 = 4'd16;
@(posedge clk_i);
a_mant0 = 8'd87; a_mant1 = 8'd145; a_mant2 = 8'd149; a_mant3 = 8'd133;
b_mant0 = 8'd146; b_mant1 = 8'd8; b_mant2 = 8'd188; b_mant3 = 8'd0;
a_exp0 = 10'd520; a_exp1 = 10'd723; a_exp2 = 10'd667; a_exp3 = 10'd252;
b_exp0 = 10'd729; b_exp1 = 10'd16; b_exp2 = 10'd39; b_exp3 = 10'd296;
a_sign0 = 4'd3; a_sign1 = 4'd5; a_sign2 = 4'd12; a_sign3 = 4'd10;
b_sign0 = 4'd11; b_sign1 = 4'd4; b_sign2 = 4'd11; b_sign3 = 4'd6;
@(posedge clk_i);
shared_exps0 = 8'd153;
shared_exps1 = 8'd114;
rstn = 0;
@(posedge clk_i);
rstn = 1;
a_mant0 = 8'd254; a_mant1 = 8'd157; a_mant2 = 8'd220; a_mant3 = 8'd17;
b_mant0 = 8'd153; b_mant1 = 8'd52; b_mant2 = 8'd81; b_mant3 = 8'd200;
a_exp0 = 10'd887; a_exp1 = 10'd675; a_exp2 = 10'd249; a_exp3 = 10'd130;
b_exp0 = 10'd566; b_exp1 = 10'd378; b_exp2 = 10'd987; b_exp3 = 10'd785;
a_sign0 = 4'd9; a_sign1 = 4'd16; a_sign2 = 4'd16; a_sign3 = 4'd12;
b_sign0 = 4'd4; b_sign1 = 4'd2; b_sign2 = 4'd10; b_sign3 = 4'd13;
@(posedge clk_i);
a_mant0 = 8'd32; a_mant1 = 8'd26; a_mant2 = 8'd19; a_mant3 = 8'd50;
b_mant0 = 8'd61; b_mant1 = 8'd13; b_mant2 = 8'd143; b_mant3 = 8'd91;
a_exp0 = 10'd317; a_exp1 = 10'd964; a_exp2 = 10'd26; a_exp3 = 10'd445;
b_exp0 = 10'd499; b_exp1 = 10'd720; b_exp2 = 10'd916; b_exp3 = 10'd26;
a_sign0 = 4'd6; a_sign1 = 4'd0; a_sign2 = 4'd12; a_sign3 = 4'd4;
b_sign0 = 4'd15; b_sign1 = 4'd16; b_sign2 = 4'd8; b_sign3 = 4'd1;
@(posedge clk_i);
a_mant0 = 8'd174; a_mant1 = 8'd150; a_mant2 = 8'd133; a_mant3 = 8'd160;
b_mant0 = 8'd134; b_mant1 = 8'd12; b_mant2 = 8'd225; b_mant3 = 8'd132;
a_exp0 = 10'd265; a_exp1 = 10'd831; a_exp2 = 10'd280; a_exp3 = 10'd723;
b_exp0 = 10'd525; b_exp1 = 10'd696; b_exp2 = 10'd889; b_exp3 = 10'd825;
a_sign0 = 4'd1; a_sign1 = 4'd5; a_sign2 = 4'd7; a_sign3 = 4'd16;
b_sign0 = 4'd2; b_sign1 = 4'd10; b_sign2 = 4'd3; b_sign3 = 4'd9;
@(posedge clk_i);
a_mant0 = 8'd244; a_mant1 = 8'd254; a_mant2 = 8'd236; a_mant3 = 8'd204;
b_mant0 = 8'd135; b_mant1 = 8'd63; b_mant2 = 8'd238; b_mant3 = 8'd207;
a_exp0 = 10'd314; a_exp1 = 10'd695; a_exp2 = 10'd558; a_exp3 = 10'd382;
b_exp0 = 10'd581; b_exp1 = 10'd970; b_exp2 = 10'd188; b_exp3 = 10'd868;
a_sign0 = 4'd1; a_sign1 = 4'd4; a_sign2 = 4'd14; a_sign3 = 4'd1;
b_sign0 = 4'd5; b_sign1 = 4'd6; b_sign2 = 4'd16; b_sign3 = 4'd14;
@(posedge clk_i);
a_mant0 = 8'd148; a_mant1 = 8'd65; a_mant2 = 8'd97; a_mant3 = 8'd25;
b_mant0 = 8'd157; b_mant1 = 8'd32; b_mant2 = 8'd195; b_mant3 = 8'd147;
a_exp0 = 10'd504; a_exp1 = 10'd714; a_exp2 = 10'd209; a_exp3 = 10'd731;
b_exp0 = 10'd163; b_exp1 = 10'd680; b_exp2 = 10'd301; b_exp3 = 10'd545;
a_sign0 = 4'd8; a_sign1 = 4'd10; a_sign2 = 4'd11; a_sign3 = 4'd11;
b_sign0 = 4'd6; b_sign1 = 4'd5; b_sign2 = 4'd12; b_sign3 = 4'd8;
@(posedge clk_i);
a_mant0 = 8'd240; a_mant1 = 8'd43; a_mant2 = 8'd245; a_mant3 = 8'd186;
b_mant0 = 8'd222; b_mant1 = 8'd240; b_mant2 = 8'd6; b_mant3 = 8'd67;
a_exp0 = 10'd710; a_exp1 = 10'd568; a_exp2 = 10'd951; a_exp3 = 10'd148;
b_exp0 = 10'd140; b_exp1 = 10'd899; b_exp2 = 10'd176; b_exp3 = 10'd317;
a_sign0 = 4'd7; a_sign1 = 4'd5; a_sign2 = 4'd16; a_sign3 = 4'd7;
b_sign0 = 4'd1; b_sign1 = 4'd6; b_sign2 = 4'd1; b_sign3 = 4'd13;
@(posedge clk_i);
a_mant0 = 8'd183; a_mant1 = 8'd183; a_mant2 = 8'd214; a_mant3 = 8'd102;
b_mant0 = 8'd200; b_mant1 = 8'd43; b_mant2 = 8'd145; b_mant3 = 8'd7;
a_exp0 = 10'd775; a_exp1 = 10'd708; a_exp2 = 10'd374; a_exp3 = 10'd439;
b_exp0 = 10'd198; b_exp1 = 10'd896; b_exp2 = 10'd678; b_exp3 = 10'd1022;
a_sign0 = 4'd8; a_sign1 = 4'd10; a_sign2 = 4'd1; a_sign3 = 4'd6;
b_sign0 = 4'd11; b_sign1 = 4'd1; b_sign2 = 4'd0; b_sign3 = 4'd9;
@(posedge clk_i);
shared_exps0 = 8'd146;
shared_exps1 = 8'd144;
a_mant0 = 8'd68; a_mant1 = 8'd161; a_mant2 = 8'd125; a_mant3 = 8'd246;
b_mant0 = 8'd220; b_mant1 = 8'd251; b_mant2 = 8'd4; b_mant3 = 8'd148;
a_exp0 = 10'd773; a_exp1 = 10'd425; a_exp2 = 10'd963; a_exp3 = 10'd827;
b_exp0 = 10'd203; b_exp1 = 10'd394; b_exp2 = 10'd282; b_exp3 = 10'd765;
a_sign0 = 4'd3; a_sign1 = 4'd8; a_sign2 = 4'd11; a_sign3 = 4'd12;
b_sign0 = 4'd13; b_sign1 = 4'd8; b_sign2 = 4'd14; b_sign3 = 4'd9;
@(posedge clk_i);
a_mant0 = 8'd70; a_mant1 = 8'd195; a_mant2 = 8'd252; a_mant3 = 8'd3;
b_mant0 = 8'd87; b_mant1 = 8'd139; b_mant2 = 8'd52; b_mant3 = 8'd67;
a_exp0 = 10'd200; a_exp1 = 10'd186; a_exp2 = 10'd665; a_exp3 = 10'd859;
b_exp0 = 10'd386; b_exp1 = 10'd455; b_exp2 = 10'd712; b_exp3 = 10'd38;
a_sign0 = 4'd11; a_sign1 = 4'd7; a_sign2 = 4'd11; a_sign3 = 4'd6;
b_sign0 = 4'd15; b_sign1 = 4'd10; b_sign2 = 4'd3; b_sign3 = 4'd10;
@(posedge clk_i);
a_mant0 = 8'd175; a_mant1 = 8'd180; a_mant2 = 8'd121; a_mant3 = 8'd46;
b_mant0 = 8'd184; b_mant1 = 8'd40; b_mant2 = 8'd153; b_mant3 = 8'd226;
a_exp0 = 10'd686; a_exp1 = 10'd66; a_exp2 = 10'd308; a_exp3 = 10'd117;
b_exp0 = 10'd849; b_exp1 = 10'd977; b_exp2 = 10'd991; b_exp3 = 10'd111;
a_sign0 = 4'd8; a_sign1 = 4'd2; a_sign2 = 4'd9; a_sign3 = 4'd7;
b_sign0 = 4'd8; b_sign1 = 4'd5; b_sign2 = 4'd8; b_sign3 = 4'd4;
@(posedge clk_i);
a_mant0 = 8'd154; a_mant1 = 8'd248; a_mant2 = 8'd104; a_mant3 = 8'd24;
b_mant0 = 8'd210; b_mant1 = 8'd229; b_mant2 = 8'd94; b_mant3 = 8'd186;
a_exp0 = 10'd993; a_exp1 = 10'd848; a_exp2 = 10'd963; a_exp3 = 10'd4;
b_exp0 = 10'd911; b_exp1 = 10'd305; b_exp2 = 10'd488; b_exp3 = 10'd395;
a_sign0 = 4'd5; a_sign1 = 4'd7; a_sign2 = 4'd11; a_sign3 = 4'd14;
b_sign0 = 4'd10; b_sign1 = 4'd0; b_sign2 = 4'd13; b_sign3 = 4'd5;
@(posedge clk_i);
a_mant0 = 8'd167; a_mant1 = 8'd241; a_mant2 = 8'd67; a_mant3 = 8'd35;
b_mant0 = 8'd88; b_mant1 = 8'd52; b_mant2 = 8'd200; b_mant3 = 8'd23;
a_exp0 = 10'd1001; a_exp1 = 10'd108; a_exp2 = 10'd765; a_exp3 = 10'd505;
b_exp0 = 10'd326; b_exp1 = 10'd148; b_exp2 = 10'd855; b_exp3 = 10'd264;
a_sign0 = 4'd5; a_sign1 = 4'd11; a_sign2 = 4'd5; a_sign3 = 4'd8;
b_sign0 = 4'd8; b_sign1 = 4'd0; b_sign2 = 4'd9; b_sign3 = 4'd8;
@(posedge clk_i);
a_mant0 = 8'd110; a_mant1 = 8'd41; a_mant2 = 8'd12; a_mant3 = 8'd161;
b_mant0 = 8'd202; b_mant1 = 8'd84; b_mant2 = 8'd174; b_mant3 = 8'd155;
a_exp0 = 10'd449; a_exp1 = 10'd685; a_exp2 = 10'd594; a_exp3 = 10'd524;
b_exp0 = 10'd939; b_exp1 = 10'd803; b_exp2 = 10'd232; b_exp3 = 10'd487;
a_sign0 = 4'd7; a_sign1 = 4'd1; a_sign2 = 4'd14; a_sign3 = 4'd9;
b_sign0 = 4'd14; b_sign1 = 4'd2; b_sign2 = 4'd15; b_sign3 = 4'd9;
@(posedge clk_i);
a_mant0 = 8'd231; a_mant1 = 8'd43; a_mant2 = 8'd231; a_mant3 = 8'd242;
b_mant0 = 8'd156; b_mant1 = 8'd158; b_mant2 = 8'd150; b_mant3 = 8'd124;
a_exp0 = 10'd38; a_exp1 = 10'd857; a_exp2 = 10'd231; a_exp3 = 10'd110;
b_exp0 = 10'd915; b_exp1 = 10'd367; b_exp2 = 10'd57; b_exp3 = 10'd334;
a_sign0 = 4'd5; a_sign1 = 4'd2; a_sign2 = 4'd1; a_sign3 = 4'd6;
b_sign0 = 4'd1; b_sign1 = 4'd12; b_sign2 = 4'd1; b_sign3 = 4'd4;
@(posedge clk_i);
a_mant0 = 8'd216; a_mant1 = 8'd24; a_mant2 = 8'd245; a_mant3 = 8'd225;
b_mant0 = 8'd215; b_mant1 = 8'd4; b_mant2 = 8'd193; b_mant3 = 8'd205;
a_exp0 = 10'd740; a_exp1 = 10'd817; a_exp2 = 10'd1000; a_exp3 = 10'd446;
b_exp0 = 10'd388; b_exp1 = 10'd374; b_exp2 = 10'd22; b_exp3 = 10'd30;
a_sign0 = 4'd13; a_sign1 = 4'd9; a_sign2 = 4'd2; a_sign3 = 4'd16;
b_sign0 = 4'd2; b_sign1 = 4'd5; b_sign2 = 4'd4; b_sign3 = 4'd6;
@(posedge clk_i);
shared_exps0 = 8'd136;
shared_exps1 = 8'd129;
a_mant0 = 8'd13; a_mant1 = 8'd61; a_mant2 = 8'd254; a_mant3 = 8'd4;
b_mant0 = 8'd98; b_mant1 = 8'd148; b_mant2 = 8'd4; b_mant3 = 8'd15;
a_exp0 = 10'd121; a_exp1 = 10'd686; a_exp2 = 10'd117; a_exp3 = 10'd879;
b_exp0 = 10'd380; b_exp1 = 10'd911; b_exp2 = 10'd415; b_exp3 = 10'd213;
a_sign0 = 4'd12; a_sign1 = 4'd11; a_sign2 = 4'd15; a_sign3 = 4'd6;
b_sign0 = 4'd12; b_sign1 = 4'd1; b_sign2 = 4'd4; b_sign3 = 4'd12;
@(posedge clk_i);
a_mant0 = 8'd169; a_mant1 = 8'd140; a_mant2 = 8'd231; a_mant3 = 8'd112;
b_mant0 = 8'd130; b_mant1 = 8'd179; b_mant2 = 8'd26; b_mant3 = 8'd225;
a_exp0 = 10'd21; a_exp1 = 10'd923; a_exp2 = 10'd379; a_exp3 = 10'd554;
b_exp0 = 10'd554; b_exp1 = 10'd714; b_exp2 = 10'd355; b_exp3 = 10'd846;
a_sign0 = 4'd12; a_sign1 = 4'd10; a_sign2 = 4'd2; a_sign3 = 4'd16;
b_sign0 = 4'd0; b_sign1 = 4'd7; b_sign2 = 4'd6; b_sign3 = 4'd13;
@(posedge clk_i);
a_mant0 = 8'd75; a_mant1 = 8'd240; a_mant2 = 8'd235; a_mant3 = 8'd200;
b_mant0 = 8'd122; b_mant1 = 8'd151; b_mant2 = 8'd59; b_mant3 = 8'd224;
a_exp0 = 10'd457; a_exp1 = 10'd37; a_exp2 = 10'd819; a_exp3 = 10'd352;
b_exp0 = 10'd791; b_exp1 = 10'd861; b_exp2 = 10'd547; b_exp3 = 10'd197;
a_sign0 = 4'd5; a_sign1 = 4'd13; a_sign2 = 4'd9; a_sign3 = 4'd6;
b_sign0 = 4'd3; b_sign1 = 4'd5; b_sign2 = 4'd5; b_sign3 = 4'd10;
@(posedge clk_i);
a_mant0 = 8'd220; a_mant1 = 8'd48; a_mant2 = 8'd173; a_mant3 = 8'd10;
b_mant0 = 8'd52; b_mant1 = 8'd193; b_mant2 = 8'd202; b_mant3 = 8'd244;
a_exp0 = 10'd148; a_exp1 = 10'd699; a_exp2 = 10'd795; a_exp3 = 10'd976;
b_exp0 = 10'd666; b_exp1 = 10'd1017; b_exp2 = 10'd1004; b_exp3 = 10'd984;
a_sign0 = 4'd1; a_sign1 = 4'd13; a_sign2 = 4'd0; a_sign3 = 4'd9;
b_sign0 = 4'd6; b_sign1 = 4'd3; b_sign2 = 4'd11; b_sign3 = 4'd8;
@(posedge clk_i);
a_mant0 = 8'd17; a_mant1 = 8'd84; a_mant2 = 8'd96; a_mant3 = 8'd161;
b_mant0 = 8'd221; b_mant1 = 8'd243; b_mant2 = 8'd49; b_mant3 = 8'd74;
a_exp0 = 10'd68; a_exp1 = 10'd513; a_exp2 = 10'd613; a_exp3 = 10'd679;
b_exp0 = 10'd670; b_exp1 = 10'd349; b_exp2 = 10'd156; b_exp3 = 10'd803;
a_sign0 = 4'd5; a_sign1 = 4'd9; a_sign2 = 4'd13; a_sign3 = 4'd10;
b_sign0 = 4'd12; b_sign1 = 4'd12; b_sign2 = 4'd9; b_sign3 = 4'd8;
@(posedge clk_i);
a_mant0 = 8'd168; a_mant1 = 8'd16; a_mant2 = 8'd232; a_mant3 = 8'd201;
b_mant0 = 8'd6; b_mant1 = 8'd178; b_mant2 = 8'd6; b_mant3 = 8'd210;
a_exp0 = 10'd722; a_exp1 = 10'd967; a_exp2 = 10'd635; a_exp3 = 10'd910;
b_exp0 = 10'd446; b_exp1 = 10'd220; b_exp2 = 10'd593; b_exp3 = 10'd555;
a_sign0 = 4'd16; a_sign1 = 4'd14; a_sign2 = 4'd16; a_sign3 = 4'd5;
b_sign0 = 4'd16; b_sign1 = 4'd5; b_sign2 = 4'd1; b_sign3 = 4'd16;
@(posedge clk_i);
a_mant0 = 8'd198; a_mant1 = 8'd188; a_mant2 = 8'd243; a_mant3 = 8'd240;
b_mant0 = 8'd26; b_mant1 = 8'd36; b_mant2 = 8'd211; b_mant3 = 8'd44;
a_exp0 = 10'd854; a_exp1 = 10'd72; a_exp2 = 10'd758; a_exp3 = 10'd123;
b_exp0 = 10'd140; b_exp1 = 10'd93; b_exp2 = 10'd163; b_exp3 = 10'd713;
a_sign0 = 4'd9; a_sign1 = 4'd16; a_sign2 = 4'd3; a_sign3 = 4'd4;
b_sign0 = 4'd1; b_sign1 = 4'd14; b_sign2 = 4'd13; b_sign3 = 4'd2;
@(posedge clk_i);
a_mant0 = 8'd246; a_mant1 = 8'd223; a_mant2 = 8'd138; a_mant3 = 8'd139;
b_mant0 = 8'd150; b_mant1 = 8'd31; b_mant2 = 8'd76; b_mant3 = 8'd203;
a_exp0 = 10'd279; a_exp1 = 10'd366; a_exp2 = 10'd647; a_exp3 = 10'd850;
b_exp0 = 10'd967; b_exp1 = 10'd298; b_exp2 = 10'd193; b_exp3 = 10'd951;
a_sign0 = 4'd9; a_sign1 = 4'd2; a_sign2 = 4'd2; a_sign3 = 4'd6;
b_sign0 = 4'd13; b_sign1 = 4'd11; b_sign2 = 4'd13; b_sign3 = 4'd3;
@(posedge clk_i);
shared_exps0 = 8'd157;
shared_exps1 = 8'd116;
a_mant0 = 8'd207; a_mant1 = 8'd13; a_mant2 = 8'd196; a_mant3 = 8'd112;
b_mant0 = 8'd142; b_mant1 = 8'd109; b_mant2 = 8'd37; b_mant3 = 8'd83;
a_exp0 = 10'd216; a_exp1 = 10'd92; a_exp2 = 10'd837; a_exp3 = 10'd886;
b_exp0 = 10'd876; b_exp1 = 10'd300; b_exp2 = 10'd830; b_exp3 = 10'd611;
a_sign0 = 4'd10; a_sign1 = 4'd7; a_sign2 = 4'd3; a_sign3 = 4'd0;
b_sign0 = 4'd1; b_sign1 = 4'd2; b_sign2 = 4'd14; b_sign3 = 4'd16;
@(posedge clk_i);
a_mant0 = 8'd203; a_mant1 = 8'd150; a_mant2 = 8'd89; a_mant3 = 8'd2;
b_mant0 = 8'd200; b_mant1 = 8'd38; b_mant2 = 8'd97; b_mant3 = 8'd40;
a_exp0 = 10'd884; a_exp1 = 10'd287; a_exp2 = 10'd1; a_exp3 = 10'd753;
b_exp0 = 10'd686; b_exp1 = 10'd494; b_exp2 = 10'd90; b_exp3 = 10'd791;
a_sign0 = 4'd3; a_sign1 = 4'd11; a_sign2 = 4'd12; a_sign3 = 4'd7;
b_sign0 = 4'd0; b_sign1 = 4'd7; b_sign2 = 4'd9; b_sign3 = 4'd15;
@(posedge clk_i);
a_mant0 = 8'd124; a_mant1 = 8'd105; a_mant2 = 8'd242; a_mant3 = 8'd11;
b_mant0 = 8'd172; b_mant1 = 8'd143; b_mant2 = 8'd17; b_mant3 = 8'd64;
a_exp0 = 10'd586; a_exp1 = 10'd387; a_exp2 = 10'd721; a_exp3 = 10'd477;
b_exp0 = 10'd38; b_exp1 = 10'd10; b_exp2 = 10'd439; b_exp3 = 10'd906;
a_sign0 = 4'd3; a_sign1 = 4'd14; a_sign2 = 4'd3; a_sign3 = 4'd13;
b_sign0 = 4'd7; b_sign1 = 4'd5; b_sign2 = 4'd8; b_sign3 = 4'd12;
@(posedge clk_i);
a_mant0 = 8'd106; a_mant1 = 8'd185; a_mant2 = 8'd51; a_mant3 = 8'd198;
b_mant0 = 8'd116; b_mant1 = 8'd36; b_mant2 = 8'd102; b_mant3 = 8'd15;
a_exp0 = 10'd35; a_exp1 = 10'd472; a_exp2 = 10'd473; a_exp3 = 10'd302;
b_exp0 = 10'd610; b_exp1 = 10'd392; b_exp2 = 10'd496; b_exp3 = 10'd946;
a_sign0 = 4'd14; a_sign1 = 4'd6; a_sign2 = 4'd12; a_sign3 = 4'd4;
b_sign0 = 4'd10; b_sign1 = 4'd6; b_sign2 = 4'd15; b_sign3 = 4'd12;
@(posedge clk_i);
a_mant0 = 8'd244; a_mant1 = 8'd111; a_mant2 = 8'd248; a_mant3 = 8'd175;
b_mant0 = 8'd108; b_mant1 = 8'd73; b_mant2 = 8'd164; b_mant3 = 8'd51;
a_exp0 = 10'd676; a_exp1 = 10'd518; a_exp2 = 10'd802; a_exp3 = 10'd235;
b_exp0 = 10'd1006; b_exp1 = 10'd181; b_exp2 = 10'd740; b_exp3 = 10'd896;
a_sign0 = 4'd8; a_sign1 = 4'd2; a_sign2 = 4'd15; a_sign3 = 4'd10;
b_sign0 = 4'd13; b_sign1 = 4'd8; b_sign2 = 4'd9; b_sign3 = 4'd11;
@(posedge clk_i);
a_mant0 = 8'd102; a_mant1 = 8'd88; a_mant2 = 8'd173; a_mant3 = 8'd250;
b_mant0 = 8'd109; b_mant1 = 8'd213; b_mant2 = 8'd10; b_mant3 = 8'd56;
a_exp0 = 10'd946; a_exp1 = 10'd461; a_exp2 = 10'd113; a_exp3 = 10'd940;
b_exp0 = 10'd736; b_exp1 = 10'd550; b_exp2 = 10'd141; b_exp3 = 10'd602;
a_sign0 = 4'd3; a_sign1 = 4'd10; a_sign2 = 4'd4; a_sign3 = 4'd3;
b_sign0 = 4'd11; b_sign1 = 4'd1; b_sign2 = 4'd8; b_sign3 = 4'd3;
@(posedge clk_i);
a_mant0 = 8'd47; a_mant1 = 8'd28; a_mant2 = 8'd246; a_mant3 = 8'd79;
b_mant0 = 8'd124; b_mant1 = 8'd143; b_mant2 = 8'd155; b_mant3 = 8'd255;
a_exp0 = 10'd76; a_exp1 = 10'd597; a_exp2 = 10'd752; a_exp3 = 10'd491;
b_exp0 = 10'd566; b_exp1 = 10'd913; b_exp2 = 10'd277; b_exp3 = 10'd334;
a_sign0 = 4'd13; a_sign1 = 4'd7; a_sign2 = 4'd2; a_sign3 = 4'd10;
b_sign0 = 4'd6; b_sign1 = 4'd7; b_sign2 = 4'd15; b_sign3 = 4'd6;
@(posedge clk_i);
a_mant0 = 8'd59; a_mant1 = 8'd117; a_mant2 = 8'd246; a_mant3 = 8'd160;
b_mant0 = 8'd111; b_mant1 = 8'd165; b_mant2 = 8'd119; b_mant3 = 8'd160;
a_exp0 = 10'd930; a_exp1 = 10'd795; a_exp2 = 10'd184; a_exp3 = 10'd889;
b_exp0 = 10'd860; b_exp1 = 10'd1007; b_exp2 = 10'd286; b_exp3 = 10'd678;
a_sign0 = 4'd11; a_sign1 = 4'd14; a_sign2 = 4'd10; a_sign3 = 4'd5;
b_sign0 = 4'd9; b_sign1 = 4'd1; b_sign2 = 4'd2; b_sign3 = 4'd2;
@(posedge clk_i);
shared_exps0 = 8'd131;
shared_exps1 = 8'd132;
rstn = 0;
@(posedge clk_i);
rstn = 1;
a_mant0 = 8'd15; a_mant1 = 8'd111; a_mant2 = 8'd243; a_mant3 = 8'd151;
b_mant0 = 8'd0; b_mant1 = 8'd210; b_mant2 = 8'd58; b_mant3 = 8'd55;
a_exp0 = 10'd405; a_exp1 = 10'd751; a_exp2 = 10'd321; a_exp3 = 10'd66;
b_exp0 = 10'd736; b_exp1 = 10'd554; b_exp2 = 10'd414; b_exp3 = 10'd591;
a_sign0 = 4'd13; a_sign1 = 4'd7; a_sign2 = 4'd4; a_sign3 = 4'd12;
b_sign0 = 4'd15; b_sign1 = 4'd10; b_sign2 = 4'd0; b_sign3 = 4'd8;
@(posedge clk_i);
a_mant0 = 8'd29; a_mant1 = 8'd211; a_mant2 = 8'd200; a_mant3 = 8'd206;
b_mant0 = 8'd199; b_mant1 = 8'd180; b_mant2 = 8'd104; b_mant3 = 8'd114;
a_exp0 = 10'd164; a_exp1 = 10'd118; a_exp2 = 10'd932; a_exp3 = 10'd999;
b_exp0 = 10'd739; b_exp1 = 10'd7; b_exp2 = 10'd551; b_exp3 = 10'd498;
a_sign0 = 4'd4; a_sign1 = 4'd6; a_sign2 = 4'd7; a_sign3 = 4'd14;
b_sign0 = 4'd3; b_sign1 = 4'd14; b_sign2 = 4'd1; b_sign3 = 4'd2;
@(posedge clk_i);
a_mant0 = 8'd196; a_mant1 = 8'd134; a_mant2 = 8'd0; a_mant3 = 8'd154;
b_mant0 = 8'd184; b_mant1 = 8'd162; b_mant2 = 8'd203; b_mant3 = 8'd67;
a_exp0 = 10'd295; a_exp1 = 10'd884; a_exp2 = 10'd290; a_exp3 = 10'd945;
b_exp0 = 10'd349; b_exp1 = 10'd158; b_exp2 = 10'd858; b_exp3 = 10'd651;
a_sign0 = 4'd8; a_sign1 = 4'd3; a_sign2 = 4'd6; a_sign3 = 4'd9;
b_sign0 = 4'd16; b_sign1 = 4'd5; b_sign2 = 4'd13; b_sign3 = 4'd13;
@(posedge clk_i);
a_mant0 = 8'd47; a_mant1 = 8'd225; a_mant2 = 8'd219; a_mant3 = 8'd168;
b_mant0 = 8'd194; b_mant1 = 8'd223; b_mant2 = 8'd86; b_mant3 = 8'd237;
a_exp0 = 10'd4; a_exp1 = 10'd394; a_exp2 = 10'd819; a_exp3 = 10'd126;
b_exp0 = 10'd716; b_exp1 = 10'd658; b_exp2 = 10'd1006; b_exp3 = 10'd411;
a_sign0 = 4'd6; a_sign1 = 4'd11; a_sign2 = 4'd4; a_sign3 = 4'd5;
b_sign0 = 4'd10; b_sign1 = 4'd8; b_sign2 = 4'd0; b_sign3 = 4'd13;
@(posedge clk_i);
a_mant0 = 8'd210; a_mant1 = 8'd118; a_mant2 = 8'd131; a_mant3 = 8'd117;
b_mant0 = 8'd5; b_mant1 = 8'd54; b_mant2 = 8'd99; b_mant3 = 8'd246;
a_exp0 = 10'd664; a_exp1 = 10'd120; a_exp2 = 10'd73; a_exp3 = 10'd567;
b_exp0 = 10'd624; b_exp1 = 10'd967; b_exp2 = 10'd53; b_exp3 = 10'd906;
a_sign0 = 4'd10; a_sign1 = 4'd6; a_sign2 = 4'd7; a_sign3 = 4'd11;
b_sign0 = 4'd5; b_sign1 = 4'd10; b_sign2 = 4'd13; b_sign3 = 4'd6;
@(posedge clk_i);
a_mant0 = 8'd201; a_mant1 = 8'd38; a_mant2 = 8'd29; a_mant3 = 8'd23;
b_mant0 = 8'd202; b_mant1 = 8'd181; b_mant2 = 8'd1; b_mant3 = 8'd61;
a_exp0 = 10'd225; a_exp1 = 10'd62; a_exp2 = 10'd51; a_exp3 = 10'd805;
b_exp0 = 10'd774; b_exp1 = 10'd496; b_exp2 = 10'd95; b_exp3 = 10'd665;
a_sign0 = 4'd8; a_sign1 = 4'd3; a_sign2 = 4'd12; a_sign3 = 4'd15;
b_sign0 = 4'd15; b_sign1 = 4'd16; b_sign2 = 4'd11; b_sign3 = 4'd5;
@(posedge clk_i);
a_mant0 = 8'd27; a_mant1 = 8'd183; a_mant2 = 8'd199; a_mant3 = 8'd104;
b_mant0 = 8'd98; b_mant1 = 8'd47; b_mant2 = 8'd192; b_mant3 = 8'd223;
a_exp0 = 10'd472; a_exp1 = 10'd123; a_exp2 = 10'd149; a_exp3 = 10'd932;
b_exp0 = 10'd264; b_exp1 = 10'd405; b_exp2 = 10'd631; b_exp3 = 10'd966;
a_sign0 = 4'd0; a_sign1 = 4'd8; a_sign2 = 4'd9; a_sign3 = 4'd4;
b_sign0 = 4'd7; b_sign1 = 4'd16; b_sign2 = 4'd4; b_sign3 = 4'd12;
@(posedge clk_i);
shared_exps0 = 8'd120;
shared_exps1 = 8'd126;
a_mant0 = 8'd240; a_mant1 = 8'd115; a_mant2 = 8'd42; a_mant3 = 8'd254;
b_mant0 = 8'd113; b_mant1 = 8'd46; b_mant2 = 8'd32; b_mant3 = 8'd128;
a_exp0 = 10'd808; a_exp1 = 10'd958; a_exp2 = 10'd843; a_exp3 = 10'd445;
b_exp0 = 10'd815; b_exp1 = 10'd735; b_exp2 = 10'd625; b_exp3 = 10'd399;
a_sign0 = 4'd5; a_sign1 = 4'd4; a_sign2 = 4'd6; a_sign3 = 4'd0;
b_sign0 = 4'd16; b_sign1 = 4'd15; b_sign2 = 4'd7; b_sign3 = 4'd6;
@(posedge clk_i);
a_mant0 = 8'd166; a_mant1 = 8'd135; a_mant2 = 8'd4; a_mant3 = 8'd205;
b_mant0 = 8'd20; b_mant1 = 8'd42; b_mant2 = 8'd185; b_mant3 = 8'd21;
a_exp0 = 10'd95; a_exp1 = 10'd512; a_exp2 = 10'd271; a_exp3 = 10'd513;
b_exp0 = 10'd667; b_exp1 = 10'd210; b_exp2 = 10'd741; b_exp3 = 10'd416;
a_sign0 = 4'd11; a_sign1 = 4'd5; a_sign2 = 4'd5; a_sign3 = 4'd14;
b_sign0 = 4'd0; b_sign1 = 4'd15; b_sign2 = 4'd6; b_sign3 = 4'd5;
@(posedge clk_i);
a_mant0 = 8'd26; a_mant1 = 8'd20; a_mant2 = 8'd187; a_mant3 = 8'd91;
b_mant0 = 8'd95; b_mant1 = 8'd144; b_mant2 = 8'd212; b_mant3 = 8'd86;
a_exp0 = 10'd923; a_exp1 = 10'd254; a_exp2 = 10'd275; a_exp3 = 10'd616;
b_exp0 = 10'd250; b_exp1 = 10'd867; b_exp2 = 10'd523; b_exp3 = 10'd20;
a_sign0 = 4'd10; a_sign1 = 4'd14; a_sign2 = 4'd1; a_sign3 = 4'd8;
b_sign0 = 4'd11; b_sign1 = 4'd3; b_sign2 = 4'd12; b_sign3 = 4'd6;
@(posedge clk_i);
a_mant0 = 8'd213; a_mant1 = 8'd96; a_mant2 = 8'd141; a_mant3 = 8'd77;
b_mant0 = 8'd38; b_mant1 = 8'd79; b_mant2 = 8'd162; b_mant3 = 8'd132;
a_exp0 = 10'd795; a_exp1 = 10'd190; a_exp2 = 10'd571; a_exp3 = 10'd975;
b_exp0 = 10'd61; b_exp1 = 10'd99; b_exp2 = 10'd344; b_exp3 = 10'd690;
a_sign0 = 4'd2; a_sign1 = 4'd13; a_sign2 = 4'd4; a_sign3 = 4'd6;
b_sign0 = 4'd12; b_sign1 = 4'd14; b_sign2 = 4'd10; b_sign3 = 4'd12;
@(posedge clk_i);
a_mant0 = 8'd138; a_mant1 = 8'd48; a_mant2 = 8'd62; a_mant3 = 8'd49;
b_mant0 = 8'd171; b_mant1 = 8'd102; b_mant2 = 8'd115; b_mant3 = 8'd226;
a_exp0 = 10'd438; a_exp1 = 10'd671; a_exp2 = 10'd503; a_exp3 = 10'd906;
b_exp0 = 10'd435; b_exp1 = 10'd16; b_exp2 = 10'd216; b_exp3 = 10'd318;
a_sign0 = 4'd15; a_sign1 = 4'd9; a_sign2 = 4'd1; a_sign3 = 4'd12;
b_sign0 = 4'd6; b_sign1 = 4'd14; b_sign2 = 4'd3; b_sign3 = 4'd11;
@(posedge clk_i);
a_mant0 = 8'd219; a_mant1 = 8'd182; a_mant2 = 8'd161; a_mant3 = 8'd158;
b_mant0 = 8'd116; b_mant1 = 8'd238; b_mant2 = 8'd196; b_mant3 = 8'd113;
a_exp0 = 10'd434; a_exp1 = 10'd405; a_exp2 = 10'd546; a_exp3 = 10'd69;
b_exp0 = 10'd846; b_exp1 = 10'd944; b_exp2 = 10'd424; b_exp3 = 10'd343;
a_sign0 = 4'd12; a_sign1 = 4'd4; a_sign2 = 4'd15; a_sign3 = 4'd6;
b_sign0 = 4'd16; b_sign1 = 4'd14; b_sign2 = 4'd9; b_sign3 = 4'd13;
@(posedge clk_i);
a_mant0 = 8'd106; a_mant1 = 8'd191; a_mant2 = 8'd250; a_mant3 = 8'd197;
b_mant0 = 8'd13; b_mant1 = 8'd25; b_mant2 = 8'd93; b_mant3 = 8'd45;
a_exp0 = 10'd355; a_exp1 = 10'd996; a_exp2 = 10'd742; a_exp3 = 10'd138;
b_exp0 = 10'd1005; b_exp1 = 10'd39; b_exp2 = 10'd939; b_exp3 = 10'd14;
a_sign0 = 4'd0; a_sign1 = 4'd13; a_sign2 = 4'd15; a_sign3 = 4'd8;
b_sign0 = 4'd3; b_sign1 = 4'd1; b_sign2 = 4'd13; b_sign3 = 4'd8;
@(posedge clk_i);
a_mant0 = 8'd211; a_mant1 = 8'd60; a_mant2 = 8'd11; a_mant3 = 8'd141;
b_mant0 = 8'd209; b_mant1 = 8'd50; b_mant2 = 8'd33; b_mant3 = 8'd43;
a_exp0 = 10'd771; a_exp1 = 10'd314; a_exp2 = 10'd216; a_exp3 = 10'd21;
b_exp0 = 10'd9; b_exp1 = 10'd272; b_exp2 = 10'd681; b_exp3 = 10'd79;
a_sign0 = 4'd6; a_sign1 = 4'd4; a_sign2 = 4'd1; a_sign3 = 4'd0;
b_sign0 = 4'd8; b_sign1 = 4'd7; b_sign2 = 4'd11; b_sign3 = 4'd1;
@(posedge clk_i);
shared_exps0 = 8'd132;
shared_exps1 = 8'd125;
a_mant0 = 8'd32; a_mant1 = 8'd184; a_mant2 = 8'd115; a_mant3 = 8'd235;
b_mant0 = 8'd127; b_mant1 = 8'd20; b_mant2 = 8'd80; b_mant3 = 8'd201;
a_exp0 = 10'd506; a_exp1 = 10'd752; a_exp2 = 10'd639; a_exp3 = 10'd565;
b_exp0 = 10'd418; b_exp1 = 10'd388; b_exp2 = 10'd814; b_exp3 = 10'd789;
a_sign0 = 4'd0; a_sign1 = 4'd14; a_sign2 = 4'd15; a_sign3 = 4'd8;
b_sign0 = 4'd2; b_sign1 = 4'd4; b_sign2 = 4'd4; b_sign3 = 4'd6;
@(posedge clk_i);
a_mant0 = 8'd76; a_mant1 = 8'd146; a_mant2 = 8'd200; a_mant3 = 8'd255;
b_mant0 = 8'd6; b_mant1 = 8'd48; b_mant2 = 8'd174; b_mant3 = 8'd191;
a_exp0 = 10'd873; a_exp1 = 10'd947; a_exp2 = 10'd426; a_exp3 = 10'd642;
b_exp0 = 10'd711; b_exp1 = 10'd549; b_exp2 = 10'd763; b_exp3 = 10'd44;
a_sign0 = 4'd15; a_sign1 = 4'd12; a_sign2 = 4'd1; a_sign3 = 4'd7;
b_sign0 = 4'd13; b_sign1 = 4'd13; b_sign2 = 4'd12; b_sign3 = 4'd13;
@(posedge clk_i);
a_mant0 = 8'd217; a_mant1 = 8'd217; a_mant2 = 8'd183; a_mant3 = 8'd171;
b_mant0 = 8'd207; b_mant1 = 8'd207; b_mant2 = 8'd121; b_mant3 = 8'd195;
a_exp0 = 10'd881; a_exp1 = 10'd387; a_exp2 = 10'd164; a_exp3 = 10'd315;
b_exp0 = 10'd469; b_exp1 = 10'd575; b_exp2 = 10'd350; b_exp3 = 10'd774;
a_sign0 = 4'd8; a_sign1 = 4'd1; a_sign2 = 4'd14; a_sign3 = 4'd3;
b_sign0 = 4'd15; b_sign1 = 4'd4; b_sign2 = 4'd2; b_sign3 = 4'd6;
@(posedge clk_i);
a_mant0 = 8'd143; a_mant1 = 8'd136; a_mant2 = 8'd178; a_mant3 = 8'd228;
b_mant0 = 8'd133; b_mant1 = 8'd97; b_mant2 = 8'd6; b_mant3 = 8'd37;
a_exp0 = 10'd515; a_exp1 = 10'd341; a_exp2 = 10'd43; a_exp3 = 10'd647;
b_exp0 = 10'd380; b_exp1 = 10'd349; b_exp2 = 10'd384; b_exp3 = 10'd886;
a_sign0 = 4'd4; a_sign1 = 4'd1; a_sign2 = 4'd1; a_sign3 = 4'd15;
b_sign0 = 4'd4; b_sign1 = 4'd12; b_sign2 = 4'd9; b_sign3 = 4'd13;
@(posedge clk_i);
a_mant0 = 8'd56; a_mant1 = 8'd194; a_mant2 = 8'd137; a_mant3 = 8'd57;
b_mant0 = 8'd185; b_mant1 = 8'd142; b_mant2 = 8'd194; b_mant3 = 8'd160;
a_exp0 = 10'd96; a_exp1 = 10'd869; a_exp2 = 10'd657; a_exp3 = 10'd977;
b_exp0 = 10'd1020; b_exp1 = 10'd462; b_exp2 = 10'd1023; b_exp3 = 10'd566;
a_sign0 = 4'd1; a_sign1 = 4'd8; a_sign2 = 4'd1; a_sign3 = 4'd12;
b_sign0 = 4'd13; b_sign1 = 4'd16; b_sign2 = 4'd0; b_sign3 = 4'd6;
@(posedge clk_i);
a_mant0 = 8'd200; a_mant1 = 8'd83; a_mant2 = 8'd99; a_mant3 = 8'd243;
b_mant0 = 8'd42; b_mant1 = 8'd195; b_mant2 = 8'd32; b_mant3 = 8'd70;
a_exp0 = 10'd126; a_exp1 = 10'd955; a_exp2 = 10'd10; a_exp3 = 10'd956;
b_exp0 = 10'd651; b_exp1 = 10'd876; b_exp2 = 10'd930; b_exp3 = 10'd423;
a_sign0 = 4'd10; a_sign1 = 4'd7; a_sign2 = 4'd3; a_sign3 = 4'd16;
b_sign0 = 4'd1; b_sign1 = 4'd3; b_sign2 = 4'd15; b_sign3 = 4'd7;
@(posedge clk_i);
a_mant0 = 8'd51; a_mant1 = 8'd2; a_mant2 = 8'd12; a_mant3 = 8'd213;
b_mant0 = 8'd240; b_mant1 = 8'd75; b_mant2 = 8'd240; b_mant3 = 8'd237;
a_exp0 = 10'd579; a_exp1 = 10'd941; a_exp2 = 10'd707; a_exp3 = 10'd249;
b_exp0 = 10'd433; b_exp1 = 10'd777; b_exp2 = 10'd1008; b_exp3 = 10'd857;
a_sign0 = 4'd16; a_sign1 = 4'd7; a_sign2 = 4'd4; a_sign3 = 4'd7;
b_sign0 = 4'd10; b_sign1 = 4'd9; b_sign2 = 4'd5; b_sign3 = 4'd8;
@(posedge clk_i);
a_mant0 = 8'd193; a_mant1 = 8'd10; a_mant2 = 8'd86; a_mant3 = 8'd63;
b_mant0 = 8'd245; b_mant1 = 8'd145; b_mant2 = 8'd135; b_mant3 = 8'd240;
a_exp0 = 10'd480; a_exp1 = 10'd471; a_exp2 = 10'd688; a_exp3 = 10'd144;
b_exp0 = 10'd329; b_exp1 = 10'd685; b_exp2 = 10'd659; b_exp3 = 10'd646;
a_sign0 = 4'd8; a_sign1 = 4'd16; a_sign2 = 4'd11; a_sign3 = 4'd10;
b_sign0 = 4'd2; b_sign1 = 4'd1; b_sign2 = 4'd0; b_sign3 = 4'd10;
@(posedge clk_i);
shared_exps0 = 8'd106;
shared_exps1 = 8'd144;
a_mant0 = 8'd40; a_mant1 = 8'd255; a_mant2 = 8'd240; a_mant3 = 8'd238;
b_mant0 = 8'd248; b_mant1 = 8'd102; b_mant2 = 8'd123; b_mant3 = 8'd162;
a_exp0 = 10'd314; a_exp1 = 10'd538; a_exp2 = 10'd91; a_exp3 = 10'd580;
b_exp0 = 10'd198; b_exp1 = 10'd764; b_exp2 = 10'd680; b_exp3 = 10'd657;
a_sign0 = 4'd12; a_sign1 = 4'd14; a_sign2 = 4'd14; a_sign3 = 4'd11;
b_sign0 = 4'd2; b_sign1 = 4'd1; b_sign2 = 4'd6; b_sign3 = 4'd15;
@(posedge clk_i);
a_mant0 = 8'd182; a_mant1 = 8'd17; a_mant2 = 8'd141; a_mant3 = 8'd161;
b_mant0 = 8'd206; b_mant1 = 8'd222; b_mant2 = 8'd8; b_mant3 = 8'd77;
a_exp0 = 10'd705; a_exp1 = 10'd403; a_exp2 = 10'd920; a_exp3 = 10'd416;
b_exp0 = 10'd636; b_exp1 = 10'd873; b_exp2 = 10'd847; b_exp3 = 10'd355;
a_sign0 = 4'd3; a_sign1 = 4'd8; a_sign2 = 4'd1; a_sign3 = 4'd2;
b_sign0 = 4'd4; b_sign1 = 4'd16; b_sign2 = 4'd3; b_sign3 = 4'd16;
@(posedge clk_i);
a_mant0 = 8'd14; a_mant1 = 8'd28; a_mant2 = 8'd245; a_mant3 = 8'd170;
b_mant0 = 8'd131; b_mant1 = 8'd97; b_mant2 = 8'd62; b_mant3 = 8'd94;
a_exp0 = 10'd85; a_exp1 = 10'd216; a_exp2 = 10'd830; a_exp3 = 10'd585;
b_exp0 = 10'd224; b_exp1 = 10'd882; b_exp2 = 10'd916; b_exp3 = 10'd162;
a_sign0 = 4'd5; a_sign1 = 4'd6; a_sign2 = 4'd13; a_sign3 = 4'd9;
b_sign0 = 4'd11; b_sign1 = 4'd5; b_sign2 = 4'd9; b_sign3 = 4'd9;
@(posedge clk_i);
a_mant0 = 8'd227; a_mant1 = 8'd46; a_mant2 = 8'd51; a_mant3 = 8'd9;
b_mant0 = 8'd196; b_mant1 = 8'd177; b_mant2 = 8'd227; b_mant3 = 8'd28;
a_exp0 = 10'd718; a_exp1 = 10'd204; a_exp2 = 10'd894; a_exp3 = 10'd553;
b_exp0 = 10'd335; b_exp1 = 10'd710; b_exp2 = 10'd894; b_exp3 = 10'd992;
a_sign0 = 4'd15; a_sign1 = 4'd16; a_sign2 = 4'd16; a_sign3 = 4'd9;
b_sign0 = 4'd13; b_sign1 = 4'd0; b_sign2 = 4'd14; b_sign3 = 4'd9;
@(posedge clk_i);
a_mant0 = 8'd117; a_mant1 = 8'd153; a_mant2 = 8'd43; a_mant3 = 8'd216;
b_mant0 = 8'd187; b_mant1 = 8'd147; b_mant2 = 8'd187; b_mant3 = 8'd212;
a_exp0 = 10'd574; a_exp1 = 10'd729; a_exp2 = 10'd479; a_exp3 = 10'd168;
b_exp0 = 10'd201; b_exp1 = 10'd769; b_exp2 = 10'd301; b_exp3 = 10'd403;
a_sign0 = 4'd2; a_sign1 = 4'd11; a_sign2 = 4'd4; a_sign3 = 4'd13;
b_sign0 = 4'd15; b_sign1 = 4'd15; b_sign2 = 4'd1; b_sign3 = 4'd4;
@(posedge clk_i);
a_mant0 = 8'd190; a_mant1 = 8'd213; a_mant2 = 8'd142; a_mant3 = 8'd179;
b_mant0 = 8'd89; b_mant1 = 8'd215; b_mant2 = 8'd94; b_mant3 = 8'd9;
a_exp0 = 10'd81; a_exp1 = 10'd661; a_exp2 = 10'd509; a_exp3 = 10'd178;
b_exp0 = 10'd977; b_exp1 = 10'd859; b_exp2 = 10'd350; b_exp3 = 10'd309;
a_sign0 = 4'd12; a_sign1 = 4'd5; a_sign2 = 4'd12; a_sign3 = 4'd14;
b_sign0 = 4'd3; b_sign1 = 4'd7; b_sign2 = 4'd7; b_sign3 = 4'd0;
@(posedge clk_i);
a_mant0 = 8'd208; a_mant1 = 8'd0; a_mant2 = 8'd123; a_mant3 = 8'd41;
b_mant0 = 8'd167; b_mant1 = 8'd85; b_mant2 = 8'd212; b_mant3 = 8'd2;
a_exp0 = 10'd641; a_exp1 = 10'd278; a_exp2 = 10'd327; a_exp3 = 10'd69;
b_exp0 = 10'd286; b_exp1 = 10'd317; b_exp2 = 10'd924; b_exp3 = 10'd558;
a_sign0 = 4'd2; a_sign1 = 4'd14; a_sign2 = 4'd12; a_sign3 = 4'd7;
b_sign0 = 4'd12; b_sign1 = 4'd11; b_sign2 = 4'd4; b_sign3 = 4'd5;
@(posedge clk_i);
a_mant0 = 8'd196; a_mant1 = 8'd141; a_mant2 = 8'd62; a_mant3 = 8'd55;
b_mant0 = 8'd49; b_mant1 = 8'd76; b_mant2 = 8'd166; b_mant3 = 8'd156;
a_exp0 = 10'd350; a_exp1 = 10'd279; a_exp2 = 10'd801; a_exp3 = 10'd653;
b_exp0 = 10'd823; b_exp1 = 10'd497; b_exp2 = 10'd309; b_exp3 = 10'd805;
a_sign0 = 4'd3; a_sign1 = 4'd6; a_sign2 = 4'd8; a_sign3 = 4'd11;
b_sign0 = 4'd6; b_sign1 = 4'd3; b_sign2 = 4'd1; b_sign3 = 4'd0;
@(posedge clk_i);
shared_exps0 = 8'd143;
shared_exps1 = 8'd112;
rstn = 0;
@(posedge clk_i);
rstn = 1;
a_mant0 = 8'd22; a_mant1 = 8'd25; a_mant2 = 8'd208; a_mant3 = 8'd74;
b_mant0 = 8'd44; b_mant1 = 8'd1; b_mant2 = 8'd186; b_mant3 = 8'd133;
a_exp0 = 10'd693; a_exp1 = 10'd317; a_exp2 = 10'd453; a_exp3 = 10'd672;
b_exp0 = 10'd316; b_exp1 = 10'd1000; b_exp2 = 10'd675; b_exp3 = 10'd375;
a_sign0 = 4'd14; a_sign1 = 4'd9; a_sign2 = 4'd2; a_sign3 = 4'd9;
b_sign0 = 4'd12; b_sign1 = 4'd2; b_sign2 = 4'd16; b_sign3 = 4'd4;
@(posedge clk_i);
a_mant0 = 8'd170; a_mant1 = 8'd10; a_mant2 = 8'd118; a_mant3 = 8'd86;
b_mant0 = 8'd80; b_mant1 = 8'd97; b_mant2 = 8'd3; b_mant3 = 8'd3;
a_exp0 = 10'd743; a_exp1 = 10'd120; a_exp2 = 10'd513; a_exp3 = 10'd683;
b_exp0 = 10'd176; b_exp1 = 10'd962; b_exp2 = 10'd211; b_exp3 = 10'd633;
a_sign0 = 4'd12; a_sign1 = 4'd11; a_sign2 = 4'd14; a_sign3 = 4'd13;
b_sign0 = 4'd2; b_sign1 = 4'd5; b_sign2 = 4'd13; b_sign3 = 4'd15;
@(posedge clk_i);
a_mant0 = 8'd77; a_mant1 = 8'd196; a_mant2 = 8'd184; a_mant3 = 8'd226;
b_mant0 = 8'd227; b_mant1 = 8'd218; b_mant2 = 8'd191; b_mant3 = 8'd80;
a_exp0 = 10'd527; a_exp1 = 10'd21; a_exp2 = 10'd577; a_exp3 = 10'd281;
b_exp0 = 10'd386; b_exp1 = 10'd390; b_exp2 = 10'd20; b_exp3 = 10'd943;
a_sign0 = 4'd15; a_sign1 = 4'd15; a_sign2 = 4'd13; a_sign3 = 4'd1;
b_sign0 = 4'd4; b_sign1 = 4'd6; b_sign2 = 4'd13; b_sign3 = 4'd12;
@(posedge clk_i);
a_mant0 = 8'd83; a_mant1 = 8'd62; a_mant2 = 8'd240; a_mant3 = 8'd23;
b_mant0 = 8'd68; b_mant1 = 8'd208; b_mant2 = 8'd9; b_mant3 = 8'd214;
a_exp0 = 10'd407; a_exp1 = 10'd627; a_exp2 = 10'd955; a_exp3 = 10'd569;
b_exp0 = 10'd509; b_exp1 = 10'd328; b_exp2 = 10'd897; b_exp3 = 10'd48;
a_sign0 = 4'd5; a_sign1 = 4'd3; a_sign2 = 4'd4; a_sign3 = 4'd14;
b_sign0 = 4'd14; b_sign1 = 4'd13; b_sign2 = 4'd14; b_sign3 = 4'd2;
@(posedge clk_i);
a_mant0 = 8'd49; a_mant1 = 8'd212; a_mant2 = 8'd7; a_mant3 = 8'd129;
b_mant0 = 8'd131; b_mant1 = 8'd133; b_mant2 = 8'd223; b_mant3 = 8'd192;
a_exp0 = 10'd1004; a_exp1 = 10'd395; a_exp2 = 10'd963; a_exp3 = 10'd445;
b_exp0 = 10'd339; b_exp1 = 10'd633; b_exp2 = 10'd850; b_exp3 = 10'd879;
a_sign0 = 4'd6; a_sign1 = 4'd9; a_sign2 = 4'd13; a_sign3 = 4'd0;
b_sign0 = 4'd0; b_sign1 = 4'd9; b_sign2 = 4'd4; b_sign3 = 4'd6;
@(posedge clk_i);
a_mant0 = 8'd155; a_mant1 = 8'd67; a_mant2 = 8'd224; a_mant3 = 8'd31;
b_mant0 = 8'd161; b_mant1 = 8'd250; b_mant2 = 8'd168; b_mant3 = 8'd30;
a_exp0 = 10'd1022; a_exp1 = 10'd435; a_exp2 = 10'd363; a_exp3 = 10'd990;
b_exp0 = 10'd626; b_exp1 = 10'd806; b_exp2 = 10'd149; b_exp3 = 10'd391;
a_sign0 = 4'd14; a_sign1 = 4'd14; a_sign2 = 4'd11; a_sign3 = 4'd13;
b_sign0 = 4'd14; b_sign1 = 4'd4; b_sign2 = 4'd16; b_sign3 = 4'd15;
@(posedge clk_i);
a_mant0 = 8'd1; a_mant1 = 8'd83; a_mant2 = 8'd250; a_mant3 = 8'd75;
b_mant0 = 8'd19; b_mant1 = 8'd148; b_mant2 = 8'd185; b_mant3 = 8'd103;
a_exp0 = 10'd911; a_exp1 = 10'd831; a_exp2 = 10'd607; a_exp3 = 10'd594;
b_exp0 = 10'd873; b_exp1 = 10'd580; b_exp2 = 10'd597; b_exp3 = 10'd688;
a_sign0 = 4'd2; a_sign1 = 4'd13; a_sign2 = 4'd9; a_sign3 = 4'd8;
b_sign0 = 4'd2; b_sign1 = 4'd5; b_sign2 = 4'd11; b_sign3 = 4'd9;
@(posedge clk_i);
shared_exps0 = 8'd121;
shared_exps1 = 8'd151;
a_mant0 = 8'd97; a_mant1 = 8'd194; a_mant2 = 8'd43; a_mant3 = 8'd102;
b_mant0 = 8'd168; b_mant1 = 8'd11; b_mant2 = 8'd185; b_mant3 = 8'd18;
a_exp0 = 10'd182; a_exp1 = 10'd274; a_exp2 = 10'd347; a_exp3 = 10'd592;
b_exp0 = 10'd162; b_exp1 = 10'd470; b_exp2 = 10'd902; b_exp3 = 10'd260;
a_sign0 = 4'd0; a_sign1 = 4'd13; a_sign2 = 4'd16; a_sign3 = 4'd11;
b_sign0 = 4'd13; b_sign1 = 4'd4; b_sign2 = 4'd14; b_sign3 = 4'd11;
@(posedge clk_i);
a_mant0 = 8'd184; a_mant1 = 8'd131; a_mant2 = 8'd189; a_mant3 = 8'd72;
b_mant0 = 8'd101; b_mant1 = 8'd49; b_mant2 = 8'd177; b_mant3 = 8'd13;
a_exp0 = 10'd203; a_exp1 = 10'd0; a_exp2 = 10'd88; a_exp3 = 10'd414;
b_exp0 = 10'd289; b_exp1 = 10'd387; b_exp2 = 10'd625; b_exp3 = 10'd990;
a_sign0 = 4'd4; a_sign1 = 4'd11; a_sign2 = 4'd6; a_sign3 = 4'd6;
b_sign0 = 4'd7; b_sign1 = 4'd8; b_sign2 = 4'd7; b_sign3 = 4'd11;
@(posedge clk_i);
a_mant0 = 8'd99; a_mant1 = 8'd71; a_mant2 = 8'd46; a_mant3 = 8'd113;
b_mant0 = 8'd106; b_mant1 = 8'd31; b_mant2 = 8'd53; b_mant3 = 8'd25;
a_exp0 = 10'd249; a_exp1 = 10'd932; a_exp2 = 10'd905; a_exp3 = 10'd990;
b_exp0 = 10'd462; b_exp1 = 10'd799; b_exp2 = 10'd354; b_exp3 = 10'd677;
a_sign0 = 4'd9; a_sign1 = 4'd8; a_sign2 = 4'd1; a_sign3 = 4'd14;
b_sign0 = 4'd2; b_sign1 = 4'd10; b_sign2 = 4'd6; b_sign3 = 4'd12;
@(posedge clk_i);
a_mant0 = 8'd118; a_mant1 = 8'd206; a_mant2 = 8'd48; a_mant3 = 8'd143;
b_mant0 = 8'd87; b_mant1 = 8'd83; b_mant2 = 8'd55; b_mant3 = 8'd154;
a_exp0 = 10'd735; a_exp1 = 10'd186; a_exp2 = 10'd325; a_exp3 = 10'd135;
b_exp0 = 10'd631; b_exp1 = 10'd57; b_exp2 = 10'd817; b_exp3 = 10'd2;
a_sign0 = 4'd14; a_sign1 = 4'd6; a_sign2 = 4'd1; a_sign3 = 4'd15;
b_sign0 = 4'd4; b_sign1 = 4'd2; b_sign2 = 4'd7; b_sign3 = 4'd3;
@(posedge clk_i);
a_mant0 = 8'd203; a_mant1 = 8'd106; a_mant2 = 8'd176; a_mant3 = 8'd183;
b_mant0 = 8'd174; b_mant1 = 8'd57; b_mant2 = 8'd216; b_mant3 = 8'd167;
a_exp0 = 10'd754; a_exp1 = 10'd782; a_exp2 = 10'd43; a_exp3 = 10'd129;
b_exp0 = 10'd112; b_exp1 = 10'd750; b_exp2 = 10'd365; b_exp3 = 10'd440;
a_sign0 = 4'd3; a_sign1 = 4'd7; a_sign2 = 4'd4; a_sign3 = 4'd15;
b_sign0 = 4'd8; b_sign1 = 4'd16; b_sign2 = 4'd5; b_sign3 = 4'd1;
@(posedge clk_i);
a_mant0 = 8'd95; a_mant1 = 8'd251; a_mant2 = 8'd193; a_mant3 = 8'd41;
b_mant0 = 8'd20; b_mant1 = 8'd226; b_mant2 = 8'd48; b_mant3 = 8'd234;
a_exp0 = 10'd638; a_exp1 = 10'd622; a_exp2 = 10'd55; a_exp3 = 10'd985;
b_exp0 = 10'd314; b_exp1 = 10'd454; b_exp2 = 10'd603; b_exp3 = 10'd907;
a_sign0 = 4'd13; a_sign1 = 4'd0; a_sign2 = 4'd6; a_sign3 = 4'd16;
b_sign0 = 4'd10; b_sign1 = 4'd10; b_sign2 = 4'd12; b_sign3 = 4'd15;
@(posedge clk_i);
a_mant0 = 8'd8; a_mant1 = 8'd98; a_mant2 = 8'd128; a_mant3 = 8'd74;
b_mant0 = 8'd47; b_mant1 = 8'd220; b_mant2 = 8'd108; b_mant3 = 8'd5;
a_exp0 = 10'd914; a_exp1 = 10'd305; a_exp2 = 10'd118; a_exp3 = 10'd974;
b_exp0 = 10'd555; b_exp1 = 10'd969; b_exp2 = 10'd560; b_exp3 = 10'd359;
a_sign0 = 4'd14; a_sign1 = 4'd0; a_sign2 = 4'd7; a_sign3 = 4'd13;
b_sign0 = 4'd3; b_sign1 = 4'd3; b_sign2 = 4'd14; b_sign3 = 4'd4;
@(posedge clk_i);
a_mant0 = 8'd113; a_mant1 = 8'd50; a_mant2 = 8'd108; a_mant3 = 8'd131;
b_mant0 = 8'd163; b_mant1 = 8'd60; b_mant2 = 8'd57; b_mant3 = 8'd35;
a_exp0 = 10'd347; a_exp1 = 10'd389; a_exp2 = 10'd449; a_exp3 = 10'd16;
b_exp0 = 10'd865; b_exp1 = 10'd906; b_exp2 = 10'd501; b_exp3 = 10'd683;
a_sign0 = 4'd8; a_sign1 = 4'd11; a_sign2 = 4'd5; a_sign3 = 4'd15;
b_sign0 = 4'd16; b_sign1 = 4'd10; b_sign2 = 4'd12; b_sign3 = 4'd0;
@(posedge clk_i);
shared_exps0 = 8'd124;
shared_exps1 = 8'd132;
a_mant0 = 8'd140; a_mant1 = 8'd34; a_mant2 = 8'd67; a_mant3 = 8'd119;
b_mant0 = 8'd178; b_mant1 = 8'd114; b_mant2 = 8'd99; b_mant3 = 8'd114;
a_exp0 = 10'd262; a_exp1 = 10'd9; a_exp2 = 10'd622; a_exp3 = 10'd584;
b_exp0 = 10'd773; b_exp1 = 10'd502; b_exp2 = 10'd440; b_exp3 = 10'd791;
a_sign0 = 4'd11; a_sign1 = 4'd1; a_sign2 = 4'd5; a_sign3 = 4'd15;
b_sign0 = 4'd0; b_sign1 = 4'd14; b_sign2 = 4'd11; b_sign3 = 4'd10;
@(posedge clk_i);
a_mant0 = 8'd224; a_mant1 = 8'd17; a_mant2 = 8'd127; a_mant3 = 8'd227;
b_mant0 = 8'd169; b_mant1 = 8'd51; b_mant2 = 8'd211; b_mant3 = 8'd3;
a_exp0 = 10'd471; a_exp1 = 10'd271; a_exp2 = 10'd730; a_exp3 = 10'd566;
b_exp0 = 10'd776; b_exp1 = 10'd41; b_exp2 = 10'd782; b_exp3 = 10'd121;
a_sign0 = 4'd10; a_sign1 = 4'd6; a_sign2 = 4'd5; a_sign3 = 4'd5;
b_sign0 = 4'd12; b_sign1 = 4'd7; b_sign2 = 4'd2; b_sign3 = 4'd1;
@(posedge clk_i);
a_mant0 = 8'd231; a_mant1 = 8'd153; a_mant2 = 8'd186; a_mant3 = 8'd8;
b_mant0 = 8'd253; b_mant1 = 8'd9; b_mant2 = 8'd146; b_mant3 = 8'd91;
a_exp0 = 10'd985; a_exp1 = 10'd680; a_exp2 = 10'd7; a_exp3 = 10'd591;
b_exp0 = 10'd270; b_exp1 = 10'd753; b_exp2 = 10'd177; b_exp3 = 10'd352;
a_sign0 = 4'd15; a_sign1 = 4'd4; a_sign2 = 4'd8; a_sign3 = 4'd6;
b_sign0 = 4'd5; b_sign1 = 4'd1; b_sign2 = 4'd4; b_sign3 = 4'd10;
@(posedge clk_i);
a_mant0 = 8'd156; a_mant1 = 8'd71; a_mant2 = 8'd64; a_mant3 = 8'd0;
b_mant0 = 8'd178; b_mant1 = 8'd242; b_mant2 = 8'd242; b_mant3 = 8'd18;
a_exp0 = 10'd509; a_exp1 = 10'd893; a_exp2 = 10'd859; a_exp3 = 10'd88;
b_exp0 = 10'd243; b_exp1 = 10'd1007; b_exp2 = 10'd435; b_exp3 = 10'd866;
a_sign0 = 4'd9; a_sign1 = 4'd5; a_sign2 = 4'd4; a_sign3 = 4'd0;
b_sign0 = 4'd8; b_sign1 = 4'd11; b_sign2 = 4'd3; b_sign3 = 4'd8;
@(posedge clk_i);
a_mant0 = 8'd20; a_mant1 = 8'd156; a_mant2 = 8'd101; a_mant3 = 8'd169;
b_mant0 = 8'd168; b_mant1 = 8'd134; b_mant2 = 8'd21; b_mant3 = 8'd32;
a_exp0 = 10'd206; a_exp1 = 10'd328; a_exp2 = 10'd519; a_exp3 = 10'd56;
b_exp0 = 10'd586; b_exp1 = 10'd196; b_exp2 = 10'd145; b_exp3 = 10'd310;
a_sign0 = 4'd4; a_sign1 = 4'd6; a_sign2 = 4'd10; a_sign3 = 4'd9;
b_sign0 = 4'd11; b_sign1 = 4'd1; b_sign2 = 4'd3; b_sign3 = 4'd0;
@(posedge clk_i);
a_mant0 = 8'd58; a_mant1 = 8'd65; a_mant2 = 8'd41; a_mant3 = 8'd109;
b_mant0 = 8'd35; b_mant1 = 8'd31; b_mant2 = 8'd123; b_mant3 = 8'd88;
a_exp0 = 10'd147; a_exp1 = 10'd233; a_exp2 = 10'd441; a_exp3 = 10'd541;
b_exp0 = 10'd396; b_exp1 = 10'd768; b_exp2 = 10'd789; b_exp3 = 10'd973;
a_sign0 = 4'd9; a_sign1 = 4'd0; a_sign2 = 4'd13; a_sign3 = 4'd12;
b_sign0 = 4'd5; b_sign1 = 4'd4; b_sign2 = 4'd16; b_sign3 = 4'd13;
@(posedge clk_i);
a_mant0 = 8'd173; a_mant1 = 8'd103; a_mant2 = 8'd218; a_mant3 = 8'd144;
b_mant0 = 8'd17; b_mant1 = 8'd171; b_mant2 = 8'd200; b_mant3 = 8'd241;
a_exp0 = 10'd276; a_exp1 = 10'd980; a_exp2 = 10'd248; a_exp3 = 10'd688;
b_exp0 = 10'd14; b_exp1 = 10'd942; b_exp2 = 10'd909; b_exp3 = 10'd564;
a_sign0 = 4'd10; a_sign1 = 4'd9; a_sign2 = 4'd0; a_sign3 = 4'd15;
b_sign0 = 4'd13; b_sign1 = 4'd11; b_sign2 = 4'd7; b_sign3 = 4'd1;
@(posedge clk_i);
a_mant0 = 8'd143; a_mant1 = 8'd209; a_mant2 = 8'd111; a_mant3 = 8'd7;
b_mant0 = 8'd161; b_mant1 = 8'd202; b_mant2 = 8'd181; b_mant3 = 8'd218;
a_exp0 = 10'd984; a_exp1 = 10'd91; a_exp2 = 10'd996; a_exp3 = 10'd744;
b_exp0 = 10'd856; b_exp1 = 10'd429; b_exp2 = 10'd243; b_exp3 = 10'd723;
a_sign0 = 4'd8; a_sign1 = 4'd14; a_sign2 = 4'd2; a_sign3 = 4'd13;
b_sign0 = 4'd16; b_sign1 = 4'd0; b_sign2 = 4'd15; b_sign3 = 4'd15;
@(posedge clk_i);
shared_exps0 = 8'd117;
shared_exps1 = 8'd118;
a_mant0 = 8'd198; a_mant1 = 8'd64; a_mant2 = 8'd89; a_mant3 = 8'd208;
b_mant0 = 8'd174; b_mant1 = 8'd199; b_mant2 = 8'd64; b_mant3 = 8'd3;
a_exp0 = 10'd180; a_exp1 = 10'd900; a_exp2 = 10'd484; a_exp3 = 10'd530;
b_exp0 = 10'd13; b_exp1 = 10'd513; b_exp2 = 10'd671; b_exp3 = 10'd899;
a_sign0 = 4'd0; a_sign1 = 4'd4; a_sign2 = 4'd10; a_sign3 = 4'd9;
b_sign0 = 4'd14; b_sign1 = 4'd14; b_sign2 = 4'd5; b_sign3 = 4'd2;
@(posedge clk_i);
a_mant0 = 8'd206; a_mant1 = 8'd234; a_mant2 = 8'd113; a_mant3 = 8'd215;
b_mant0 = 8'd121; b_mant1 = 8'd17; b_mant2 = 8'd244; b_mant3 = 8'd198;
a_exp0 = 10'd418; a_exp1 = 10'd104; a_exp2 = 10'd1018; a_exp3 = 10'd86;
b_exp0 = 10'd145; b_exp1 = 10'd160; b_exp2 = 10'd449; b_exp3 = 10'd363;
a_sign0 = 4'd9; a_sign1 = 4'd6; a_sign2 = 4'd1; a_sign3 = 4'd12;
b_sign0 = 4'd12; b_sign1 = 4'd9; b_sign2 = 4'd13; b_sign3 = 4'd16;
@(posedge clk_i);
a_mant0 = 8'd60; a_mant1 = 8'd108; a_mant2 = 8'd196; a_mant3 = 8'd12;
b_mant0 = 8'd179; b_mant1 = 8'd115; b_mant2 = 8'd153; b_mant3 = 8'd35;
a_exp0 = 10'd110; a_exp1 = 10'd1008; a_exp2 = 10'd324; a_exp3 = 10'd401;
b_exp0 = 10'd763; b_exp1 = 10'd721; b_exp2 = 10'd1002; b_exp3 = 10'd527;
a_sign0 = 4'd8; a_sign1 = 4'd3; a_sign2 = 4'd13; a_sign3 = 4'd9;
b_sign0 = 4'd15; b_sign1 = 4'd13; b_sign2 = 4'd13; b_sign3 = 4'd8;
@(posedge clk_i);
a_mant0 = 8'd215; a_mant1 = 8'd17; a_mant2 = 8'd123; a_mant3 = 8'd213;
b_mant0 = 8'd101; b_mant1 = 8'd72; b_mant2 = 8'd219; b_mant3 = 8'd49;
a_exp0 = 10'd560; a_exp1 = 10'd907; a_exp2 = 10'd84; a_exp3 = 10'd126;
b_exp0 = 10'd837; b_exp1 = 10'd893; b_exp2 = 10'd702; b_exp3 = 10'd661;
a_sign0 = 4'd3; a_sign1 = 4'd10; a_sign2 = 4'd2; a_sign3 = 4'd16;
b_sign0 = 4'd13; b_sign1 = 4'd9; b_sign2 = 4'd16; b_sign3 = 4'd15;
@(posedge clk_i);
a_mant0 = 8'd228; a_mant1 = 8'd201; a_mant2 = 8'd109; a_mant3 = 8'd71;
b_mant0 = 8'd118; b_mant1 = 8'd178; b_mant2 = 8'd0; b_mant3 = 8'd231;
a_exp0 = 10'd348; a_exp1 = 10'd751; a_exp2 = 10'd793; a_exp3 = 10'd200;
b_exp0 = 10'd407; b_exp1 = 10'd955; b_exp2 = 10'd648; b_exp3 = 10'd574;
a_sign0 = 4'd3; a_sign1 = 4'd2; a_sign2 = 4'd15; a_sign3 = 4'd10;
b_sign0 = 4'd9; b_sign1 = 4'd9; b_sign2 = 4'd9; b_sign3 = 4'd7;
@(posedge clk_i);
a_mant0 = 8'd18; a_mant1 = 8'd207; a_mant2 = 8'd144; a_mant3 = 8'd134;
b_mant0 = 8'd36; b_mant1 = 8'd201; b_mant2 = 8'd172; b_mant3 = 8'd73;
a_exp0 = 10'd895; a_exp1 = 10'd785; a_exp2 = 10'd750; a_exp3 = 10'd149;
b_exp0 = 10'd367; b_exp1 = 10'd59; b_exp2 = 10'd130; b_exp3 = 10'd675;
a_sign0 = 4'd16; a_sign1 = 4'd12; a_sign2 = 4'd14; a_sign3 = 4'd6;
b_sign0 = 4'd10; b_sign1 = 4'd11; b_sign2 = 4'd7; b_sign3 = 4'd2;
@(posedge clk_i);
a_mant0 = 8'd138; a_mant1 = 8'd69; a_mant2 = 8'd230; a_mant3 = 8'd67;
b_mant0 = 8'd226; b_mant1 = 8'd131; b_mant2 = 8'd48; b_mant3 = 8'd68;
a_exp0 = 10'd704; a_exp1 = 10'd700; a_exp2 = 10'd69; a_exp3 = 10'd694;
b_exp0 = 10'd316; b_exp1 = 10'd242; b_exp2 = 10'd371; b_exp3 = 10'd311;
a_sign0 = 4'd7; a_sign1 = 4'd0; a_sign2 = 4'd4; a_sign3 = 4'd14;
b_sign0 = 4'd11; b_sign1 = 4'd8; b_sign2 = 4'd3; b_sign3 = 4'd3;
@(posedge clk_i);
a_mant0 = 8'd118; a_mant1 = 8'd213; a_mant2 = 8'd149; a_mant3 = 8'd194;
b_mant0 = 8'd47; b_mant1 = 8'd153; b_mant2 = 8'd57; b_mant3 = 8'd61;
a_exp0 = 10'd636; a_exp1 = 10'd655; a_exp2 = 10'd816; a_exp3 = 10'd800;
b_exp0 = 10'd746; b_exp1 = 10'd259; b_exp2 = 10'd338; b_exp3 = 10'd417;
a_sign0 = 4'd13; a_sign1 = 4'd13; a_sign2 = 4'd15; a_sign3 = 4'd0;
b_sign0 = 4'd12; b_sign1 = 4'd10; b_sign2 = 4'd12; b_sign3 = 4'd6;
@(posedge clk_i);
shared_exps0 = 8'd124;
shared_exps1 = 8'd104;
rstn = 0;
@(posedge clk_i);
rstn = 1;
a_mant0 = 8'd120; a_mant1 = 8'd155; a_mant2 = 8'd89; a_mant3 = 8'd220;
b_mant0 = 8'd176; b_mant1 = 8'd172; b_mant2 = 8'd238; b_mant3 = 8'd24;
a_exp0 = 10'd375; a_exp1 = 10'd363; a_exp2 = 10'd551; a_exp3 = 10'd434;
b_exp0 = 10'd147; b_exp1 = 10'd299; b_exp2 = 10'd301; b_exp3 = 10'd414;
a_sign0 = 4'd16; a_sign1 = 4'd7; a_sign2 = 4'd10; a_sign3 = 4'd3;
b_sign0 = 4'd7; b_sign1 = 4'd6; b_sign2 = 4'd1; b_sign3 = 4'd11;
@(posedge clk_i);
a_mant0 = 8'd50; a_mant1 = 8'd124; a_mant2 = 8'd25; a_mant3 = 8'd142;
b_mant0 = 8'd177; b_mant1 = 8'd205; b_mant2 = 8'd105; b_mant3 = 8'd102;
a_exp0 = 10'd196; a_exp1 = 10'd843; a_exp2 = 10'd247; a_exp3 = 10'd990;
b_exp0 = 10'd589; b_exp1 = 10'd375; b_exp2 = 10'd162; b_exp3 = 10'd883;
a_sign0 = 4'd2; a_sign1 = 4'd1; a_sign2 = 4'd14; a_sign3 = 4'd8;
b_sign0 = 4'd16; b_sign1 = 4'd0; b_sign2 = 4'd8; b_sign3 = 4'd10;
@(posedge clk_i);
a_mant0 = 8'd205; a_mant1 = 8'd171; a_mant2 = 8'd242; a_mant3 = 8'd204;
b_mant0 = 8'd52; b_mant1 = 8'd254; b_mant2 = 8'd86; b_mant3 = 8'd150;
a_exp0 = 10'd270; a_exp1 = 10'd15; a_exp2 = 10'd726; a_exp3 = 10'd435;
b_exp0 = 10'd879; b_exp1 = 10'd695; b_exp2 = 10'd1000; b_exp3 = 10'd371;
a_sign0 = 4'd16; a_sign1 = 4'd5; a_sign2 = 4'd7; a_sign3 = 4'd8;
b_sign0 = 4'd10; b_sign1 = 4'd9; b_sign2 = 4'd6; b_sign3 = 4'd1;
@(posedge clk_i);
a_mant0 = 8'd44; a_mant1 = 8'd70; a_mant2 = 8'd114; a_mant3 = 8'd64;
b_mant0 = 8'd134; b_mant1 = 8'd88; b_mant2 = 8'd101; b_mant3 = 8'd175;
a_exp0 = 10'd588; a_exp1 = 10'd276; a_exp2 = 10'd93; a_exp3 = 10'd378;
b_exp0 = 10'd279; b_exp1 = 10'd544; b_exp2 = 10'd311; b_exp3 = 10'd917;
a_sign0 = 4'd7; a_sign1 = 4'd6; a_sign2 = 4'd4; a_sign3 = 4'd10;
b_sign0 = 4'd5; b_sign1 = 4'd3; b_sign2 = 4'd3; b_sign3 = 4'd0;
@(posedge clk_i);
a_mant0 = 8'd30; a_mant1 = 8'd253; a_mant2 = 8'd37; a_mant3 = 8'd78;
b_mant0 = 8'd100; b_mant1 = 8'd196; b_mant2 = 8'd177; b_mant3 = 8'd222;
a_exp0 = 10'd418; a_exp1 = 10'd30; a_exp2 = 10'd25; a_exp3 = 10'd364;
b_exp0 = 10'd708; b_exp1 = 10'd602; b_exp2 = 10'd220; b_exp3 = 10'd1015;
a_sign0 = 4'd12; a_sign1 = 4'd7; a_sign2 = 4'd11; a_sign3 = 4'd12;
b_sign0 = 4'd13; b_sign1 = 4'd16; b_sign2 = 4'd0; b_sign3 = 4'd10;
@(posedge clk_i);
a_mant0 = 8'd184; a_mant1 = 8'd201; a_mant2 = 8'd129; a_mant3 = 8'd118;
b_mant0 = 8'd194; b_mant1 = 8'd97; b_mant2 = 8'd98; b_mant3 = 8'd82;
a_exp0 = 10'd613; a_exp1 = 10'd1007; a_exp2 = 10'd648; a_exp3 = 10'd804;
b_exp0 = 10'd594; b_exp1 = 10'd571; b_exp2 = 10'd241; b_exp3 = 10'd353;
a_sign0 = 4'd13; a_sign1 = 4'd2; a_sign2 = 4'd8; a_sign3 = 4'd5;
b_sign0 = 4'd16; b_sign1 = 4'd8; b_sign2 = 4'd0; b_sign3 = 4'd7;
@(posedge clk_i);
a_mant0 = 8'd244; a_mant1 = 8'd108; a_mant2 = 8'd135; a_mant3 = 8'd77;
b_mant0 = 8'd249; b_mant1 = 8'd118; b_mant2 = 8'd113; b_mant3 = 8'd106;
a_exp0 = 10'd589; a_exp1 = 10'd339; a_exp2 = 10'd496; a_exp3 = 10'd737;
b_exp0 = 10'd503; b_exp1 = 10'd313; b_exp2 = 10'd773; b_exp3 = 10'd222;
a_sign0 = 4'd2; a_sign1 = 4'd7; a_sign2 = 4'd8; a_sign3 = 4'd12;
b_sign0 = 4'd15; b_sign1 = 4'd10; b_sign2 = 4'd10; b_sign3 = 4'd4;
@(posedge clk_i);
shared_exps0 = 8'd137;
shared_exps1 = 8'd133;
a_mant0 = 8'd132; a_mant1 = 8'd27; a_mant2 = 8'd131; a_mant3 = 8'd216;
b_mant0 = 8'd189; b_mant1 = 8'd215; b_mant2 = 8'd72; b_mant3 = 8'd108;
a_exp0 = 10'd161; a_exp1 = 10'd830; a_exp2 = 10'd587; a_exp3 = 10'd719;
b_exp0 = 10'd290; b_exp1 = 10'd594; b_exp2 = 10'd432; b_exp3 = 10'd472;
a_sign0 = 4'd15; a_sign1 = 4'd13; a_sign2 = 4'd11; a_sign3 = 4'd16;
b_sign0 = 4'd13; b_sign1 = 4'd6; b_sign2 = 4'd11; b_sign3 = 4'd6;
@(posedge clk_i);
a_mant0 = 8'd36; a_mant1 = 8'd74; a_mant2 = 8'd43; a_mant3 = 8'd64;
b_mant0 = 8'd200; b_mant1 = 8'd24; b_mant2 = 8'd136; b_mant3 = 8'd231;
a_exp0 = 10'd891; a_exp1 = 10'd692; a_exp2 = 10'd333; a_exp3 = 10'd791;
b_exp0 = 10'd168; b_exp1 = 10'd83; b_exp2 = 10'd525; b_exp3 = 10'd100;
a_sign0 = 4'd1; a_sign1 = 4'd6; a_sign2 = 4'd2; a_sign3 = 4'd3;
b_sign0 = 4'd8; b_sign1 = 4'd6; b_sign2 = 4'd12; b_sign3 = 4'd4;
@(posedge clk_i);
a_mant0 = 8'd125; a_mant1 = 8'd149; a_mant2 = 8'd1; a_mant3 = 8'd94;
b_mant0 = 8'd167; b_mant1 = 8'd26; b_mant2 = 8'd217; b_mant3 = 8'd36;
a_exp0 = 10'd839; a_exp1 = 10'd872; a_exp2 = 10'd284; a_exp3 = 10'd50;
b_exp0 = 10'd117; b_exp1 = 10'd606; b_exp2 = 10'd364; b_exp3 = 10'd720;
a_sign0 = 4'd4; a_sign1 = 4'd12; a_sign2 = 4'd12; a_sign3 = 4'd2;
b_sign0 = 4'd9; b_sign1 = 4'd8; b_sign2 = 4'd15; b_sign3 = 4'd3;
@(posedge clk_i);
a_mant0 = 8'd73; a_mant1 = 8'd139; a_mant2 = 8'd157; a_mant3 = 8'd20;
b_mant0 = 8'd139; b_mant1 = 8'd38; b_mant2 = 8'd69; b_mant3 = 8'd120;
a_exp0 = 10'd625; a_exp1 = 10'd967; a_exp2 = 10'd633; a_exp3 = 10'd354;
b_exp0 = 10'd1011; b_exp1 = 10'd549; b_exp2 = 10'd439; b_exp3 = 10'd32;
a_sign0 = 4'd8; a_sign1 = 4'd2; a_sign2 = 4'd0; a_sign3 = 4'd16;
b_sign0 = 4'd14; b_sign1 = 4'd4; b_sign2 = 4'd14; b_sign3 = 4'd0;
@(posedge clk_i);
a_mant0 = 8'd40; a_mant1 = 8'd168; a_mant2 = 8'd254; a_mant3 = 8'd108;
b_mant0 = 8'd158; b_mant1 = 8'd95; b_mant2 = 8'd22; b_mant3 = 8'd192;
a_exp0 = 10'd998; a_exp1 = 10'd239; a_exp2 = 10'd575; a_exp3 = 10'd951;
b_exp0 = 10'd642; b_exp1 = 10'd865; b_exp2 = 10'd406; b_exp3 = 10'd344;
a_sign0 = 4'd4; a_sign1 = 4'd13; a_sign2 = 4'd3; a_sign3 = 4'd6;
b_sign0 = 4'd14; b_sign1 = 4'd5; b_sign2 = 4'd12; b_sign3 = 4'd2;
@(posedge clk_i);
a_mant0 = 8'd7; a_mant1 = 8'd59; a_mant2 = 8'd241; a_mant3 = 8'd253;
b_mant0 = 8'd178; b_mant1 = 8'd206; b_mant2 = 8'd93; b_mant3 = 8'd133;
a_exp0 = 10'd184; a_exp1 = 10'd883; a_exp2 = 10'd301; a_exp3 = 10'd607;
b_exp0 = 10'd553; b_exp1 = 10'd312; b_exp2 = 10'd367; b_exp3 = 10'd912;
a_sign0 = 4'd6; a_sign1 = 4'd12; a_sign2 = 4'd4; a_sign3 = 4'd11;
b_sign0 = 4'd12; b_sign1 = 4'd5; b_sign2 = 4'd13; b_sign3 = 4'd2;
@(posedge clk_i);
a_mant0 = 8'd155; a_mant1 = 8'd179; a_mant2 = 8'd197; a_mant3 = 8'd40;
b_mant0 = 8'd12; b_mant1 = 8'd142; b_mant2 = 8'd59; b_mant3 = 8'd219;
a_exp0 = 10'd367; a_exp1 = 10'd872; a_exp2 = 10'd405; a_exp3 = 10'd834;
b_exp0 = 10'd689; b_exp1 = 10'd129; b_exp2 = 10'd373; b_exp3 = 10'd964;
a_sign0 = 4'd1; a_sign1 = 4'd5; a_sign2 = 4'd2; a_sign3 = 4'd0;
b_sign0 = 4'd12; b_sign1 = 4'd7; b_sign2 = 4'd15; b_sign3 = 4'd10;
@(posedge clk_i);
a_mant0 = 8'd233; a_mant1 = 8'd80; a_mant2 = 8'd208; a_mant3 = 8'd161;
b_mant0 = 8'd87; b_mant1 = 8'd160; b_mant2 = 8'd127; b_mant3 = 8'd84;
a_exp0 = 10'd364; a_exp1 = 10'd905; a_exp2 = 10'd1008; a_exp3 = 10'd586;
b_exp0 = 10'd187; b_exp1 = 10'd770; b_exp2 = 10'd1005; b_exp3 = 10'd448;
a_sign0 = 4'd14; a_sign1 = 4'd8; a_sign2 = 4'd2; a_sign3 = 4'd4;
b_sign0 = 4'd9; b_sign1 = 4'd13; b_sign2 = 4'd8; b_sign3 = 4'd15;
@(posedge clk_i);
shared_exps0 = 8'd131;
shared_exps1 = 8'd114;
a_mant0 = 8'd47; a_mant1 = 8'd222; a_mant2 = 8'd63; a_mant3 = 8'd30;
b_mant0 = 8'd85; b_mant1 = 8'd118; b_mant2 = 8'd229; b_mant3 = 8'd212;
a_exp0 = 10'd502; a_exp1 = 10'd127; a_exp2 = 10'd988; a_exp3 = 10'd141;
b_exp0 = 10'd237; b_exp1 = 10'd877; b_exp2 = 10'd3; b_exp3 = 10'd458;
a_sign0 = 4'd16; a_sign1 = 4'd13; a_sign2 = 4'd6; a_sign3 = 4'd14;
b_sign0 = 4'd3; b_sign1 = 4'd5; b_sign2 = 4'd12; b_sign3 = 4'd1;
@(posedge clk_i);
a_mant0 = 8'd73; a_mant1 = 8'd104; a_mant2 = 8'd84; a_mant3 = 8'd82;
b_mant0 = 8'd118; b_mant1 = 8'd176; b_mant2 = 8'd154; b_mant3 = 8'd217;
a_exp0 = 10'd692; a_exp1 = 10'd751; a_exp2 = 10'd307; a_exp3 = 10'd506;
b_exp0 = 10'd706; b_exp1 = 10'd872; b_exp2 = 10'd521; b_exp3 = 10'd586;
a_sign0 = 4'd13; a_sign1 = 4'd14; a_sign2 = 4'd14; a_sign3 = 4'd10;
b_sign0 = 4'd13; b_sign1 = 4'd12; b_sign2 = 4'd12; b_sign3 = 4'd15;
@(posedge clk_i);
a_mant0 = 8'd42; a_mant1 = 8'd160; a_mant2 = 8'd120; a_mant3 = 8'd76;
b_mant0 = 8'd158; b_mant1 = 8'd204; b_mant2 = 8'd235; b_mant3 = 8'd205;
a_exp0 = 10'd725; a_exp1 = 10'd132; a_exp2 = 10'd797; a_exp3 = 10'd122;
b_exp0 = 10'd310; b_exp1 = 10'd324; b_exp2 = 10'd709; b_exp3 = 10'd437;
a_sign0 = 4'd8; a_sign1 = 4'd4; a_sign2 = 4'd12; a_sign3 = 4'd10;
b_sign0 = 4'd6; b_sign1 = 4'd12; b_sign2 = 4'd13; b_sign3 = 4'd4;
@(posedge clk_i);
a_mant0 = 8'd175; a_mant1 = 8'd59; a_mant2 = 8'd200; a_mant3 = 8'd239;
b_mant0 = 8'd185; b_mant1 = 8'd176; b_mant2 = 8'd229; b_mant3 = 8'd192;
a_exp0 = 10'd978; a_exp1 = 10'd251; a_exp2 = 10'd952; a_exp3 = 10'd494;
b_exp0 = 10'd430; b_exp1 = 10'd598; b_exp2 = 10'd941; b_exp3 = 10'd68;
a_sign0 = 4'd11; a_sign1 = 4'd5; a_sign2 = 4'd8; a_sign3 = 4'd9;
b_sign0 = 4'd6; b_sign1 = 4'd12; b_sign2 = 4'd16; b_sign3 = 4'd10;
@(posedge clk_i);
a_mant0 = 8'd152; a_mant1 = 8'd35; a_mant2 = 8'd170; a_mant3 = 8'd185;
b_mant0 = 8'd90; b_mant1 = 8'd170; b_mant2 = 8'd73; b_mant3 = 8'd142;
a_exp0 = 10'd841; a_exp1 = 10'd31; a_exp2 = 10'd556; a_exp3 = 10'd171;
b_exp0 = 10'd943; b_exp1 = 10'd14; b_exp2 = 10'd892; b_exp3 = 10'd1000;
a_sign0 = 4'd1; a_sign1 = 4'd12; a_sign2 = 4'd13; a_sign3 = 4'd7;
b_sign0 = 4'd6; b_sign1 = 4'd13; b_sign2 = 4'd5; b_sign3 = 4'd2;
@(posedge clk_i);
a_mant0 = 8'd190; a_mant1 = 8'd216; a_mant2 = 8'd109; a_mant3 = 8'd105;
b_mant0 = 8'd207; b_mant1 = 8'd5; b_mant2 = 8'd95; b_mant3 = 8'd235;
a_exp0 = 10'd434; a_exp1 = 10'd11; a_exp2 = 10'd296; a_exp3 = 10'd124;
b_exp0 = 10'd204; b_exp1 = 10'd673; b_exp2 = 10'd753; b_exp3 = 10'd787;
a_sign0 = 4'd14; a_sign1 = 4'd12; a_sign2 = 4'd9; a_sign3 = 4'd10;
b_sign0 = 4'd9; b_sign1 = 4'd11; b_sign2 = 4'd13; b_sign3 = 4'd7;
@(posedge clk_i);
a_mant0 = 8'd60; a_mant1 = 8'd113; a_mant2 = 8'd215; a_mant3 = 8'd136;
b_mant0 = 8'd102; b_mant1 = 8'd38; b_mant2 = 8'd128; b_mant3 = 8'd51;
a_exp0 = 10'd611; a_exp1 = 10'd454; a_exp2 = 10'd343; a_exp3 = 10'd542;
b_exp0 = 10'd806; b_exp1 = 10'd120; b_exp2 = 10'd702; b_exp3 = 10'd2;
a_sign0 = 4'd2; a_sign1 = 4'd9; a_sign2 = 4'd16; a_sign3 = 4'd0;
b_sign0 = 4'd8; b_sign1 = 4'd15; b_sign2 = 4'd6; b_sign3 = 4'd12;
@(posedge clk_i);
a_mant0 = 8'd128; a_mant1 = 8'd17; a_mant2 = 8'd226; a_mant3 = 8'd117;
b_mant0 = 8'd121; b_mant1 = 8'd174; b_mant2 = 8'd123; b_mant3 = 8'd226;
a_exp0 = 10'd991; a_exp1 = 10'd161; a_exp2 = 10'd728; a_exp3 = 10'd939;
b_exp0 = 10'd963; b_exp1 = 10'd628; b_exp2 = 10'd525; b_exp3 = 10'd580;
a_sign0 = 4'd12; a_sign1 = 4'd10; a_sign2 = 4'd7; a_sign3 = 4'd1;
b_sign0 = 4'd12; b_sign1 = 4'd8; b_sign2 = 4'd10; b_sign3 = 4'd14;
@(posedge clk_i);
shared_exps0 = 8'd83;
shared_exps1 = 8'd130;
a_mant0 = 8'd72; a_mant1 = 8'd205; a_mant2 = 8'd107; a_mant3 = 8'd223;
b_mant0 = 8'd33; b_mant1 = 8'd31; b_mant2 = 8'd8; b_mant3 = 8'd124;
a_exp0 = 10'd959; a_exp1 = 10'd800; a_exp2 = 10'd933; a_exp3 = 10'd600;
b_exp0 = 10'd606; b_exp1 = 10'd221; b_exp2 = 10'd353; b_exp3 = 10'd1016;
a_sign0 = 4'd8; a_sign1 = 4'd3; a_sign2 = 4'd0; a_sign3 = 4'd16;
b_sign0 = 4'd12; b_sign1 = 4'd9; b_sign2 = 4'd11; b_sign3 = 4'd12;
@(posedge clk_i);
a_mant0 = 8'd237; a_mant1 = 8'd148; a_mant2 = 8'd98; a_mant3 = 8'd121;
b_mant0 = 8'd124; b_mant1 = 8'd130; b_mant2 = 8'd253; b_mant3 = 8'd202;
a_exp0 = 10'd515; a_exp1 = 10'd578; a_exp2 = 10'd246; a_exp3 = 10'd159;
b_exp0 = 10'd699; b_exp1 = 10'd493; b_exp2 = 10'd734; b_exp3 = 10'd242;
a_sign0 = 4'd11; a_sign1 = 4'd8; a_sign2 = 4'd4; a_sign3 = 4'd0;
b_sign0 = 4'd0; b_sign1 = 4'd5; b_sign2 = 4'd1; b_sign3 = 4'd2;
@(posedge clk_i);
a_mant0 = 8'd105; a_mant1 = 8'd196; a_mant2 = 8'd100; a_mant3 = 8'd156;
b_mant0 = 8'd210; b_mant1 = 8'd97; b_mant2 = 8'd96; b_mant3 = 8'd80;
a_exp0 = 10'd296; a_exp1 = 10'd779; a_exp2 = 10'd572; a_exp3 = 10'd227;
b_exp0 = 10'd149; b_exp1 = 10'd877; b_exp2 = 10'd125; b_exp3 = 10'd285;
a_sign0 = 4'd15; a_sign1 = 4'd14; a_sign2 = 4'd4; a_sign3 = 4'd6;
b_sign0 = 4'd1; b_sign1 = 4'd1; b_sign2 = 4'd8; b_sign3 = 4'd7;
@(posedge clk_i);
a_mant0 = 8'd21; a_mant1 = 8'd79; a_mant2 = 8'd198; a_mant3 = 8'd80;
b_mant0 = 8'd53; b_mant1 = 8'd238; b_mant2 = 8'd233; b_mant3 = 8'd247;
a_exp0 = 10'd416; a_exp1 = 10'd38; a_exp2 = 10'd787; a_exp3 = 10'd691;
b_exp0 = 10'd992; b_exp1 = 10'd575; b_exp2 = 10'd142; b_exp3 = 10'd443;
a_sign0 = 4'd15; a_sign1 = 4'd13; a_sign2 = 4'd14; a_sign3 = 4'd9;
b_sign0 = 4'd0; b_sign1 = 4'd15; b_sign2 = 4'd11; b_sign3 = 4'd1;
@(posedge clk_i);
a_mant0 = 8'd57; a_mant1 = 8'd184; a_mant2 = 8'd47; a_mant3 = 8'd232;
b_mant0 = 8'd243; b_mant1 = 8'd153; b_mant2 = 8'd220; b_mant3 = 8'd35;
a_exp0 = 10'd877; a_exp1 = 10'd519; a_exp2 = 10'd712; a_exp3 = 10'd787;
b_exp0 = 10'd263; b_exp1 = 10'd653; b_exp2 = 10'd366; b_exp3 = 10'd118;
a_sign0 = 4'd13; a_sign1 = 4'd10; a_sign2 = 4'd11; a_sign3 = 4'd10;
b_sign0 = 4'd11; b_sign1 = 4'd14; b_sign2 = 4'd11; b_sign3 = 4'd9;
@(posedge clk_i);
a_mant0 = 8'd80; a_mant1 = 8'd146; a_mant2 = 8'd47; a_mant3 = 8'd187;
b_mant0 = 8'd67; b_mant1 = 8'd215; b_mant2 = 8'd66; b_mant3 = 8'd13;
a_exp0 = 10'd113; a_exp1 = 10'd940; a_exp2 = 10'd277; a_exp3 = 10'd26;
b_exp0 = 10'd950; b_exp1 = 10'd851; b_exp2 = 10'd170; b_exp3 = 10'd151;
a_sign0 = 4'd5; a_sign1 = 4'd14; a_sign2 = 4'd15; a_sign3 = 4'd5;
b_sign0 = 4'd14; b_sign1 = 4'd4; b_sign2 = 4'd11; b_sign3 = 4'd8;
@(posedge clk_i);
a_mant0 = 8'd222; a_mant1 = 8'd26; a_mant2 = 8'd149; a_mant3 = 8'd55;
b_mant0 = 8'd13; b_mant1 = 8'd168; b_mant2 = 8'd120; b_mant3 = 8'd233;
a_exp0 = 10'd120; a_exp1 = 10'd132; a_exp2 = 10'd725; a_exp3 = 10'd498;
b_exp0 = 10'd251; b_exp1 = 10'd466; b_exp2 = 10'd1022; b_exp3 = 10'd150;
a_sign0 = 4'd14; a_sign1 = 4'd7; a_sign2 = 4'd15; a_sign3 = 4'd9;
b_sign0 = 4'd0; b_sign1 = 4'd8; b_sign2 = 4'd13; b_sign3 = 4'd0;
@(posedge clk_i);
a_mant0 = 8'd125; a_mant1 = 8'd79; a_mant2 = 8'd51; a_mant3 = 8'd26;
b_mant0 = 8'd216; b_mant1 = 8'd56; b_mant2 = 8'd171; b_mant3 = 8'd103;
a_exp0 = 10'd447; a_exp1 = 10'd907; a_exp2 = 10'd316; a_exp3 = 10'd727;
b_exp0 = 10'd410; b_exp1 = 10'd31; b_exp2 = 10'd540; b_exp3 = 10'd3;
a_sign0 = 4'd1; a_sign1 = 4'd6; a_sign2 = 4'd2; a_sign3 = 4'd6;
b_sign0 = 4'd4; b_sign1 = 4'd16; b_sign2 = 4'd2; b_sign3 = 4'd7;
@(posedge clk_i);
shared_exps0 = 8'd139;
shared_exps1 = 8'd119;
rstn = 0;
@(posedge clk_i);
rstn = 1;
a_mant0 = 8'd162; a_mant1 = 8'd26; a_mant2 = 8'd44; a_mant3 = 8'd251;
b_mant0 = 8'd84; b_mant1 = 8'd87; b_mant2 = 8'd0; b_mant3 = 8'd209;
a_exp0 = 10'd797; a_exp1 = 10'd137; a_exp2 = 10'd619; a_exp3 = 10'd621;
b_exp0 = 10'd151; b_exp1 = 10'd676; b_exp2 = 10'd375; b_exp3 = 10'd9;
a_sign0 = 4'd3; a_sign1 = 4'd3; a_sign2 = 4'd11; a_sign3 = 4'd13;
b_sign0 = 4'd0; b_sign1 = 4'd14; b_sign2 = 4'd2; b_sign3 = 4'd14;
@(posedge clk_i);
a_mant0 = 8'd150; a_mant1 = 8'd76; a_mant2 = 8'd77; a_mant3 = 8'd116;
b_mant0 = 8'd226; b_mant1 = 8'd252; b_mant2 = 8'd136; b_mant3 = 8'd116;
a_exp0 = 10'd715; a_exp1 = 10'd860; a_exp2 = 10'd368; a_exp3 = 10'd104;
b_exp0 = 10'd127; b_exp1 = 10'd63; b_exp2 = 10'd575; b_exp3 = 10'd158;
a_sign0 = 4'd5; a_sign1 = 4'd7; a_sign2 = 4'd16; a_sign3 = 4'd9;
b_sign0 = 4'd3; b_sign1 = 4'd8; b_sign2 = 4'd8; b_sign3 = 4'd13;
@(posedge clk_i);
a_mant0 = 8'd153; a_mant1 = 8'd29; a_mant2 = 8'd240; a_mant3 = 8'd170;
b_mant0 = 8'd212; b_mant1 = 8'd197; b_mant2 = 8'd49; b_mant3 = 8'd194;
a_exp0 = 10'd795; a_exp1 = 10'd331; a_exp2 = 10'd358; a_exp3 = 10'd907;
b_exp0 = 10'd142; b_exp1 = 10'd189; b_exp2 = 10'd683; b_exp3 = 10'd124;
a_sign0 = 4'd15; a_sign1 = 4'd13; a_sign2 = 4'd1; a_sign3 = 4'd2;
b_sign0 = 4'd12; b_sign1 = 4'd8; b_sign2 = 4'd11; b_sign3 = 4'd0;
@(posedge clk_i);
a_mant0 = 8'd150; a_mant1 = 8'd18; a_mant2 = 8'd64; a_mant3 = 8'd121;
b_mant0 = 8'd91; b_mant1 = 8'd75; b_mant2 = 8'd255; b_mant3 = 8'd113;
a_exp0 = 10'd49; a_exp1 = 10'd526; a_exp2 = 10'd68; a_exp3 = 10'd500;
b_exp0 = 10'd698; b_exp1 = 10'd443; b_exp2 = 10'd553; b_exp3 = 10'd431;
a_sign0 = 4'd5; a_sign1 = 4'd4; a_sign2 = 4'd9; a_sign3 = 4'd3;
b_sign0 = 4'd6; b_sign1 = 4'd5; b_sign2 = 4'd7; b_sign3 = 4'd5;
@(posedge clk_i);
a_mant0 = 8'd30; a_mant1 = 8'd227; a_mant2 = 8'd24; a_mant3 = 8'd188;
b_mant0 = 8'd236; b_mant1 = 8'd215; b_mant2 = 8'd41; b_mant3 = 8'd194;
a_exp0 = 10'd683; a_exp1 = 10'd245; a_exp2 = 10'd628; a_exp3 = 10'd106;
b_exp0 = 10'd899; b_exp1 = 10'd397; b_exp2 = 10'd578; b_exp3 = 10'd698;
a_sign0 = 4'd12; a_sign1 = 4'd4; a_sign2 = 4'd2; a_sign3 = 4'd9;
b_sign0 = 4'd14; b_sign1 = 4'd16; b_sign2 = 4'd11; b_sign3 = 4'd15;
@(posedge clk_i);
a_mant0 = 8'd125; a_mant1 = 8'd66; a_mant2 = 8'd199; a_mant3 = 8'd31;
b_mant0 = 8'd215; b_mant1 = 8'd183; b_mant2 = 8'd79; b_mant3 = 8'd5;
a_exp0 = 10'd435; a_exp1 = 10'd754; a_exp2 = 10'd263; a_exp3 = 10'd279;
b_exp0 = 10'd677; b_exp1 = 10'd979; b_exp2 = 10'd59; b_exp3 = 10'd328;
a_sign0 = 4'd5; a_sign1 = 4'd1; a_sign2 = 4'd14; a_sign3 = 4'd7;
b_sign0 = 4'd16; b_sign1 = 4'd11; b_sign2 = 4'd16; b_sign3 = 4'd12;
@(posedge clk_i);
a_mant0 = 8'd219; a_mant1 = 8'd106; a_mant2 = 8'd83; a_mant3 = 8'd149;
b_mant0 = 8'd177; b_mant1 = 8'd219; b_mant2 = 8'd52; b_mant3 = 8'd224;
a_exp0 = 10'd357; a_exp1 = 10'd745; a_exp2 = 10'd1000; a_exp3 = 10'd274;
b_exp0 = 10'd32; b_exp1 = 10'd483; b_exp2 = 10'd658; b_exp3 = 10'd345;
a_sign0 = 4'd2; a_sign1 = 4'd15; a_sign2 = 4'd6; a_sign3 = 4'd7;
b_sign0 = 4'd16; b_sign1 = 4'd12; b_sign2 = 4'd1; b_sign3 = 4'd3;
@(posedge clk_i);
shared_exps0 = 8'd127;
shared_exps1 = 8'd123;
a_mant0 = 8'd229; a_mant1 = 8'd204; a_mant2 = 8'd174; a_mant3 = 8'd64;
b_mant0 = 8'd123; b_mant1 = 8'd45; b_mant2 = 8'd48; b_mant3 = 8'd171;
a_exp0 = 10'd128; a_exp1 = 10'd542; a_exp2 = 10'd516; a_exp3 = 10'd403;
b_exp0 = 10'd887; b_exp1 = 10'd385; b_exp2 = 10'd15; b_exp3 = 10'd840;
a_sign0 = 4'd6; a_sign1 = 4'd14; a_sign2 = 4'd9; a_sign3 = 4'd12;
b_sign0 = 4'd9; b_sign1 = 4'd13; b_sign2 = 4'd0; b_sign3 = 4'd12;
@(posedge clk_i);
a_mant0 = 8'd34; a_mant1 = 8'd69; a_mant2 = 8'd222; a_mant3 = 8'd53;
b_mant0 = 8'd108; b_mant1 = 8'd242; b_mant2 = 8'd29; b_mant3 = 8'd215;
a_exp0 = 10'd502; a_exp1 = 10'd240; a_exp2 = 10'd905; a_exp3 = 10'd230;
b_exp0 = 10'd49; b_exp1 = 10'd259; b_exp2 = 10'd383; b_exp3 = 10'd623;
a_sign0 = 4'd2; a_sign1 = 4'd7; a_sign2 = 4'd8; a_sign3 = 4'd11;
b_sign0 = 4'd4; b_sign1 = 4'd7; b_sign2 = 4'd1; b_sign3 = 4'd9;
@(posedge clk_i);
a_mant0 = 8'd221; a_mant1 = 8'd233; a_mant2 = 8'd82; a_mant3 = 8'd92;
b_mant0 = 8'd30; b_mant1 = 8'd51; b_mant2 = 8'd103; b_mant3 = 8'd61;
a_exp0 = 10'd846; a_exp1 = 10'd1010; a_exp2 = 10'd185; a_exp3 = 10'd502;
b_exp0 = 10'd346; b_exp1 = 10'd780; b_exp2 = 10'd402; b_exp3 = 10'd225;
a_sign0 = 4'd0; a_sign1 = 4'd5; a_sign2 = 4'd5; a_sign3 = 4'd8;
b_sign0 = 4'd9; b_sign1 = 4'd11; b_sign2 = 4'd2; b_sign3 = 4'd16;
@(posedge clk_i);
a_mant0 = 8'd100; a_mant1 = 8'd210; a_mant2 = 8'd146; a_mant3 = 8'd183;
b_mant0 = 8'd81; b_mant1 = 8'd23; b_mant2 = 8'd166; b_mant3 = 8'd35;
a_exp0 = 10'd881; a_exp1 = 10'd625; a_exp2 = 10'd736; a_exp3 = 10'd820;
b_exp0 = 10'd739; b_exp1 = 10'd238; b_exp2 = 10'd720; b_exp3 = 10'd119;
a_sign0 = 4'd7; a_sign1 = 4'd5; a_sign2 = 4'd9; a_sign3 = 4'd15;
b_sign0 = 4'd4; b_sign1 = 4'd9; b_sign2 = 4'd5; b_sign3 = 4'd9;
@(posedge clk_i);
a_mant0 = 8'd61; a_mant1 = 8'd230; a_mant2 = 8'd143; a_mant3 = 8'd237;
b_mant0 = 8'd73; b_mant1 = 8'd3; b_mant2 = 8'd45; b_mant3 = 8'd35;
a_exp0 = 10'd542; a_exp1 = 10'd422; a_exp2 = 10'd213; a_exp3 = 10'd779;
b_exp0 = 10'd949; b_exp1 = 10'd457; b_exp2 = 10'd263; b_exp3 = 10'd902;
a_sign0 = 4'd3; a_sign1 = 4'd1; a_sign2 = 4'd1; a_sign3 = 4'd7;
b_sign0 = 4'd13; b_sign1 = 4'd2; b_sign2 = 4'd1; b_sign3 = 4'd5;
@(posedge clk_i);
a_mant0 = 8'd11; a_mant1 = 8'd181; a_mant2 = 8'd140; a_mant3 = 8'd109;
b_mant0 = 8'd240; b_mant1 = 8'd213; b_mant2 = 8'd72; b_mant3 = 8'd225;
a_exp0 = 10'd155; a_exp1 = 10'd685; a_exp2 = 10'd58; a_exp3 = 10'd82;
b_exp0 = 10'd103; b_exp1 = 10'd376; b_exp2 = 10'd171; b_exp3 = 10'd675;
a_sign0 = 4'd14; a_sign1 = 4'd1; a_sign2 = 4'd3; a_sign3 = 4'd10;
b_sign0 = 4'd11; b_sign1 = 4'd12; b_sign2 = 4'd5; b_sign3 = 4'd14;
@(posedge clk_i);
a_mant0 = 8'd177; a_mant1 = 8'd89; a_mant2 = 8'd33; a_mant3 = 8'd194;
b_mant0 = 8'd113; b_mant1 = 8'd28; b_mant2 = 8'd37; b_mant3 = 8'd41;
a_exp0 = 10'd686; a_exp1 = 10'd720; a_exp2 = 10'd48; a_exp3 = 10'd610;
b_exp0 = 10'd450; b_exp1 = 10'd141; b_exp2 = 10'd939; b_exp3 = 10'd833;
a_sign0 = 4'd8; a_sign1 = 4'd16; a_sign2 = 4'd14; a_sign3 = 4'd6;
b_sign0 = 4'd14; b_sign1 = 4'd16; b_sign2 = 4'd0; b_sign3 = 4'd8;
@(posedge clk_i);
a_mant0 = 8'd97; a_mant1 = 8'd219; a_mant2 = 8'd168; a_mant3 = 8'd127;
b_mant0 = 8'd44; b_mant1 = 8'd64; b_mant2 = 8'd63; b_mant3 = 8'd198;
a_exp0 = 10'd234; a_exp1 = 10'd342; a_exp2 = 10'd957; a_exp3 = 10'd884;
b_exp0 = 10'd817; b_exp1 = 10'd614; b_exp2 = 10'd486; b_exp3 = 10'd368;
a_sign0 = 4'd12; a_sign1 = 4'd10; a_sign2 = 4'd8; a_sign3 = 4'd7;
b_sign0 = 4'd10; b_sign1 = 4'd9; b_sign2 = 4'd8; b_sign3 = 4'd15;
@(posedge clk_i);
shared_exps0 = 8'd132;
shared_exps1 = 8'd144;
a_mant0 = 8'd132; a_mant1 = 8'd226; a_mant2 = 8'd27; a_mant3 = 8'd206;
b_mant0 = 8'd178; b_mant1 = 8'd50; b_mant2 = 8'd167; b_mant3 = 8'd52;
a_exp0 = 10'd272; a_exp1 = 10'd1012; a_exp2 = 10'd605; a_exp3 = 10'd697;
b_exp0 = 10'd784; b_exp1 = 10'd388; b_exp2 = 10'd381; b_exp3 = 10'd648;
a_sign0 = 4'd16; a_sign1 = 4'd10; a_sign2 = 4'd5; a_sign3 = 4'd3;
b_sign0 = 4'd5; b_sign1 = 4'd14; b_sign2 = 4'd11; b_sign3 = 4'd15;
@(posedge clk_i);
a_mant0 = 8'd151; a_mant1 = 8'd107; a_mant2 = 8'd23; a_mant3 = 8'd88;
b_mant0 = 8'd4; b_mant1 = 8'd147; b_mant2 = 8'd132; b_mant3 = 8'd188;
a_exp0 = 10'd982; a_exp1 = 10'd22; a_exp2 = 10'd643; a_exp3 = 10'd102;
b_exp0 = 10'd113; b_exp1 = 10'd692; b_exp2 = 10'd948; b_exp3 = 10'd694;
a_sign0 = 4'd3; a_sign1 = 4'd10; a_sign2 = 4'd5; a_sign3 = 4'd4;
b_sign0 = 4'd3; b_sign1 = 4'd0; b_sign2 = 4'd9; b_sign3 = 4'd1;
@(posedge clk_i);
a_mant0 = 8'd205; a_mant1 = 8'd162; a_mant2 = 8'd114; a_mant3 = 8'd87;
b_mant0 = 8'd55; b_mant1 = 8'd35; b_mant2 = 8'd165; b_mant3 = 8'd255;
a_exp0 = 10'd232; a_exp1 = 10'd391; a_exp2 = 10'd328; a_exp3 = 10'd892;
b_exp0 = 10'd678; b_exp1 = 10'd811; b_exp2 = 10'd574; b_exp3 = 10'd907;
a_sign0 = 4'd5; a_sign1 = 4'd14; a_sign2 = 4'd16; a_sign3 = 4'd15;
b_sign0 = 4'd14; b_sign1 = 4'd8; b_sign2 = 4'd4; b_sign3 = 4'd12;
@(posedge clk_i);
a_mant0 = 8'd141; a_mant1 = 8'd233; a_mant2 = 8'd210; a_mant3 = 8'd85;
b_mant0 = 8'd42; b_mant1 = 8'd132; b_mant2 = 8'd38; b_mant3 = 8'd143;
a_exp0 = 10'd20; a_exp1 = 10'd502; a_exp2 = 10'd758; a_exp3 = 10'd865;
b_exp0 = 10'd449; b_exp1 = 10'd707; b_exp2 = 10'd310; b_exp3 = 10'd257;
a_sign0 = 4'd2; a_sign1 = 4'd0; a_sign2 = 4'd4; a_sign3 = 4'd15;
b_sign0 = 4'd1; b_sign1 = 4'd9; b_sign2 = 4'd8; b_sign3 = 4'd15;
@(posedge clk_i);
a_mant0 = 8'd192; a_mant1 = 8'd15; a_mant2 = 8'd186; a_mant3 = 8'd239;
b_mant0 = 8'd19; b_mant1 = 8'd123; b_mant2 = 8'd103; b_mant3 = 8'd31;
a_exp0 = 10'd911; a_exp1 = 10'd712; a_exp2 = 10'd549; a_exp3 = 10'd188;
b_exp0 = 10'd949; b_exp1 = 10'd697; b_exp2 = 10'd448; b_exp3 = 10'd173;
a_sign0 = 4'd9; a_sign1 = 4'd14; a_sign2 = 4'd3; a_sign3 = 4'd11;
b_sign0 = 4'd0; b_sign1 = 4'd11; b_sign2 = 4'd9; b_sign3 = 4'd0;
@(posedge clk_i);
a_mant0 = 8'd120; a_mant1 = 8'd4; a_mant2 = 8'd138; a_mant3 = 8'd168;
b_mant0 = 8'd189; b_mant1 = 8'd140; b_mant2 = 8'd4; b_mant3 = 8'd191;
a_exp0 = 10'd877; a_exp1 = 10'd200; a_exp2 = 10'd735; a_exp3 = 10'd770;
b_exp0 = 10'd65; b_exp1 = 10'd543; b_exp2 = 10'd21; b_exp3 = 10'd541;
a_sign0 = 4'd5; a_sign1 = 4'd7; a_sign2 = 4'd3; a_sign3 = 4'd1;
b_sign0 = 4'd6; b_sign1 = 4'd2; b_sign2 = 4'd3; b_sign3 = 4'd0;
@(posedge clk_i);
a_mant0 = 8'd71; a_mant1 = 8'd251; a_mant2 = 8'd124; a_mant3 = 8'd224;
b_mant0 = 8'd168; b_mant1 = 8'd40; b_mant2 = 8'd135; b_mant3 = 8'd110;
a_exp0 = 10'd408; a_exp1 = 10'd484; a_exp2 = 10'd314; a_exp3 = 10'd176;
b_exp0 = 10'd918; b_exp1 = 10'd426; b_exp2 = 10'd361; b_exp3 = 10'd686;
a_sign0 = 4'd0; a_sign1 = 4'd2; a_sign2 = 4'd6; a_sign3 = 4'd13;
b_sign0 = 4'd7; b_sign1 = 4'd16; b_sign2 = 4'd14; b_sign3 = 4'd16;
@(posedge clk_i);
a_mant0 = 8'd254; a_mant1 = 8'd170; a_mant2 = 8'd44; a_mant3 = 8'd47;
b_mant0 = 8'd75; b_mant1 = 8'd156; b_mant2 = 8'd71; b_mant3 = 8'd229;
a_exp0 = 10'd378; a_exp1 = 10'd472; a_exp2 = 10'd501; a_exp3 = 10'd854;
b_exp0 = 10'd706; b_exp1 = 10'd102; b_exp2 = 10'd177; b_exp3 = 10'd924;
a_sign0 = 4'd12; a_sign1 = 4'd1; a_sign2 = 4'd8; a_sign3 = 4'd1;
b_sign0 = 4'd9; b_sign1 = 4'd0; b_sign2 = 4'd5; b_sign3 = 4'd8;
@(posedge clk_i);
shared_exps0 = 8'd136;
shared_exps1 = 8'd136;
a_mant0 = 8'd189; a_mant1 = 8'd206; a_mant2 = 8'd66; a_mant3 = 8'd188;
b_mant0 = 8'd58; b_mant1 = 8'd47; b_mant2 = 8'd169; b_mant3 = 8'd105;
a_exp0 = 10'd841; a_exp1 = 10'd618; a_exp2 = 10'd593; a_exp3 = 10'd520;
b_exp0 = 10'd795; b_exp1 = 10'd314; b_exp2 = 10'd868; b_exp3 = 10'd728;
a_sign0 = 4'd5; a_sign1 = 4'd11; a_sign2 = 4'd11; a_sign3 = 4'd16;
b_sign0 = 4'd4; b_sign1 = 4'd4; b_sign2 = 4'd10; b_sign3 = 4'd7;
@(posedge clk_i);
a_mant0 = 8'd5; a_mant1 = 8'd196; a_mant2 = 8'd52; a_mant3 = 8'd149;
b_mant0 = 8'd74; b_mant1 = 8'd175; b_mant2 = 8'd227; b_mant3 = 8'd186;
a_exp0 = 10'd273; a_exp1 = 10'd306; a_exp2 = 10'd566; a_exp3 = 10'd12;
b_exp0 = 10'd967; b_exp1 = 10'd943; b_exp2 = 10'd419; b_exp3 = 10'd880;
a_sign0 = 4'd14; a_sign1 = 4'd14; a_sign2 = 4'd13; a_sign3 = 4'd10;
b_sign0 = 4'd2; b_sign1 = 4'd5; b_sign2 = 4'd4; b_sign3 = 4'd10;
@(posedge clk_i);
a_mant0 = 8'd87; a_mant1 = 8'd180; a_mant2 = 8'd57; a_mant3 = 8'd179;
b_mant0 = 8'd153; b_mant1 = 8'd135; b_mant2 = 8'd230; b_mant3 = 8'd216;
a_exp0 = 10'd4; a_exp1 = 10'd363; a_exp2 = 10'd809; a_exp3 = 10'd516;
b_exp0 = 10'd570; b_exp1 = 10'd659; b_exp2 = 10'd944; b_exp3 = 10'd342;
a_sign0 = 4'd11; a_sign1 = 4'd0; a_sign2 = 4'd7; a_sign3 = 4'd4;
b_sign0 = 4'd11; b_sign1 = 4'd1; b_sign2 = 4'd2; b_sign3 = 4'd8;
@(posedge clk_i);
a_mant0 = 8'd156; a_mant1 = 8'd112; a_mant2 = 8'd31; a_mant3 = 8'd234;
b_mant0 = 8'd108; b_mant1 = 8'd35; b_mant2 = 8'd146; b_mant3 = 8'd96;
a_exp0 = 10'd426; a_exp1 = 10'd272; a_exp2 = 10'd378; a_exp3 = 10'd115;
b_exp0 = 10'd78; b_exp1 = 10'd554; b_exp2 = 10'd772; b_exp3 = 10'd690;
a_sign0 = 4'd9; a_sign1 = 4'd12; a_sign2 = 4'd4; a_sign3 = 4'd10;
b_sign0 = 4'd10; b_sign1 = 4'd16; b_sign2 = 4'd2; b_sign3 = 4'd13;
@(posedge clk_i);
a_mant0 = 8'd227; a_mant1 = 8'd230; a_mant2 = 8'd140; a_mant3 = 8'd50;
b_mant0 = 8'd52; b_mant1 = 8'd59; b_mant2 = 8'd139; b_mant3 = 8'd209;
a_exp0 = 10'd224; a_exp1 = 10'd809; a_exp2 = 10'd585; a_exp3 = 10'd194;
b_exp0 = 10'd216; b_exp1 = 10'd688; b_exp2 = 10'd383; b_exp3 = 10'd428;
a_sign0 = 4'd12; a_sign1 = 4'd15; a_sign2 = 4'd9; a_sign3 = 4'd9;
b_sign0 = 4'd10; b_sign1 = 4'd10; b_sign2 = 4'd1; b_sign3 = 4'd13;
@(posedge clk_i);
a_mant0 = 8'd59; a_mant1 = 8'd148; a_mant2 = 8'd62; a_mant3 = 8'd227;
b_mant0 = 8'd140; b_mant1 = 8'd233; b_mant2 = 8'd233; b_mant3 = 8'd222;
a_exp0 = 10'd635; a_exp1 = 10'd328; a_exp2 = 10'd495; a_exp3 = 10'd325;
b_exp0 = 10'd132; b_exp1 = 10'd997; b_exp2 = 10'd496; b_exp3 = 10'd732;
a_sign0 = 4'd0; a_sign1 = 4'd5; a_sign2 = 4'd0; a_sign3 = 4'd14;
b_sign0 = 4'd1; b_sign1 = 4'd8; b_sign2 = 4'd11; b_sign3 = 4'd3;
@(posedge clk_i);
a_mant0 = 8'd2; a_mant1 = 8'd35; a_mant2 = 8'd241; a_mant3 = 8'd1;
b_mant0 = 8'd0; b_mant1 = 8'd124; b_mant2 = 8'd74; b_mant3 = 8'd231;
a_exp0 = 10'd292; a_exp1 = 10'd393; a_exp2 = 10'd56; a_exp3 = 10'd260;
b_exp0 = 10'd605; b_exp1 = 10'd774; b_exp2 = 10'd143; b_exp3 = 10'd812;
a_sign0 = 4'd3; a_sign1 = 4'd9; a_sign2 = 4'd6; a_sign3 = 4'd10;
b_sign0 = 4'd6; b_sign1 = 4'd1; b_sign2 = 4'd13; b_sign3 = 4'd13;
@(posedge clk_i);
a_mant0 = 8'd239; a_mant1 = 8'd163; a_mant2 = 8'd193; a_mant3 = 8'd235;
b_mant0 = 8'd170; b_mant1 = 8'd167; b_mant2 = 8'd69; b_mant3 = 8'd227;
a_exp0 = 10'd544; a_exp1 = 10'd136; a_exp2 = 10'd575; a_exp3 = 10'd814;
b_exp0 = 10'd887; b_exp1 = 10'd21; b_exp2 = 10'd635; b_exp3 = 10'd508;
a_sign0 = 4'd8; a_sign1 = 4'd8; a_sign2 = 4'd5; a_sign3 = 4'd11;
b_sign0 = 4'd12; b_sign1 = 4'd12; b_sign2 = 4'd11; b_sign3 = 4'd7;
@(posedge clk_i);
shared_exps0 = 8'd125;
shared_exps1 = 8'd110;
rstn = 0;
@(posedge clk_i);
rstn = 1;
a_mant0 = 8'd109; a_mant1 = 8'd145; a_mant2 = 8'd75; a_mant3 = 8'd136;
b_mant0 = 8'd173; b_mant1 = 8'd137; b_mant2 = 8'd253; b_mant3 = 8'd27;
a_exp0 = 10'd523; a_exp1 = 10'd112; a_exp2 = 10'd525; a_exp3 = 10'd174;
b_exp0 = 10'd288; b_exp1 = 10'd96; b_exp2 = 10'd564; b_exp3 = 10'd55;
a_sign0 = 4'd14; a_sign1 = 4'd9; a_sign2 = 4'd13; a_sign3 = 4'd12;
b_sign0 = 4'd0; b_sign1 = 4'd5; b_sign2 = 4'd2; b_sign3 = 4'd5;
@(posedge clk_i);
a_mant0 = 8'd8; a_mant1 = 8'd149; a_mant2 = 8'd212; a_mant3 = 8'd8;
b_mant0 = 8'd240; b_mant1 = 8'd171; b_mant2 = 8'd216; b_mant3 = 8'd247;
a_exp0 = 10'd891; a_exp1 = 10'd141; a_exp2 = 10'd533; a_exp3 = 10'd522;
b_exp0 = 10'd987; b_exp1 = 10'd546; b_exp2 = 10'd771; b_exp3 = 10'd393;
a_sign0 = 4'd2; a_sign1 = 4'd10; a_sign2 = 4'd12; a_sign3 = 4'd16;
b_sign0 = 4'd8; b_sign1 = 4'd13; b_sign2 = 4'd7; b_sign3 = 4'd12;
@(posedge clk_i);
a_mant0 = 8'd226; a_mant1 = 8'd19; a_mant2 = 8'd157; a_mant3 = 8'd127;
b_mant0 = 8'd180; b_mant1 = 8'd70; b_mant2 = 8'd135; b_mant3 = 8'd51;
a_exp0 = 10'd27; a_exp1 = 10'd66; a_exp2 = 10'd101; a_exp3 = 10'd187;
b_exp0 = 10'd21; b_exp1 = 10'd941; b_exp2 = 10'd382; b_exp3 = 10'd887;
a_sign0 = 4'd7; a_sign1 = 4'd5; a_sign2 = 4'd14; a_sign3 = 4'd9;
b_sign0 = 4'd16; b_sign1 = 4'd0; b_sign2 = 4'd6; b_sign3 = 4'd9;
@(posedge clk_i);
a_mant0 = 8'd158; a_mant1 = 8'd185; a_mant2 = 8'd25; a_mant3 = 8'd60;
b_mant0 = 8'd232; b_mant1 = 8'd223; b_mant2 = 8'd23; b_mant3 = 8'd105;
a_exp0 = 10'd729; a_exp1 = 10'd874; a_exp2 = 10'd406; a_exp3 = 10'd173;
b_exp0 = 10'd759; b_exp1 = 10'd540; b_exp2 = 10'd896; b_exp3 = 10'd731;
a_sign0 = 4'd8; a_sign1 = 4'd9; a_sign2 = 4'd16; a_sign3 = 4'd7;
b_sign0 = 4'd13; b_sign1 = 4'd5; b_sign2 = 4'd13; b_sign3 = 4'd10;
@(posedge clk_i);
a_mant0 = 8'd222; a_mant1 = 8'd80; a_mant2 = 8'd171; a_mant3 = 8'd32;
b_mant0 = 8'd43; b_mant1 = 8'd85; b_mant2 = 8'd60; b_mant3 = 8'd1;
a_exp0 = 10'd73; a_exp1 = 10'd567; a_exp2 = 10'd615; a_exp3 = 10'd448;
b_exp0 = 10'd149; b_exp1 = 10'd593; b_exp2 = 10'd104; b_exp3 = 10'd429;
a_sign0 = 4'd10; a_sign1 = 4'd10; a_sign2 = 4'd2; a_sign3 = 4'd10;
b_sign0 = 4'd8; b_sign1 = 4'd1; b_sign2 = 4'd8; b_sign3 = 4'd13;
@(posedge clk_i);
a_mant0 = 8'd179; a_mant1 = 8'd111; a_mant2 = 8'd8; a_mant3 = 8'd76;
b_mant0 = 8'd212; b_mant1 = 8'd76; b_mant2 = 8'd107; b_mant3 = 8'd56;
a_exp0 = 10'd857; a_exp1 = 10'd376; a_exp2 = 10'd8; a_exp3 = 10'd290;
b_exp0 = 10'd873; b_exp1 = 10'd403; b_exp2 = 10'd596; b_exp3 = 10'd288;
a_sign0 = 4'd10; a_sign1 = 4'd9; a_sign2 = 4'd8; a_sign3 = 4'd16;
b_sign0 = 4'd7; b_sign1 = 4'd13; b_sign2 = 4'd7; b_sign3 = 4'd11;
@(posedge clk_i);
a_mant0 = 8'd103; a_mant1 = 8'd1; a_mant2 = 8'd118; a_mant3 = 8'd137;
b_mant0 = 8'd21; b_mant1 = 8'd75; b_mant2 = 8'd21; b_mant3 = 8'd254;
a_exp0 = 10'd782; a_exp1 = 10'd304; a_exp2 = 10'd884; a_exp3 = 10'd451;
b_exp0 = 10'd197; b_exp1 = 10'd581; b_exp2 = 10'd595; b_exp3 = 10'd383;
a_sign0 = 4'd9; a_sign1 = 4'd6; a_sign2 = 4'd0; a_sign3 = 4'd9;
b_sign0 = 4'd0; b_sign1 = 4'd7; b_sign2 = 4'd5; b_sign3 = 4'd9;
@(posedge clk_i);
shared_exps0 = 8'd118;
shared_exps1 = 8'd127;
a_mant0 = 8'd103; a_mant1 = 8'd214; a_mant2 = 8'd138; a_mant3 = 8'd95;
b_mant0 = 8'd153; b_mant1 = 8'd175; b_mant2 = 8'd205; b_mant3 = 8'd82;
a_exp0 = 10'd267; a_exp1 = 10'd965; a_exp2 = 10'd832; a_exp3 = 10'd264;
b_exp0 = 10'd586; b_exp1 = 10'd768; b_exp2 = 10'd587; b_exp3 = 10'd318;
a_sign0 = 4'd3; a_sign1 = 4'd2; a_sign2 = 4'd6; a_sign3 = 4'd2;
b_sign0 = 4'd0; b_sign1 = 4'd3; b_sign2 = 4'd3; b_sign3 = 4'd4;
@(posedge clk_i);
a_mant0 = 8'd212; a_mant1 = 8'd180; a_mant2 = 8'd196; a_mant3 = 8'd131;
b_mant0 = 8'd246; b_mant1 = 8'd162; b_mant2 = 8'd140; b_mant3 = 8'd21;
a_exp0 = 10'd297; a_exp1 = 10'd18; a_exp2 = 10'd404; a_exp3 = 10'd708;
b_exp0 = 10'd177; b_exp1 = 10'd401; b_exp2 = 10'd339; b_exp3 = 10'd955;
a_sign0 = 4'd15; a_sign1 = 4'd0; a_sign2 = 4'd1; a_sign3 = 4'd2;
b_sign0 = 4'd12; b_sign1 = 4'd4; b_sign2 = 4'd11; b_sign3 = 4'd13;
@(posedge clk_i);
a_mant0 = 8'd1; a_mant1 = 8'd135; a_mant2 = 8'd86; a_mant3 = 8'd26;
b_mant0 = 8'd127; b_mant1 = 8'd110; b_mant2 = 8'd89; b_mant3 = 8'd152;
a_exp0 = 10'd43; a_exp1 = 10'd375; a_exp2 = 10'd417; a_exp3 = 10'd339;
b_exp0 = 10'd346; b_exp1 = 10'd943; b_exp2 = 10'd799; b_exp3 = 10'd182;
a_sign0 = 4'd8; a_sign1 = 4'd12; a_sign2 = 4'd13; a_sign3 = 4'd8;
b_sign0 = 4'd12; b_sign1 = 4'd9; b_sign2 = 4'd12; b_sign3 = 4'd6;
@(posedge clk_i);
a_mant0 = 8'd150; a_mant1 = 8'd238; a_mant2 = 8'd80; a_mant3 = 8'd85;
b_mant0 = 8'd143; b_mant1 = 8'd32; b_mant2 = 8'd103; b_mant3 = 8'd220;
a_exp0 = 10'd953; a_exp1 = 10'd436; a_exp2 = 10'd440; a_exp3 = 10'd356;
b_exp0 = 10'd782; b_exp1 = 10'd536; b_exp2 = 10'd581; b_exp3 = 10'd271;
a_sign0 = 4'd15; a_sign1 = 4'd0; a_sign2 = 4'd3; a_sign3 = 4'd8;
b_sign0 = 4'd5; b_sign1 = 4'd12; b_sign2 = 4'd7; b_sign3 = 4'd16;
@(posedge clk_i);
a_mant0 = 8'd122; a_mant1 = 8'd90; a_mant2 = 8'd110; a_mant3 = 8'd234;
b_mant0 = 8'd190; b_mant1 = 8'd181; b_mant2 = 8'd168; b_mant3 = 8'd76;
a_exp0 = 10'd547; a_exp1 = 10'd922; a_exp2 = 10'd209; a_exp3 = 10'd534;
b_exp0 = 10'd933; b_exp1 = 10'd332; b_exp2 = 10'd57; b_exp3 = 10'd760;
a_sign0 = 4'd13; a_sign1 = 4'd7; a_sign2 = 4'd12; a_sign3 = 4'd5;
b_sign0 = 4'd5; b_sign1 = 4'd16; b_sign2 = 4'd7; b_sign3 = 4'd10;
@(posedge clk_i);
a_mant0 = 8'd31; a_mant1 = 8'd42; a_mant2 = 8'd140; a_mant3 = 8'd26;
b_mant0 = 8'd19; b_mant1 = 8'd228; b_mant2 = 8'd9; b_mant3 = 8'd211;
a_exp0 = 10'd47; a_exp1 = 10'd512; a_exp2 = 10'd201; a_exp3 = 10'd653;
b_exp0 = 10'd642; b_exp1 = 10'd240; b_exp2 = 10'd911; b_exp3 = 10'd99;
a_sign0 = 4'd15; a_sign1 = 4'd16; a_sign2 = 4'd1; a_sign3 = 4'd1;
b_sign0 = 4'd13; b_sign1 = 4'd3; b_sign2 = 4'd7; b_sign3 = 4'd16;
@(posedge clk_i);
a_mant0 = 8'd222; a_mant1 = 8'd221; a_mant2 = 8'd180; a_mant3 = 8'd247;
b_mant0 = 8'd111; b_mant1 = 8'd145; b_mant2 = 8'd204; b_mant3 = 8'd145;
a_exp0 = 10'd538; a_exp1 = 10'd29; a_exp2 = 10'd497; a_exp3 = 10'd22;
b_exp0 = 10'd295; b_exp1 = 10'd629; b_exp2 = 10'd105; b_exp3 = 10'd139;
a_sign0 = 4'd4; a_sign1 = 4'd13; a_sign2 = 4'd15; a_sign3 = 4'd15;
b_sign0 = 4'd1; b_sign1 = 4'd16; b_sign2 = 4'd16; b_sign3 = 4'd1;
@(posedge clk_i);
a_mant0 = 8'd77; a_mant1 = 8'd130; a_mant2 = 8'd183; a_mant3 = 8'd76;
b_mant0 = 8'd181; b_mant1 = 8'd75; b_mant2 = 8'd195; b_mant3 = 8'd16;
a_exp0 = 10'd677; a_exp1 = 10'd581; a_exp2 = 10'd449; a_exp3 = 10'd297;
b_exp0 = 10'd309; b_exp1 = 10'd280; b_exp2 = 10'd376; b_exp3 = 10'd587;
a_sign0 = 4'd11; a_sign1 = 4'd7; a_sign2 = 4'd12; a_sign3 = 4'd4;
b_sign0 = 4'd2; b_sign1 = 4'd12; b_sign2 = 4'd14; b_sign3 = 4'd4;
@(posedge clk_i);
shared_exps0 = 8'd111;
shared_exps1 = 8'd145;
a_mant0 = 8'd234; a_mant1 = 8'd105; a_mant2 = 8'd96; a_mant3 = 8'd213;
b_mant0 = 8'd32; b_mant1 = 8'd95; b_mant2 = 8'd60; b_mant3 = 8'd34;
a_exp0 = 10'd374; a_exp1 = 10'd705; a_exp2 = 10'd784; a_exp3 = 10'd276;
b_exp0 = 10'd938; b_exp1 = 10'd482; b_exp2 = 10'd681; b_exp3 = 10'd778;
a_sign0 = 4'd12; a_sign1 = 4'd0; a_sign2 = 4'd14; a_sign3 = 4'd16;
b_sign0 = 4'd15; b_sign1 = 4'd3; b_sign2 = 4'd16; b_sign3 = 4'd12;
@(posedge clk_i);
a_mant0 = 8'd10; a_mant1 = 8'd1; a_mant2 = 8'd94; a_mant3 = 8'd16;
b_mant0 = 8'd28; b_mant1 = 8'd120; b_mant2 = 8'd120; b_mant3 = 8'd15;
a_exp0 = 10'd506; a_exp1 = 10'd294; a_exp2 = 10'd436; a_exp3 = 10'd619;
b_exp0 = 10'd225; b_exp1 = 10'd738; b_exp2 = 10'd587; b_exp3 = 10'd289;
a_sign0 = 4'd10; a_sign1 = 4'd2; a_sign2 = 4'd5; a_sign3 = 4'd2;
b_sign0 = 4'd13; b_sign1 = 4'd9; b_sign2 = 4'd1; b_sign3 = 4'd0;
@(posedge clk_i);
a_mant0 = 8'd122; a_mant1 = 8'd113; a_mant2 = 8'd203; a_mant3 = 8'd57;
b_mant0 = 8'd199; b_mant1 = 8'd163; b_mant2 = 8'd219; b_mant3 = 8'd248;
a_exp0 = 10'd851; a_exp1 = 10'd449; a_exp2 = 10'd224; a_exp3 = 10'd815;
b_exp0 = 10'd706; b_exp1 = 10'd836; b_exp2 = 10'd812; b_exp3 = 10'd35;
a_sign0 = 4'd2; a_sign1 = 4'd9; a_sign2 = 4'd13; a_sign3 = 4'd10;
b_sign0 = 4'd8; b_sign1 = 4'd13; b_sign2 = 4'd5; b_sign3 = 4'd9;
@(posedge clk_i);
a_mant0 = 8'd99; a_mant1 = 8'd108; a_mant2 = 8'd46; a_mant3 = 8'd152;
b_mant0 = 8'd249; b_mant1 = 8'd29; b_mant2 = 8'd254; b_mant3 = 8'd154;
a_exp0 = 10'd679; a_exp1 = 10'd366; a_exp2 = 10'd923; a_exp3 = 10'd287;
b_exp0 = 10'd880; b_exp1 = 10'd254; b_exp2 = 10'd44; b_exp3 = 10'd192;
a_sign0 = 4'd7; a_sign1 = 4'd1; a_sign2 = 4'd13; a_sign3 = 4'd15;
b_sign0 = 4'd12; b_sign1 = 4'd7; b_sign2 = 4'd11; b_sign3 = 4'd10;
@(posedge clk_i);
a_mant0 = 8'd177; a_mant1 = 8'd186; a_mant2 = 8'd217; a_mant3 = 8'd215;
b_mant0 = 8'd150; b_mant1 = 8'd12; b_mant2 = 8'd134; b_mant3 = 8'd0;
a_exp0 = 10'd841; a_exp1 = 10'd67; a_exp2 = 10'd539; a_exp3 = 10'd705;
b_exp0 = 10'd205; b_exp1 = 10'd636; b_exp2 = 10'd774; b_exp3 = 10'd475;
a_sign0 = 4'd15; a_sign1 = 4'd9; a_sign2 = 4'd9; a_sign3 = 4'd2;
b_sign0 = 4'd13; b_sign1 = 4'd10; b_sign2 = 4'd0; b_sign3 = 4'd10;
@(posedge clk_i);
a_mant0 = 8'd119; a_mant1 = 8'd167; a_mant2 = 8'd4; a_mant3 = 8'd28;
b_mant0 = 8'd47; b_mant1 = 8'd100; b_mant2 = 8'd214; b_mant3 = 8'd91;
a_exp0 = 10'd550; a_exp1 = 10'd684; a_exp2 = 10'd561; a_exp3 = 10'd315;
b_exp0 = 10'd983; b_exp1 = 10'd33; b_exp2 = 10'd180; b_exp3 = 10'd555;
a_sign0 = 4'd7; a_sign1 = 4'd0; a_sign2 = 4'd12; a_sign3 = 4'd3;
b_sign0 = 4'd8; b_sign1 = 4'd0; b_sign2 = 4'd0; b_sign3 = 4'd3;
@(posedge clk_i);
a_mant0 = 8'd129; a_mant1 = 8'd112; a_mant2 = 8'd244; a_mant3 = 8'd44;
b_mant0 = 8'd161; b_mant1 = 8'd78; b_mant2 = 8'd22; b_mant3 = 8'd88;
a_exp0 = 10'd757; a_exp1 = 10'd943; a_exp2 = 10'd238; a_exp3 = 10'd188;
b_exp0 = 10'd620; b_exp1 = 10'd759; b_exp2 = 10'd102; b_exp3 = 10'd622;
a_sign0 = 4'd15; a_sign1 = 4'd6; a_sign2 = 4'd11; a_sign3 = 4'd3;
b_sign0 = 4'd2; b_sign1 = 4'd3; b_sign2 = 4'd8; b_sign3 = 4'd11;
@(posedge clk_i);
a_mant0 = 8'd59; a_mant1 = 8'd251; a_mant2 = 8'd38; a_mant3 = 8'd24;
b_mant0 = 8'd217; b_mant1 = 8'd95; b_mant2 = 8'd174; b_mant3 = 8'd35;
a_exp0 = 10'd821; a_exp1 = 10'd739; a_exp2 = 10'd523; a_exp3 = 10'd208;
b_exp0 = 10'd73; b_exp1 = 10'd562; b_exp2 = 10'd103; b_exp3 = 10'd944;
a_sign0 = 4'd11; a_sign1 = 4'd4; a_sign2 = 4'd1; a_sign3 = 4'd5;
b_sign0 = 4'd11; b_sign1 = 4'd6; b_sign2 = 4'd8; b_sign3 = 4'd11;
@(posedge clk_i);
shared_exps0 = 8'd147;
shared_exps1 = 8'd96;
a_mant0 = 8'd49; a_mant1 = 8'd101; a_mant2 = 8'd55; a_mant3 = 8'd86;
b_mant0 = 8'd65; b_mant1 = 8'd116; b_mant2 = 8'd139; b_mant3 = 8'd177;
a_exp0 = 10'd798; a_exp1 = 10'd267; a_exp2 = 10'd558; a_exp3 = 10'd939;
b_exp0 = 10'd483; b_exp1 = 10'd483; b_exp2 = 10'd992; b_exp3 = 10'd577;
a_sign0 = 4'd16; a_sign1 = 4'd15; a_sign2 = 4'd3; a_sign3 = 4'd9;
b_sign0 = 4'd10; b_sign1 = 4'd0; b_sign2 = 4'd16; b_sign3 = 4'd16;
@(posedge clk_i);
a_mant0 = 8'd20; a_mant1 = 8'd241; a_mant2 = 8'd25; a_mant3 = 8'd82;
b_mant0 = 8'd184; b_mant1 = 8'd117; b_mant2 = 8'd132; b_mant3 = 8'd66;
a_exp0 = 10'd540; a_exp1 = 10'd178; a_exp2 = 10'd663; a_exp3 = 10'd502;
b_exp0 = 10'd609; b_exp1 = 10'd842; b_exp2 = 10'd736; b_exp3 = 10'd847;
a_sign0 = 4'd10; a_sign1 = 4'd8; a_sign2 = 4'd13; a_sign3 = 4'd0;
b_sign0 = 4'd12; b_sign1 = 4'd13; b_sign2 = 4'd16; b_sign3 = 4'd14;
@(posedge clk_i);
a_mant0 = 8'd133; a_mant1 = 8'd161; a_mant2 = 8'd99; a_mant3 = 8'd83;
b_mant0 = 8'd223; b_mant1 = 8'd138; b_mant2 = 8'd85; b_mant3 = 8'd206;
a_exp0 = 10'd934; a_exp1 = 10'd454; a_exp2 = 10'd180; a_exp3 = 10'd924;
b_exp0 = 10'd908; b_exp1 = 10'd337; b_exp2 = 10'd267; b_exp3 = 10'd39;
a_sign0 = 4'd13; a_sign1 = 4'd15; a_sign2 = 4'd11; a_sign3 = 4'd6;
b_sign0 = 4'd11; b_sign1 = 4'd14; b_sign2 = 4'd9; b_sign3 = 4'd9;
@(posedge clk_i);
a_mant0 = 8'd98; a_mant1 = 8'd121; a_mant2 = 8'd14; a_mant3 = 8'd169;
b_mant0 = 8'd227; b_mant1 = 8'd141; b_mant2 = 8'd98; b_mant3 = 8'd139;
a_exp0 = 10'd54; a_exp1 = 10'd687; a_exp2 = 10'd759; a_exp3 = 10'd946;
b_exp0 = 10'd95; b_exp1 = 10'd231; b_exp2 = 10'd548; b_exp3 = 10'd980;
a_sign0 = 4'd10; a_sign1 = 4'd15; a_sign2 = 4'd7; a_sign3 = 4'd13;
b_sign0 = 4'd16; b_sign1 = 4'd10; b_sign2 = 4'd5; b_sign3 = 4'd8;
@(posedge clk_i);
a_mant0 = 8'd190; a_mant1 = 8'd47; a_mant2 = 8'd206; a_mant3 = 8'd116;
b_mant0 = 8'd135; b_mant1 = 8'd24; b_mant2 = 8'd193; b_mant3 = 8'd145;
a_exp0 = 10'd804; a_exp1 = 10'd35; a_exp2 = 10'd402; a_exp3 = 10'd970;
b_exp0 = 10'd147; b_exp1 = 10'd104; b_exp2 = 10'd109; b_exp3 = 10'd990;
a_sign0 = 4'd9; a_sign1 = 4'd2; a_sign2 = 4'd8; a_sign3 = 4'd8;
b_sign0 = 4'd5; b_sign1 = 4'd5; b_sign2 = 4'd8; b_sign3 = 4'd6;
@(posedge clk_i);
a_mant0 = 8'd237; a_mant1 = 8'd137; a_mant2 = 8'd154; a_mant3 = 8'd205;
b_mant0 = 8'd14; b_mant1 = 8'd157; b_mant2 = 8'd203; b_mant3 = 8'd187;
a_exp0 = 10'd799; a_exp1 = 10'd768; a_exp2 = 10'd966; a_exp3 = 10'd358;
b_exp0 = 10'd683; b_exp1 = 10'd890; b_exp2 = 10'd1017; b_exp3 = 10'd776;
a_sign0 = 4'd4; a_sign1 = 4'd0; a_sign2 = 4'd11; a_sign3 = 4'd4;
b_sign0 = 4'd15; b_sign1 = 4'd1; b_sign2 = 4'd7; b_sign3 = 4'd5;
@(posedge clk_i);
a_mant0 = 8'd30; a_mant1 = 8'd33; a_mant2 = 8'd63; a_mant3 = 8'd160;
b_mant0 = 8'd145; b_mant1 = 8'd230; b_mant2 = 8'd24; b_mant3 = 8'd248;
a_exp0 = 10'd733; a_exp1 = 10'd268; a_exp2 = 10'd993; a_exp3 = 10'd1023;
b_exp0 = 10'd37; b_exp1 = 10'd289; b_exp2 = 10'd576; b_exp3 = 10'd49;
a_sign0 = 4'd1; a_sign1 = 4'd8; a_sign2 = 4'd2; a_sign3 = 4'd11;
b_sign0 = 4'd1; b_sign1 = 4'd9; b_sign2 = 4'd16; b_sign3 = 4'd6;
@(posedge clk_i);
a_mant0 = 8'd88; a_mant1 = 8'd8; a_mant2 = 8'd107; a_mant3 = 8'd2;
b_mant0 = 8'd116; b_mant1 = 8'd157; b_mant2 = 8'd27; b_mant3 = 8'd38;
a_exp0 = 10'd978; a_exp1 = 10'd905; a_exp2 = 10'd31; a_exp3 = 10'd85;
b_exp0 = 10'd418; b_exp1 = 10'd687; b_exp2 = 10'd812; b_exp3 = 10'd58;
a_sign0 = 4'd11; a_sign1 = 4'd4; a_sign2 = 4'd13; a_sign3 = 4'd3;
b_sign0 = 4'd13; b_sign1 = 4'd15; b_sign2 = 4'd0; b_sign3 = 4'd14;
@(posedge clk_i);
shared_exps0 = 8'd135;
shared_exps1 = 8'd119;
rstn = 0;
@(posedge clk_i);
rstn = 1;
a_mant0 = 8'd66; a_mant1 = 8'd224; a_mant2 = 8'd198; a_mant3 = 8'd125;
b_mant0 = 8'd224; b_mant1 = 8'd248; b_mant2 = 8'd193; b_mant3 = 8'd60;
a_exp0 = 10'd593; a_exp1 = 10'd891; a_exp2 = 10'd487; a_exp3 = 10'd1017;
b_exp0 = 10'd585; b_exp1 = 10'd103; b_exp2 = 10'd267; b_exp3 = 10'd454;
a_sign0 = 4'd5; a_sign1 = 4'd0; a_sign2 = 4'd2; a_sign3 = 4'd3;
b_sign0 = 4'd2; b_sign1 = 4'd0; b_sign2 = 4'd1; b_sign3 = 4'd8;
@(posedge clk_i);
a_mant0 = 8'd33; a_mant1 = 8'd219; a_mant2 = 8'd213; a_mant3 = 8'd143;
b_mant0 = 8'd71; b_mant1 = 8'd5; b_mant2 = 8'd162; b_mant3 = 8'd183;
a_exp0 = 10'd449; a_exp1 = 10'd903; a_exp2 = 10'd639; a_exp3 = 10'd752;
b_exp0 = 10'd803; b_exp1 = 10'd150; b_exp2 = 10'd638; b_exp3 = 10'd913;
a_sign0 = 4'd5; a_sign1 = 4'd11; a_sign2 = 4'd15; a_sign3 = 4'd12;
b_sign0 = 4'd13; b_sign1 = 4'd0; b_sign2 = 4'd4; b_sign3 = 4'd4;
@(posedge clk_i);
a_mant0 = 8'd202; a_mant1 = 8'd14; a_mant2 = 8'd87; a_mant3 = 8'd205;
b_mant0 = 8'd157; b_mant1 = 8'd136; b_mant2 = 8'd172; b_mant3 = 8'd1;
a_exp0 = 10'd296; a_exp1 = 10'd802; a_exp2 = 10'd665; a_exp3 = 10'd599;
b_exp0 = 10'd850; b_exp1 = 10'd16; b_exp2 = 10'd601; b_exp3 = 10'd44;
a_sign0 = 4'd8; a_sign1 = 4'd11; a_sign2 = 4'd11; a_sign3 = 4'd15;
b_sign0 = 4'd14; b_sign1 = 4'd2; b_sign2 = 4'd1; b_sign3 = 4'd4;
@(posedge clk_i);
a_mant0 = 8'd98; a_mant1 = 8'd21; a_mant2 = 8'd51; a_mant3 = 8'd1;
b_mant0 = 8'd37; b_mant1 = 8'd162; b_mant2 = 8'd110; b_mant3 = 8'd171;
a_exp0 = 10'd273; a_exp1 = 10'd1005; a_exp2 = 10'd534; a_exp3 = 10'd912;
b_exp0 = 10'd286; b_exp1 = 10'd570; b_exp2 = 10'd394; b_exp3 = 10'd863;
a_sign0 = 4'd4; a_sign1 = 4'd10; a_sign2 = 4'd2; a_sign3 = 4'd14;
b_sign0 = 4'd0; b_sign1 = 4'd1; b_sign2 = 4'd16; b_sign3 = 4'd9;
@(posedge clk_i);
a_mant0 = 8'd221; a_mant1 = 8'd57; a_mant2 = 8'd193; a_mant3 = 8'd184;
b_mant0 = 8'd125; b_mant1 = 8'd108; b_mant2 = 8'd56; b_mant3 = 8'd119;
a_exp0 = 10'd537; a_exp1 = 10'd276; a_exp2 = 10'd866; a_exp3 = 10'd661;
b_exp0 = 10'd763; b_exp1 = 10'd289; b_exp2 = 10'd758; b_exp3 = 10'd240;
a_sign0 = 4'd12; a_sign1 = 4'd15; a_sign2 = 4'd2; a_sign3 = 4'd2;
b_sign0 = 4'd12; b_sign1 = 4'd0; b_sign2 = 4'd14; b_sign3 = 4'd13;
@(posedge clk_i);
a_mant0 = 8'd18; a_mant1 = 8'd2; a_mant2 = 8'd56; a_mant3 = 8'd195;
b_mant0 = 8'd56; b_mant1 = 8'd65; b_mant2 = 8'd30; b_mant3 = 8'd194;
a_exp0 = 10'd379; a_exp1 = 10'd369; a_exp2 = 10'd213; a_exp3 = 10'd662;
b_exp0 = 10'd776; b_exp1 = 10'd869; b_exp2 = 10'd936; b_exp3 = 10'd200;
a_sign0 = 4'd8; a_sign1 = 4'd4; a_sign2 = 4'd6; a_sign3 = 4'd7;
b_sign0 = 4'd3; b_sign1 = 4'd10; b_sign2 = 4'd10; b_sign3 = 4'd6;
@(posedge clk_i);
a_mant0 = 8'd87; a_mant1 = 8'd38; a_mant2 = 8'd103; a_mant3 = 8'd220;
b_mant0 = 8'd131; b_mant1 = 8'd151; b_mant2 = 8'd122; b_mant3 = 8'd22;
a_exp0 = 10'd104; a_exp1 = 10'd66; a_exp2 = 10'd30; a_exp3 = 10'd234;
b_exp0 = 10'd8; b_exp1 = 10'd14; b_exp2 = 10'd813; b_exp3 = 10'd260;
a_sign0 = 4'd6; a_sign1 = 4'd8; a_sign2 = 4'd3; a_sign3 = 4'd0;
b_sign0 = 4'd0; b_sign1 = 4'd1; b_sign2 = 4'd4; b_sign3 = 4'd5;
@(posedge clk_i);
shared_exps0 = 8'd130;
shared_exps1 = 8'd155;
a_mant0 = 8'd82; a_mant1 = 8'd6; a_mant2 = 8'd234; a_mant3 = 8'd118;
b_mant0 = 8'd146; b_mant1 = 8'd180; b_mant2 = 8'd76; b_mant3 = 8'd111;
a_exp0 = 10'd21; a_exp1 = 10'd116; a_exp2 = 10'd948; a_exp3 = 10'd837;
b_exp0 = 10'd435; b_exp1 = 10'd345; b_exp2 = 10'd78; b_exp3 = 10'd683;
a_sign0 = 4'd3; a_sign1 = 4'd10; a_sign2 = 4'd16; a_sign3 = 4'd0;
b_sign0 = 4'd16; b_sign1 = 4'd8; b_sign2 = 4'd3; b_sign3 = 4'd3;
@(posedge clk_i);
a_mant0 = 8'd182; a_mant1 = 8'd43; a_mant2 = 8'd121; a_mant3 = 8'd232;
b_mant0 = 8'd158; b_mant1 = 8'd230; b_mant2 = 8'd206; b_mant3 = 8'd61;
a_exp0 = 10'd435; a_exp1 = 10'd625; a_exp2 = 10'd618; a_exp3 = 10'd212;
b_exp0 = 10'd586; b_exp1 = 10'd181; b_exp2 = 10'd493; b_exp3 = 10'd416;
a_sign0 = 4'd4; a_sign1 = 4'd13; a_sign2 = 4'd12; a_sign3 = 4'd1;
b_sign0 = 4'd3; b_sign1 = 4'd14; b_sign2 = 4'd11; b_sign3 = 4'd9;
@(posedge clk_i);
a_mant0 = 8'd34; a_mant1 = 8'd163; a_mant2 = 8'd26; a_mant3 = 8'd224;
b_mant0 = 8'd149; b_mant1 = 8'd99; b_mant2 = 8'd253; b_mant3 = 8'd80;
a_exp0 = 10'd650; a_exp1 = 10'd314; a_exp2 = 10'd329; a_exp3 = 10'd1009;
b_exp0 = 10'd959; b_exp1 = 10'd973; b_exp2 = 10'd376; b_exp3 = 10'd943;
a_sign0 = 4'd10; a_sign1 = 4'd6; a_sign2 = 4'd15; a_sign3 = 4'd6;
b_sign0 = 4'd3; b_sign1 = 4'd6; b_sign2 = 4'd10; b_sign3 = 4'd6;
@(posedge clk_i);
a_mant0 = 8'd225; a_mant1 = 8'd133; a_mant2 = 8'd80; a_mant3 = 8'd220;
b_mant0 = 8'd182; b_mant1 = 8'd241; b_mant2 = 8'd2; b_mant3 = 8'd243;
a_exp0 = 10'd623; a_exp1 = 10'd359; a_exp2 = 10'd109; a_exp3 = 10'd757;
b_exp0 = 10'd700; b_exp1 = 10'd468; b_exp2 = 10'd455; b_exp3 = 10'd815;
a_sign0 = 4'd0; a_sign1 = 4'd8; a_sign2 = 4'd4; a_sign3 = 4'd7;
b_sign0 = 4'd0; b_sign1 = 4'd2; b_sign2 = 4'd14; b_sign3 = 4'd3;
@(posedge clk_i);
a_mant0 = 8'd221; a_mant1 = 8'd128; a_mant2 = 8'd171; a_mant3 = 8'd128;
b_mant0 = 8'd194; b_mant1 = 8'd197; b_mant2 = 8'd25; b_mant3 = 8'd73;
a_exp0 = 10'd366; a_exp1 = 10'd911; a_exp2 = 10'd577; a_exp3 = 10'd197;
b_exp0 = 10'd712; b_exp1 = 10'd803; b_exp2 = 10'd725; b_exp3 = 10'd957;
a_sign0 = 4'd9; a_sign1 = 4'd16; a_sign2 = 4'd11; a_sign3 = 4'd7;
b_sign0 = 4'd4; b_sign1 = 4'd8; b_sign2 = 4'd12; b_sign3 = 4'd0;
@(posedge clk_i);
a_mant0 = 8'd9; a_mant1 = 8'd2; a_mant2 = 8'd239; a_mant3 = 8'd60;
b_mant0 = 8'd255; b_mant1 = 8'd249; b_mant2 = 8'd15; b_mant3 = 8'd63;
a_exp0 = 10'd522; a_exp1 = 10'd314; a_exp2 = 10'd283; a_exp3 = 10'd604;
b_exp0 = 10'd878; b_exp1 = 10'd707; b_exp2 = 10'd86; b_exp3 = 10'd511;
a_sign0 = 4'd9; a_sign1 = 4'd9; a_sign2 = 4'd15; a_sign3 = 4'd15;
b_sign0 = 4'd10; b_sign1 = 4'd11; b_sign2 = 4'd11; b_sign3 = 4'd6;
@(posedge clk_i);
a_mant0 = 8'd13; a_mant1 = 8'd126; a_mant2 = 8'd208; a_mant3 = 8'd150;
b_mant0 = 8'd115; b_mant1 = 8'd23; b_mant2 = 8'd184; b_mant3 = 8'd161;
a_exp0 = 10'd942; a_exp1 = 10'd391; a_exp2 = 10'd270; a_exp3 = 10'd550;
b_exp0 = 10'd126; b_exp1 = 10'd999; b_exp2 = 10'd277; b_exp3 = 10'd925;
a_sign0 = 4'd4; a_sign1 = 4'd13; a_sign2 = 4'd1; a_sign3 = 4'd13;
b_sign0 = 4'd6; b_sign1 = 4'd4; b_sign2 = 4'd14; b_sign3 = 4'd14;
@(posedge clk_i);
a_mant0 = 8'd135; a_mant1 = 8'd151; a_mant2 = 8'd148; a_mant3 = 8'd149;
b_mant0 = 8'd47; b_mant1 = 8'd25; b_mant2 = 8'd199; b_mant3 = 8'd224;
a_exp0 = 10'd623; a_exp1 = 10'd589; a_exp2 = 10'd270; a_exp3 = 10'd784;
b_exp0 = 10'd279; b_exp1 = 10'd742; b_exp2 = 10'd355; b_exp3 = 10'd318;
a_sign0 = 4'd15; a_sign1 = 4'd1; a_sign2 = 4'd7; a_sign3 = 4'd10;
b_sign0 = 4'd6; b_sign1 = 4'd11; b_sign2 = 4'd1; b_sign3 = 4'd6;
@(posedge clk_i);
shared_exps0 = 8'd147;
shared_exps1 = 8'd118;
a_mant0 = 8'd24; a_mant1 = 8'd133; a_mant2 = 8'd72; a_mant3 = 8'd4;
b_mant0 = 8'd77; b_mant1 = 8'd1; b_mant2 = 8'd43; b_mant3 = 8'd2;
a_exp0 = 10'd85; a_exp1 = 10'd271; a_exp2 = 10'd107; a_exp3 = 10'd274;
b_exp0 = 10'd490; b_exp1 = 10'd23; b_exp2 = 10'd473; b_exp3 = 10'd29;
a_sign0 = 4'd0; a_sign1 = 4'd3; a_sign2 = 4'd11; a_sign3 = 4'd9;
b_sign0 = 4'd11; b_sign1 = 4'd2; b_sign2 = 4'd4; b_sign3 = 4'd9;
@(posedge clk_i);
a_mant0 = 8'd70; a_mant1 = 8'd232; a_mant2 = 8'd215; a_mant3 = 8'd79;
b_mant0 = 8'd66; b_mant1 = 8'd127; b_mant2 = 8'd14; b_mant3 = 8'd95;
a_exp0 = 10'd682; a_exp1 = 10'd572; a_exp2 = 10'd823; a_exp3 = 10'd243;
b_exp0 = 10'd959; b_exp1 = 10'd262; b_exp2 = 10'd62; b_exp3 = 10'd755;
a_sign0 = 4'd7; a_sign1 = 4'd1; a_sign2 = 4'd12; a_sign3 = 4'd3;
b_sign0 = 4'd15; b_sign1 = 4'd11; b_sign2 = 4'd15; b_sign3 = 4'd15;
@(posedge clk_i);
a_mant0 = 8'd149; a_mant1 = 8'd169; a_mant2 = 8'd112; a_mant3 = 8'd74;
b_mant0 = 8'd199; b_mant1 = 8'd168; b_mant2 = 8'd207; b_mant3 = 8'd113;
a_exp0 = 10'd169; a_exp1 = 10'd943; a_exp2 = 10'd766; a_exp3 = 10'd137;
b_exp0 = 10'd962; b_exp1 = 10'd42; b_exp2 = 10'd81; b_exp3 = 10'd285;
a_sign0 = 4'd3; a_sign1 = 4'd0; a_sign2 = 4'd8; a_sign3 = 4'd8;
b_sign0 = 4'd14; b_sign1 = 4'd11; b_sign2 = 4'd9; b_sign3 = 4'd0;
@(posedge clk_i);
a_mant0 = 8'd19; a_mant1 = 8'd196; a_mant2 = 8'd77; a_mant3 = 8'd63;
b_mant0 = 8'd219; b_mant1 = 8'd35; b_mant2 = 8'd12; b_mant3 = 8'd110;
a_exp0 = 10'd837; a_exp1 = 10'd439; a_exp2 = 10'd207; a_exp3 = 10'd898;
b_exp0 = 10'd753; b_exp1 = 10'd470; b_exp2 = 10'd653; b_exp3 = 10'd301;
a_sign0 = 4'd15; a_sign1 = 4'd11; a_sign2 = 4'd15; a_sign3 = 4'd7;
b_sign0 = 4'd1; b_sign1 = 4'd14; b_sign2 = 4'd8; b_sign3 = 4'd12;
@(posedge clk_i);
a_mant0 = 8'd140; a_mant1 = 8'd142; a_mant2 = 8'd19; a_mant3 = 8'd196;
b_mant0 = 8'd78; b_mant1 = 8'd177; b_mant2 = 8'd83; b_mant3 = 8'd88;
a_exp0 = 10'd817; a_exp1 = 10'd718; a_exp2 = 10'd961; a_exp3 = 10'd687;
b_exp0 = 10'd747; b_exp1 = 10'd983; b_exp2 = 10'd920; b_exp3 = 10'd916;
a_sign0 = 4'd15; a_sign1 = 4'd2; a_sign2 = 4'd2; a_sign3 = 4'd14;
b_sign0 = 4'd13; b_sign1 = 4'd7; b_sign2 = 4'd11; b_sign3 = 4'd10;
@(posedge clk_i);
a_mant0 = 8'd57; a_mant1 = 8'd50; a_mant2 = 8'd122; a_mant3 = 8'd18;
b_mant0 = 8'd64; b_mant1 = 8'd108; b_mant2 = 8'd206; b_mant3 = 8'd152;
a_exp0 = 10'd271; a_exp1 = 10'd924; a_exp2 = 10'd449; a_exp3 = 10'd302;
b_exp0 = 10'd540; b_exp1 = 10'd930; b_exp2 = 10'd704; b_exp3 = 10'd152;
a_sign0 = 4'd16; a_sign1 = 4'd12; a_sign2 = 4'd14; a_sign3 = 4'd13;
b_sign0 = 4'd11; b_sign1 = 4'd12; b_sign2 = 4'd9; b_sign3 = 4'd1;
@(posedge clk_i);
a_mant0 = 8'd177; a_mant1 = 8'd166; a_mant2 = 8'd241; a_mant3 = 8'd36;
b_mant0 = 8'd142; b_mant1 = 8'd184; b_mant2 = 8'd92; b_mant3 = 8'd235;
a_exp0 = 10'd942; a_exp1 = 10'd141; a_exp2 = 10'd344; a_exp3 = 10'd26;
b_exp0 = 10'd423; b_exp1 = 10'd760; b_exp2 = 10'd35; b_exp3 = 10'd874;
a_sign0 = 4'd12; a_sign1 = 4'd4; a_sign2 = 4'd13; a_sign3 = 4'd2;
b_sign0 = 4'd8; b_sign1 = 4'd11; b_sign2 = 4'd10; b_sign3 = 4'd5;
@(posedge clk_i);
a_mant0 = 8'd111; a_mant1 = 8'd51; a_mant2 = 8'd139; a_mant3 = 8'd218;
b_mant0 = 8'd156; b_mant1 = 8'd69; b_mant2 = 8'd36; b_mant3 = 8'd2;
a_exp0 = 10'd541; a_exp1 = 10'd31; a_exp2 = 10'd494; a_exp3 = 10'd197;
b_exp0 = 10'd240; b_exp1 = 10'd701; b_exp2 = 10'd626; b_exp3 = 10'd295;
a_sign0 = 4'd8; a_sign1 = 4'd5; a_sign2 = 4'd0; a_sign3 = 4'd9;
b_sign0 = 4'd10; b_sign1 = 4'd8; b_sign2 = 4'd0; b_sign3 = 4'd8;
@(posedge clk_i);
shared_exps0 = 8'd134;
shared_exps1 = 8'd121;
a_mant0 = 8'd154; a_mant1 = 8'd220; a_mant2 = 8'd169; a_mant3 = 8'd156;
b_mant0 = 8'd149; b_mant1 = 8'd187; b_mant2 = 8'd159; b_mant3 = 8'd128;
a_exp0 = 10'd741; a_exp1 = 10'd692; a_exp2 = 10'd122; a_exp3 = 10'd716;
b_exp0 = 10'd236; b_exp1 = 10'd129; b_exp2 = 10'd861; b_exp3 = 10'd782;
a_sign0 = 4'd0; a_sign1 = 4'd11; a_sign2 = 4'd3; a_sign3 = 4'd9;
b_sign0 = 4'd7; b_sign1 = 4'd6; b_sign2 = 4'd0; b_sign3 = 4'd4;
@(posedge clk_i);
a_mant0 = 8'd63; a_mant1 = 8'd250; a_mant2 = 8'd187; a_mant3 = 8'd196;
b_mant0 = 8'd247; b_mant1 = 8'd23; b_mant2 = 8'd225; b_mant3 = 8'd222;
a_exp0 = 10'd276; a_exp1 = 10'd414; a_exp2 = 10'd75; a_exp3 = 10'd460;
b_exp0 = 10'd475; b_exp1 = 10'd251; b_exp2 = 10'd43; b_exp3 = 10'd274;
a_sign0 = 4'd7; a_sign1 = 4'd15; a_sign2 = 4'd1; a_sign3 = 4'd0;
b_sign0 = 4'd14; b_sign1 = 4'd3; b_sign2 = 4'd0; b_sign3 = 4'd3;
@(posedge clk_i);
a_mant0 = 8'd79; a_mant1 = 8'd190; a_mant2 = 8'd228; a_mant3 = 8'd83;
b_mant0 = 8'd231; b_mant1 = 8'd131; b_mant2 = 8'd126; b_mant3 = 8'd183;
a_exp0 = 10'd687; a_exp1 = 10'd867; a_exp2 = 10'd784; a_exp3 = 10'd444;
b_exp0 = 10'd996; b_exp1 = 10'd801; b_exp2 = 10'd41; b_exp3 = 10'd345;
a_sign0 = 4'd1; a_sign1 = 4'd13; a_sign2 = 4'd13; a_sign3 = 4'd12;
b_sign0 = 4'd3; b_sign1 = 4'd1; b_sign2 = 4'd7; b_sign3 = 4'd13;
@(posedge clk_i);
a_mant0 = 8'd195; a_mant1 = 8'd164; a_mant2 = 8'd155; a_mant3 = 8'd214;
b_mant0 = 8'd34; b_mant1 = 8'd0; b_mant2 = 8'd45; b_mant3 = 8'd35;
a_exp0 = 10'd584; a_exp1 = 10'd819; a_exp2 = 10'd674; a_exp3 = 10'd593;
b_exp0 = 10'd707; b_exp1 = 10'd961; b_exp2 = 10'd671; b_exp3 = 10'd661;
a_sign0 = 4'd1; a_sign1 = 4'd9; a_sign2 = 4'd3; a_sign3 = 4'd12;
b_sign0 = 4'd1; b_sign1 = 4'd9; b_sign2 = 4'd15; b_sign3 = 4'd14;
@(posedge clk_i);
a_mant0 = 8'd214; a_mant1 = 8'd32; a_mant2 = 8'd74; a_mant3 = 8'd150;
b_mant0 = 8'd243; b_mant1 = 8'd156; b_mant2 = 8'd28; b_mant3 = 8'd14;
a_exp0 = 10'd130; a_exp1 = 10'd722; a_exp2 = 10'd722; a_exp3 = 10'd441;
b_exp0 = 10'd651; b_exp1 = 10'd675; b_exp2 = 10'd305; b_exp3 = 10'd800;
a_sign0 = 4'd5; a_sign1 = 4'd16; a_sign2 = 4'd2; a_sign3 = 4'd13;
b_sign0 = 4'd12; b_sign1 = 4'd6; b_sign2 = 4'd16; b_sign3 = 4'd6;
@(posedge clk_i);
a_mant0 = 8'd87; a_mant1 = 8'd181; a_mant2 = 8'd217; a_mant3 = 8'd104;
b_mant0 = 8'd38; b_mant1 = 8'd137; b_mant2 = 8'd140; b_mant3 = 8'd55;
a_exp0 = 10'd96; a_exp1 = 10'd459; a_exp2 = 10'd261; a_exp3 = 10'd224;
b_exp0 = 10'd351; b_exp1 = 10'd367; b_exp2 = 10'd438; b_exp3 = 10'd318;
a_sign0 = 4'd11; a_sign1 = 4'd14; a_sign2 = 4'd4; a_sign3 = 4'd1;
b_sign0 = 4'd3; b_sign1 = 4'd16; b_sign2 = 4'd12; b_sign3 = 4'd7;
@(posedge clk_i);
a_mant0 = 8'd200; a_mant1 = 8'd148; a_mant2 = 8'd98; a_mant3 = 8'd15;
b_mant0 = 8'd238; b_mant1 = 8'd229; b_mant2 = 8'd106; b_mant3 = 8'd99;
a_exp0 = 10'd483; a_exp1 = 10'd149; a_exp2 = 10'd187; a_exp3 = 10'd466;
b_exp0 = 10'd271; b_exp1 = 10'd230; b_exp2 = 10'd23; b_exp3 = 10'd19;
a_sign0 = 4'd10; a_sign1 = 4'd13; a_sign2 = 4'd11; a_sign3 = 4'd6;
b_sign0 = 4'd11; b_sign1 = 4'd0; b_sign2 = 4'd6; b_sign3 = 4'd6;
@(posedge clk_i);
a_mant0 = 8'd1; a_mant1 = 8'd74; a_mant2 = 8'd190; a_mant3 = 8'd20;
b_mant0 = 8'd121; b_mant1 = 8'd169; b_mant2 = 8'd249; b_mant3 = 8'd130;
a_exp0 = 10'd727; a_exp1 = 10'd669; a_exp2 = 10'd956; a_exp3 = 10'd990;
b_exp0 = 10'd362; b_exp1 = 10'd307; b_exp2 = 10'd666; b_exp3 = 10'd407;
a_sign0 = 4'd5; a_sign1 = 4'd6; a_sign2 = 4'd0; a_sign3 = 4'd9;
b_sign0 = 4'd2; b_sign1 = 4'd0; b_sign2 = 4'd16; b_sign3 = 4'd13;
@(posedge clk_i);
shared_exps0 = 8'd109;
shared_exps1 = 8'd150;
rstn = 0;
@(posedge clk_i);
rstn = 1;
a_mant0 = 8'd29; a_mant1 = 8'd109; a_mant2 = 8'd12; a_mant3 = 8'd159;
b_mant0 = 8'd17; b_mant1 = 8'd102; b_mant2 = 8'd236; b_mant3 = 8'd159;
a_exp0 = 10'd979; a_exp1 = 10'd636; a_exp2 = 10'd713; a_exp3 = 10'd527;
b_exp0 = 10'd308; b_exp1 = 10'd267; b_exp2 = 10'd989; b_exp3 = 10'd645;
a_sign0 = 4'd1; a_sign1 = 4'd0; a_sign2 = 4'd2; a_sign3 = 4'd6;
b_sign0 = 4'd3; b_sign1 = 4'd4; b_sign2 = 4'd0; b_sign3 = 4'd3;
@(posedge clk_i);
a_mant0 = 8'd25; a_mant1 = 8'd158; a_mant2 = 8'd183; a_mant3 = 8'd45;
b_mant0 = 8'd228; b_mant1 = 8'd34; b_mant2 = 8'd34; b_mant3 = 8'd168;
a_exp0 = 10'd895; a_exp1 = 10'd1005; a_exp2 = 10'd554; a_exp3 = 10'd630;
b_exp0 = 10'd726; b_exp1 = 10'd865; b_exp2 = 10'd799; b_exp3 = 10'd433;
a_sign0 = 4'd13; a_sign1 = 4'd8; a_sign2 = 4'd13; a_sign3 = 4'd0;
b_sign0 = 4'd1; b_sign1 = 4'd0; b_sign2 = 4'd11; b_sign3 = 4'd13;
@(posedge clk_i);
a_mant0 = 8'd168; a_mant1 = 8'd42; a_mant2 = 8'd79; a_mant3 = 8'd109;
b_mant0 = 8'd221; b_mant1 = 8'd168; b_mant2 = 8'd87; b_mant3 = 8'd64;
a_exp0 = 10'd127; a_exp1 = 10'd674; a_exp2 = 10'd327; a_exp3 = 10'd849;
b_exp0 = 10'd986; b_exp1 = 10'd938; b_exp2 = 10'd1; b_exp3 = 10'd747;
a_sign0 = 4'd0; a_sign1 = 4'd3; a_sign2 = 4'd11; a_sign3 = 4'd2;
b_sign0 = 4'd9; b_sign1 = 4'd15; b_sign2 = 4'd16; b_sign3 = 4'd14;
@(posedge clk_i);
a_mant0 = 8'd34; a_mant1 = 8'd186; a_mant2 = 8'd184; a_mant3 = 8'd108;
b_mant0 = 8'd59; b_mant1 = 8'd159; b_mant2 = 8'd188; b_mant3 = 8'd204;
a_exp0 = 10'd527; a_exp1 = 10'd486; a_exp2 = 10'd631; a_exp3 = 10'd883;
b_exp0 = 10'd753; b_exp1 = 10'd485; b_exp2 = 10'd61; b_exp3 = 10'd744;
a_sign0 = 4'd14; a_sign1 = 4'd0; a_sign2 = 4'd2; a_sign3 = 4'd0;
b_sign0 = 4'd15; b_sign1 = 4'd5; b_sign2 = 4'd10; b_sign3 = 4'd8;
@(posedge clk_i);
a_mant0 = 8'd194; a_mant1 = 8'd16; a_mant2 = 8'd114; a_mant3 = 8'd209;
b_mant0 = 8'd179; b_mant1 = 8'd76; b_mant2 = 8'd78; b_mant3 = 8'd229;
a_exp0 = 10'd436; a_exp1 = 10'd761; a_exp2 = 10'd465; a_exp3 = 10'd227;
b_exp0 = 10'd490; b_exp1 = 10'd1004; b_exp2 = 10'd554; b_exp3 = 10'd453;
a_sign0 = 4'd4; a_sign1 = 4'd14; a_sign2 = 4'd9; a_sign3 = 4'd11;
b_sign0 = 4'd4; b_sign1 = 4'd1; b_sign2 = 4'd10; b_sign3 = 4'd1;
@(posedge clk_i);
a_mant0 = 8'd222; a_mant1 = 8'd33; a_mant2 = 8'd101; a_mant3 = 8'd98;
b_mant0 = 8'd43; b_mant1 = 8'd199; b_mant2 = 8'd77; b_mant3 = 8'd198;
a_exp0 = 10'd269; a_exp1 = 10'd1013; a_exp2 = 10'd148; a_exp3 = 10'd4;
b_exp0 = 10'd771; b_exp1 = 10'd200; b_exp2 = 10'd847; b_exp3 = 10'd823;
a_sign0 = 4'd8; a_sign1 = 4'd6; a_sign2 = 4'd2; a_sign3 = 4'd15;
b_sign0 = 4'd8; b_sign1 = 4'd2; b_sign2 = 4'd0; b_sign3 = 4'd9;
@(posedge clk_i);
a_mant0 = 8'd241; a_mant1 = 8'd148; a_mant2 = 8'd84; a_mant3 = 8'd32;
b_mant0 = 8'd221; b_mant1 = 8'd32; b_mant2 = 8'd74; b_mant3 = 8'd249;
a_exp0 = 10'd633; a_exp1 = 10'd317; a_exp2 = 10'd627; a_exp3 = 10'd353;
b_exp0 = 10'd0; b_exp1 = 10'd626; b_exp2 = 10'd808; b_exp3 = 10'd50;
a_sign0 = 4'd8; a_sign1 = 4'd7; a_sign2 = 4'd0; a_sign3 = 4'd13;
b_sign0 = 4'd8; b_sign1 = 4'd13; b_sign2 = 4'd9; b_sign3 = 4'd10;
@(posedge clk_i);
shared_exps0 = 8'd127;
shared_exps1 = 8'd111;
a_mant0 = 8'd51; a_mant1 = 8'd155; a_mant2 = 8'd249; a_mant3 = 8'd30;
b_mant0 = 8'd28; b_mant1 = 8'd36; b_mant2 = 8'd19; b_mant3 = 8'd192;
a_exp0 = 10'd803; a_exp1 = 10'd698; a_exp2 = 10'd959; a_exp3 = 10'd309;
b_exp0 = 10'd625; b_exp1 = 10'd809; b_exp2 = 10'd220; b_exp3 = 10'd707;
a_sign0 = 4'd0; a_sign1 = 4'd3; a_sign2 = 4'd11; a_sign3 = 4'd4;
b_sign0 = 4'd5; b_sign1 = 4'd15; b_sign2 = 4'd3; b_sign3 = 4'd1;
@(posedge clk_i);
a_mant0 = 8'd201; a_mant1 = 8'd87; a_mant2 = 8'd22; a_mant3 = 8'd93;
b_mant0 = 8'd143; b_mant1 = 8'd148; b_mant2 = 8'd59; b_mant3 = 8'd53;
a_exp0 = 10'd587; a_exp1 = 10'd643; a_exp2 = 10'd478; a_exp3 = 10'd412;
b_exp0 = 10'd198; b_exp1 = 10'd314; b_exp2 = 10'd920; b_exp3 = 10'd890;
a_sign0 = 4'd1; a_sign1 = 4'd15; a_sign2 = 4'd1; a_sign3 = 4'd0;
b_sign0 = 4'd10; b_sign1 = 4'd1; b_sign2 = 4'd5; b_sign3 = 4'd6;
@(posedge clk_i);
a_mant0 = 8'd43; a_mant1 = 8'd231; a_mant2 = 8'd150; a_mant3 = 8'd71;
b_mant0 = 8'd162; b_mant1 = 8'd40; b_mant2 = 8'd176; b_mant3 = 8'd28;
a_exp0 = 10'd348; a_exp1 = 10'd908; a_exp2 = 10'd617; a_exp3 = 10'd551;
b_exp0 = 10'd763; b_exp1 = 10'd246; b_exp2 = 10'd320; b_exp3 = 10'd717;
a_sign0 = 4'd11; a_sign1 = 4'd6; a_sign2 = 4'd1; a_sign3 = 4'd3;
b_sign0 = 4'd1; b_sign1 = 4'd8; b_sign2 = 4'd7; b_sign3 = 4'd0;
@(posedge clk_i);
a_mant0 = 8'd234; a_mant1 = 8'd134; a_mant2 = 8'd54; a_mant3 = 8'd73;
b_mant0 = 8'd11; b_mant1 = 8'd112; b_mant2 = 8'd220; b_mant3 = 8'd93;
a_exp0 = 10'd853; a_exp1 = 10'd366; a_exp2 = 10'd39; a_exp3 = 10'd881;
b_exp0 = 10'd161; b_exp1 = 10'd360; b_exp2 = 10'd682; b_exp3 = 10'd847;
a_sign0 = 4'd15; a_sign1 = 4'd5; a_sign2 = 4'd14; a_sign3 = 4'd5;
b_sign0 = 4'd5; b_sign1 = 4'd3; b_sign2 = 4'd5; b_sign3 = 4'd2;
@(posedge clk_i);
a_mant0 = 8'd56; a_mant1 = 8'd225; a_mant2 = 8'd221; a_mant3 = 8'd46;
b_mant0 = 8'd137; b_mant1 = 8'd79; b_mant2 = 8'd136; b_mant3 = 8'd241;
a_exp0 = 10'd68; a_exp1 = 10'd4; a_exp2 = 10'd443; a_exp3 = 10'd285;
b_exp0 = 10'd924; b_exp1 = 10'd942; b_exp2 = 10'd54; b_exp3 = 10'd662;
a_sign0 = 4'd7; a_sign1 = 4'd11; a_sign2 = 4'd4; a_sign3 = 4'd1;
b_sign0 = 4'd4; b_sign1 = 4'd10; b_sign2 = 4'd0; b_sign3 = 4'd4;
@(posedge clk_i);
a_mant0 = 8'd154; a_mant1 = 8'd203; a_mant2 = 8'd243; a_mant3 = 8'd254;
b_mant0 = 8'd99; b_mant1 = 8'd178; b_mant2 = 8'd112; b_mant3 = 8'd177;
a_exp0 = 10'd158; a_exp1 = 10'd405; a_exp2 = 10'd668; a_exp3 = 10'd239;
b_exp0 = 10'd108; b_exp1 = 10'd826; b_exp2 = 10'd11; b_exp3 = 10'd239;
a_sign0 = 4'd5; a_sign1 = 4'd6; a_sign2 = 4'd9; a_sign3 = 4'd3;
b_sign0 = 4'd7; b_sign1 = 4'd8; b_sign2 = 4'd9; b_sign3 = 4'd0;
@(posedge clk_i);
a_mant0 = 8'd183; a_mant1 = 8'd130; a_mant2 = 8'd40; a_mant3 = 8'd122;
b_mant0 = 8'd208; b_mant1 = 8'd199; b_mant2 = 8'd107; b_mant3 = 8'd182;
a_exp0 = 10'd334; a_exp1 = 10'd875; a_exp2 = 10'd695; a_exp3 = 10'd238;
b_exp0 = 10'd947; b_exp1 = 10'd777; b_exp2 = 10'd224; b_exp3 = 10'd426;
a_sign0 = 4'd3; a_sign1 = 4'd16; a_sign2 = 4'd8; a_sign3 = 4'd5;
b_sign0 = 4'd1; b_sign1 = 4'd16; b_sign2 = 4'd12; b_sign3 = 4'd12;
@(posedge clk_i);
a_mant0 = 8'd112; a_mant1 = 8'd5; a_mant2 = 8'd217; a_mant3 = 8'd223;
b_mant0 = 8'd61; b_mant1 = 8'd82; b_mant2 = 8'd70; b_mant3 = 8'd97;
a_exp0 = 10'd440; a_exp1 = 10'd151; a_exp2 = 10'd295; a_exp3 = 10'd608;
b_exp0 = 10'd487; b_exp1 = 10'd927; b_exp2 = 10'd1003; b_exp3 = 10'd97;
a_sign0 = 4'd0; a_sign1 = 4'd2; a_sign2 = 4'd2; a_sign3 = 4'd8;
b_sign0 = 4'd3; b_sign1 = 4'd16; b_sign2 = 4'd0; b_sign3 = 4'd5;
@(posedge clk_i);
shared_exps0 = 8'd143;
shared_exps1 = 8'd124;
a_mant0 = 8'd33; a_mant1 = 8'd81; a_mant2 = 8'd216; a_mant3 = 8'd189;
b_mant0 = 8'd180; b_mant1 = 8'd156; b_mant2 = 8'd119; b_mant3 = 8'd20;
a_exp0 = 10'd276; a_exp1 = 10'd611; a_exp2 = 10'd668; a_exp3 = 10'd782;
b_exp0 = 10'd461; b_exp1 = 10'd867; b_exp2 = 10'd41; b_exp3 = 10'd987;
a_sign0 = 4'd4; a_sign1 = 4'd10; a_sign2 = 4'd11; a_sign3 = 4'd10;
b_sign0 = 4'd5; b_sign1 = 4'd13; b_sign2 = 4'd13; b_sign3 = 4'd5;
@(posedge clk_i);
a_mant0 = 8'd145; a_mant1 = 8'd100; a_mant2 = 8'd47; a_mant3 = 8'd140;
b_mant0 = 8'd165; b_mant1 = 8'd146; b_mant2 = 8'd197; b_mant3 = 8'd157;
a_exp0 = 10'd968; a_exp1 = 10'd563; a_exp2 = 10'd169; a_exp3 = 10'd99;
b_exp0 = 10'd362; b_exp1 = 10'd386; b_exp2 = 10'd50; b_exp3 = 10'd799;
a_sign0 = 4'd7; a_sign1 = 4'd2; a_sign2 = 4'd11; a_sign3 = 4'd8;
b_sign0 = 4'd15; b_sign1 = 4'd5; b_sign2 = 4'd0; b_sign3 = 4'd2;
@(posedge clk_i);
a_mant0 = 8'd247; a_mant1 = 8'd191; a_mant2 = 8'd188; a_mant3 = 8'd192;
b_mant0 = 8'd40; b_mant1 = 8'd23; b_mant2 = 8'd47; b_mant3 = 8'd28;
a_exp0 = 10'd336; a_exp1 = 10'd342; a_exp2 = 10'd428; a_exp3 = 10'd719;
b_exp0 = 10'd467; b_exp1 = 10'd430; b_exp2 = 10'd506; b_exp3 = 10'd732;
a_sign0 = 4'd7; a_sign1 = 4'd10; a_sign2 = 4'd0; a_sign3 = 4'd9;
b_sign0 = 4'd13; b_sign1 = 4'd10; b_sign2 = 4'd7; b_sign3 = 4'd3;
@(posedge clk_i);
a_mant0 = 8'd181; a_mant1 = 8'd139; a_mant2 = 8'd181; a_mant3 = 8'd248;
b_mant0 = 8'd1; b_mant1 = 8'd187; b_mant2 = 8'd53; b_mant3 = 8'd208;
a_exp0 = 10'd57; a_exp1 = 10'd745; a_exp2 = 10'd587; a_exp3 = 10'd25;
b_exp0 = 10'd831; b_exp1 = 10'd213; b_exp2 = 10'd166; b_exp3 = 10'd765;
a_sign0 = 4'd14; a_sign1 = 4'd6; a_sign2 = 4'd9; a_sign3 = 4'd10;
b_sign0 = 4'd0; b_sign1 = 4'd1; b_sign2 = 4'd8; b_sign3 = 4'd7;
@(posedge clk_i);
a_mant0 = 8'd243; a_mant1 = 8'd18; a_mant2 = 8'd196; a_mant3 = 8'd78;
b_mant0 = 8'd216; b_mant1 = 8'd139; b_mant2 = 8'd80; b_mant3 = 8'd230;
a_exp0 = 10'd596; a_exp1 = 10'd908; a_exp2 = 10'd242; a_exp3 = 10'd533;
b_exp0 = 10'd118; b_exp1 = 10'd837; b_exp2 = 10'd2; b_exp3 = 10'd974;
a_sign0 = 4'd5; a_sign1 = 4'd8; a_sign2 = 4'd9; a_sign3 = 4'd2;
b_sign0 = 4'd3; b_sign1 = 4'd14; b_sign2 = 4'd16; b_sign3 = 4'd8;
@(posedge clk_i);
a_mant0 = 8'd147; a_mant1 = 8'd102; a_mant2 = 8'd17; a_mant3 = 8'd234;
b_mant0 = 8'd62; b_mant1 = 8'd154; b_mant2 = 8'd170; b_mant3 = 8'd5;
a_exp0 = 10'd512; a_exp1 = 10'd673; a_exp2 = 10'd986; a_exp3 = 10'd525;
b_exp0 = 10'd385; b_exp1 = 10'd308; b_exp2 = 10'd948; b_exp3 = 10'd242;
a_sign0 = 4'd5; a_sign1 = 4'd2; a_sign2 = 4'd3; a_sign3 = 4'd1;
b_sign0 = 4'd12; b_sign1 = 4'd15; b_sign2 = 4'd0; b_sign3 = 4'd9;
@(posedge clk_i);
a_mant0 = 8'd198; a_mant1 = 8'd249; a_mant2 = 8'd130; a_mant3 = 8'd120;
b_mant0 = 8'd93; b_mant1 = 8'd131; b_mant2 = 8'd156; b_mant3 = 8'd21;
a_exp0 = 10'd647; a_exp1 = 10'd323; a_exp2 = 10'd81; a_exp3 = 10'd492;
b_exp0 = 10'd140; b_exp1 = 10'd328; b_exp2 = 10'd24; b_exp3 = 10'd408;
a_sign0 = 4'd2; a_sign1 = 4'd12; a_sign2 = 4'd6; a_sign3 = 4'd5;
b_sign0 = 4'd12; b_sign1 = 4'd15; b_sign2 = 4'd8; b_sign3 = 4'd3;
@(posedge clk_i);
a_mant0 = 8'd122; a_mant1 = 8'd212; a_mant2 = 8'd20; a_mant3 = 8'd58;
b_mant0 = 8'd30; b_mant1 = 8'd55; b_mant2 = 8'd63; b_mant3 = 8'd253;
a_exp0 = 10'd769; a_exp1 = 10'd20; a_exp2 = 10'd1010; a_exp3 = 10'd433;
b_exp0 = 10'd862; b_exp1 = 10'd821; b_exp2 = 10'd262; b_exp3 = 10'd986;
a_sign0 = 4'd4; a_sign1 = 4'd10; a_sign2 = 4'd2; a_sign3 = 4'd5;
b_sign0 = 4'd14; b_sign1 = 4'd9; b_sign2 = 4'd11; b_sign3 = 4'd3;
@(posedge clk_i);
shared_exps0 = 8'd137;
shared_exps1 = 8'd124;
a_mant0 = 8'd202; a_mant1 = 8'd184; a_mant2 = 8'd189; a_mant3 = 8'd164;
b_mant0 = 8'd126; b_mant1 = 8'd60; b_mant2 = 8'd229; b_mant3 = 8'd170;
a_exp0 = 10'd636; a_exp1 = 10'd420; a_exp2 = 10'd117; a_exp3 = 10'd155;
b_exp0 = 10'd610; b_exp1 = 10'd96; b_exp2 = 10'd126; b_exp3 = 10'd436;
a_sign0 = 4'd12; a_sign1 = 4'd1; a_sign2 = 4'd10; a_sign3 = 4'd10;
b_sign0 = 4'd4; b_sign1 = 4'd0; b_sign2 = 4'd9; b_sign3 = 4'd5;
@(posedge clk_i);
a_mant0 = 8'd55; a_mant1 = 8'd199; a_mant2 = 8'd196; a_mant3 = 8'd1;
b_mant0 = 8'd242; b_mant1 = 8'd48; b_mant2 = 8'd229; b_mant3 = 8'd88;
a_exp0 = 10'd975; a_exp1 = 10'd1018; a_exp2 = 10'd366; a_exp3 = 10'd754;
b_exp0 = 10'd797; b_exp1 = 10'd21; b_exp2 = 10'd802; b_exp3 = 10'd431;
a_sign0 = 4'd2; a_sign1 = 4'd9; a_sign2 = 4'd1; a_sign3 = 4'd16;
b_sign0 = 4'd2; b_sign1 = 4'd16; b_sign2 = 4'd10; b_sign3 = 4'd1;
@(posedge clk_i);
a_mant0 = 8'd241; a_mant1 = 8'd98; a_mant2 = 8'd228; a_mant3 = 8'd26;
b_mant0 = 8'd32; b_mant1 = 8'd98; b_mant2 = 8'd187; b_mant3 = 8'd231;
a_exp0 = 10'd337; a_exp1 = 10'd254; a_exp2 = 10'd392; a_exp3 = 10'd360;
b_exp0 = 10'd376; b_exp1 = 10'd878; b_exp2 = 10'd164; b_exp3 = 10'd304;
a_sign0 = 4'd12; a_sign1 = 4'd3; a_sign2 = 4'd13; a_sign3 = 4'd14;
b_sign0 = 4'd16; b_sign1 = 4'd14; b_sign2 = 4'd0; b_sign3 = 4'd10;
@(posedge clk_i);
a_mant0 = 8'd174; a_mant1 = 8'd174; a_mant2 = 8'd143; a_mant3 = 8'd95;
b_mant0 = 8'd142; b_mant1 = 8'd19; b_mant2 = 8'd75; b_mant3 = 8'd29;
a_exp0 = 10'd14; a_exp1 = 10'd911; a_exp2 = 10'd373; a_exp3 = 10'd334;
b_exp0 = 10'd589; b_exp1 = 10'd556; b_exp2 = 10'd487; b_exp3 = 10'd1013;
a_sign0 = 4'd2; a_sign1 = 4'd15; a_sign2 = 4'd7; a_sign3 = 4'd11;
b_sign0 = 4'd7; b_sign1 = 4'd7; b_sign2 = 4'd12; b_sign3 = 4'd7;
@(posedge clk_i);
a_mant0 = 8'd86; a_mant1 = 8'd136; a_mant2 = 8'd26; a_mant3 = 8'd15;
b_mant0 = 8'd14; b_mant1 = 8'd106; b_mant2 = 8'd246; b_mant3 = 8'd5;
a_exp0 = 10'd243; a_exp1 = 10'd535; a_exp2 = 10'd705; a_exp3 = 10'd922;
b_exp0 = 10'd722; b_exp1 = 10'd4; b_exp2 = 10'd583; b_exp3 = 10'd518;
a_sign0 = 4'd1; a_sign1 = 4'd2; a_sign2 = 4'd3; a_sign3 = 4'd12;
b_sign0 = 4'd11; b_sign1 = 4'd14; b_sign2 = 4'd14; b_sign3 = 4'd5;
@(posedge clk_i);
a_mant0 = 8'd236; a_mant1 = 8'd249; a_mant2 = 8'd157; a_mant3 = 8'd249;
b_mant0 = 8'd164; b_mant1 = 8'd62; b_mant2 = 8'd29; b_mant3 = 8'd17;
a_exp0 = 10'd0; a_exp1 = 10'd806; a_exp2 = 10'd178; a_exp3 = 10'd94;
b_exp0 = 10'd154; b_exp1 = 10'd394; b_exp2 = 10'd13; b_exp3 = 10'd236;
a_sign0 = 4'd9; a_sign1 = 4'd9; a_sign2 = 4'd6; a_sign3 = 4'd11;
b_sign0 = 4'd6; b_sign1 = 4'd9; b_sign2 = 4'd12; b_sign3 = 4'd3;
@(posedge clk_i);
a_mant0 = 8'd12; a_mant1 = 8'd41; a_mant2 = 8'd185; a_mant3 = 8'd144;
b_mant0 = 8'd244; b_mant1 = 8'd250; b_mant2 = 8'd147; b_mant3 = 8'd199;
a_exp0 = 10'd683; a_exp1 = 10'd154; a_exp2 = 10'd665; a_exp3 = 10'd109;
b_exp0 = 10'd988; b_exp1 = 10'd182; b_exp2 = 10'd43; b_exp3 = 10'd664;
a_sign0 = 4'd5; a_sign1 = 4'd4; a_sign2 = 4'd3; a_sign3 = 4'd10;
b_sign0 = 4'd0; b_sign1 = 4'd6; b_sign2 = 4'd7; b_sign3 = 4'd13;
@(posedge clk_i);
a_mant0 = 8'd144; a_mant1 = 8'd59; a_mant2 = 8'd18; a_mant3 = 8'd222;
b_mant0 = 8'd216; b_mant1 = 8'd15; b_mant2 = 8'd148; b_mant3 = 8'd69;
a_exp0 = 10'd699; a_exp1 = 10'd730; a_exp2 = 10'd809; a_exp3 = 10'd965;
b_exp0 = 10'd534; b_exp1 = 10'd718; b_exp2 = 10'd783; b_exp3 = 10'd144;
a_sign0 = 4'd11; a_sign1 = 4'd0; a_sign2 = 4'd5; a_sign3 = 4'd10;
b_sign0 = 4'd11; b_sign1 = 4'd16; b_sign2 = 4'd8; b_sign3 = 4'd2;
@(posedge clk_i);
shared_exps0 = 8'd120;
shared_exps1 = 8'd125;
rstn = 0;
@(posedge clk_i);
rstn = 1;
a_mant0 = 8'd2; a_mant1 = 8'd143; a_mant2 = 8'd34; a_mant3 = 8'd199;
b_mant0 = 8'd28; b_mant1 = 8'd251; b_mant2 = 8'd123; b_mant3 = 8'd101;
a_exp0 = 10'd223; a_exp1 = 10'd39; a_exp2 = 10'd650; a_exp3 = 10'd602;
b_exp0 = 10'd460; b_exp1 = 10'd780; b_exp2 = 10'd935; b_exp3 = 10'd113;
a_sign0 = 4'd5; a_sign1 = 4'd13; a_sign2 = 4'd15; a_sign3 = 4'd10;
b_sign0 = 4'd16; b_sign1 = 4'd7; b_sign2 = 4'd7; b_sign3 = 4'd14;
@(posedge clk_i);
a_mant0 = 8'd243; a_mant1 = 8'd150; a_mant2 = 8'd53; a_mant3 = 8'd122;
b_mant0 = 8'd159; b_mant1 = 8'd72; b_mant2 = 8'd92; b_mant3 = 8'd117;
a_exp0 = 10'd2; a_exp1 = 10'd831; a_exp2 = 10'd266; a_exp3 = 10'd985;
b_exp0 = 10'd347; b_exp1 = 10'd619; b_exp2 = 10'd620; b_exp3 = 10'd271;
a_sign0 = 4'd12; a_sign1 = 4'd16; a_sign2 = 4'd8; a_sign3 = 4'd12;
b_sign0 = 4'd15; b_sign1 = 4'd9; b_sign2 = 4'd11; b_sign3 = 4'd9;
@(posedge clk_i);
a_mant0 = 8'd75; a_mant1 = 8'd120; a_mant2 = 8'd139; a_mant3 = 8'd233;
b_mant0 = 8'd14; b_mant1 = 8'd146; b_mant2 = 8'd182; b_mant3 = 8'd136;
a_exp0 = 10'd298; a_exp1 = 10'd760; a_exp2 = 10'd190; a_exp3 = 10'd386;
b_exp0 = 10'd928; b_exp1 = 10'd438; b_exp2 = 10'd801; b_exp3 = 10'd90;
a_sign0 = 4'd1; a_sign1 = 4'd11; a_sign2 = 4'd3; a_sign3 = 4'd1;
b_sign0 = 4'd6; b_sign1 = 4'd4; b_sign2 = 4'd10; b_sign3 = 4'd1;
@(posedge clk_i);
a_mant0 = 8'd81; a_mant1 = 8'd1; a_mant2 = 8'd66; a_mant3 = 8'd196;
b_mant0 = 8'd153; b_mant1 = 8'd148; b_mant2 = 8'd54; b_mant3 = 8'd109;
a_exp0 = 10'd960; a_exp1 = 10'd374; a_exp2 = 10'd238; a_exp3 = 10'd1004;
b_exp0 = 10'd332; b_exp1 = 10'd138; b_exp2 = 10'd751; b_exp3 = 10'd141;
a_sign0 = 4'd14; a_sign1 = 4'd11; a_sign2 = 4'd6; a_sign3 = 4'd8;
b_sign0 = 4'd0; b_sign1 = 4'd5; b_sign2 = 4'd6; b_sign3 = 4'd11;
@(posedge clk_i);
a_mant0 = 8'd25; a_mant1 = 8'd95; a_mant2 = 8'd101; a_mant3 = 8'd100;
b_mant0 = 8'd132; b_mant1 = 8'd109; b_mant2 = 8'd134; b_mant3 = 8'd193;
a_exp0 = 10'd179; a_exp1 = 10'd293; a_exp2 = 10'd204; a_exp3 = 10'd340;
b_exp0 = 10'd868; b_exp1 = 10'd8; b_exp2 = 10'd102; b_exp3 = 10'd731;
a_sign0 = 4'd9; a_sign1 = 4'd10; a_sign2 = 4'd9; a_sign3 = 4'd10;
b_sign0 = 4'd12; b_sign1 = 4'd12; b_sign2 = 4'd6; b_sign3 = 4'd3;
@(posedge clk_i);
a_mant0 = 8'd80; a_mant1 = 8'd158; a_mant2 = 8'd193; a_mant3 = 8'd65;
b_mant0 = 8'd150; b_mant1 = 8'd32; b_mant2 = 8'd44; b_mant3 = 8'd148;
a_exp0 = 10'd892; a_exp1 = 10'd276; a_exp2 = 10'd222; a_exp3 = 10'd606;
b_exp0 = 10'd754; b_exp1 = 10'd481; b_exp2 = 10'd713; b_exp3 = 10'd527;
a_sign0 = 4'd12; a_sign1 = 4'd3; a_sign2 = 4'd14; a_sign3 = 4'd3;
b_sign0 = 4'd15; b_sign1 = 4'd16; b_sign2 = 4'd1; b_sign3 = 4'd2;
@(posedge clk_i);
a_mant0 = 8'd58; a_mant1 = 8'd89; a_mant2 = 8'd136; a_mant3 = 8'd73;
b_mant0 = 8'd212; b_mant1 = 8'd192; b_mant2 = 8'd139; b_mant3 = 8'd246;
a_exp0 = 10'd670; a_exp1 = 10'd745; a_exp2 = 10'd427; a_exp3 = 10'd7;
b_exp0 = 10'd576; b_exp1 = 10'd64; b_exp2 = 10'd367; b_exp3 = 10'd305;
a_sign0 = 4'd11; a_sign1 = 4'd14; a_sign2 = 4'd4; a_sign3 = 4'd1;
b_sign0 = 4'd6; b_sign1 = 4'd1; b_sign2 = 4'd10; b_sign3 = 4'd0;
@(posedge clk_i);
shared_exps0 = 8'd133;
shared_exps1 = 8'd123;
a_mant0 = 8'd115; a_mant1 = 8'd63; a_mant2 = 8'd1; a_mant3 = 8'd58;
b_mant0 = 8'd169; b_mant1 = 8'd100; b_mant2 = 8'd173; b_mant3 = 8'd162;
a_exp0 = 10'd783; a_exp1 = 10'd888; a_exp2 = 10'd492; a_exp3 = 10'd947;
b_exp0 = 10'd757; b_exp1 = 10'd436; b_exp2 = 10'd268; b_exp3 = 10'd723;
a_sign0 = 4'd3; a_sign1 = 4'd12; a_sign2 = 4'd15; a_sign3 = 4'd15;
b_sign0 = 4'd8; b_sign1 = 4'd16; b_sign2 = 4'd8; b_sign3 = 4'd8;
@(posedge clk_i);
a_mant0 = 8'd142; a_mant1 = 8'd17; a_mant2 = 8'd35; a_mant3 = 8'd18;
b_mant0 = 8'd182; b_mant1 = 8'd49; b_mant2 = 8'd103; b_mant3 = 8'd226;
a_exp0 = 10'd43; a_exp1 = 10'd430; a_exp2 = 10'd646; a_exp3 = 10'd99;
b_exp0 = 10'd972; b_exp1 = 10'd616; b_exp2 = 10'd302; b_exp3 = 10'd712;
a_sign0 = 4'd11; a_sign1 = 4'd15; a_sign2 = 4'd5; a_sign3 = 4'd16;
b_sign0 = 4'd15; b_sign1 = 4'd6; b_sign2 = 4'd5; b_sign3 = 4'd7;
@(posedge clk_i);
a_mant0 = 8'd151; a_mant1 = 8'd133; a_mant2 = 8'd40; a_mant3 = 8'd255;
b_mant0 = 8'd33; b_mant1 = 8'd12; b_mant2 = 8'd177; b_mant3 = 8'd213;
a_exp0 = 10'd11; a_exp1 = 10'd121; a_exp2 = 10'd609; a_exp3 = 10'd168;
b_exp0 = 10'd788; b_exp1 = 10'd205; b_exp2 = 10'd1004; b_exp3 = 10'd293;
a_sign0 = 4'd0; a_sign1 = 4'd13; a_sign2 = 4'd10; a_sign3 = 4'd7;
b_sign0 = 4'd9; b_sign1 = 4'd4; b_sign2 = 4'd3; b_sign3 = 4'd9;
@(posedge clk_i);
a_mant0 = 8'd245; a_mant1 = 8'd219; a_mant2 = 8'd221; a_mant3 = 8'd106;
b_mant0 = 8'd231; b_mant1 = 8'd96; b_mant2 = 8'd102; b_mant3 = 8'd82;
a_exp0 = 10'd277; a_exp1 = 10'd280; a_exp2 = 10'd525; a_exp3 = 10'd32;
b_exp0 = 10'd807; b_exp1 = 10'd339; b_exp2 = 10'd553; b_exp3 = 10'd190;
a_sign0 = 4'd15; a_sign1 = 4'd3; a_sign2 = 4'd13; a_sign3 = 4'd10;
b_sign0 = 4'd16; b_sign1 = 4'd4; b_sign2 = 4'd6; b_sign3 = 4'd11;
@(posedge clk_i);
a_mant0 = 8'd110; a_mant1 = 8'd47; a_mant2 = 8'd46; a_mant3 = 8'd245;
b_mant0 = 8'd173; b_mant1 = 8'd190; b_mant2 = 8'd100; b_mant3 = 8'd195;
a_exp0 = 10'd908; a_exp1 = 10'd743; a_exp2 = 10'd388; a_exp3 = 10'd534;
b_exp0 = 10'd741; b_exp1 = 10'd290; b_exp2 = 10'd884; b_exp3 = 10'd754;
a_sign0 = 4'd14; a_sign1 = 4'd5; a_sign2 = 4'd11; a_sign3 = 4'd8;
b_sign0 = 4'd4; b_sign1 = 4'd10; b_sign2 = 4'd1; b_sign3 = 4'd14;
@(posedge clk_i);
a_mant0 = 8'd133; a_mant1 = 8'd120; a_mant2 = 8'd153; a_mant3 = 8'd112;
b_mant0 = 8'd20; b_mant1 = 8'd211; b_mant2 = 8'd198; b_mant3 = 8'd130;
a_exp0 = 10'd75; a_exp1 = 10'd853; a_exp2 = 10'd640; a_exp3 = 10'd759;
b_exp0 = 10'd393; b_exp1 = 10'd666; b_exp2 = 10'd774; b_exp3 = 10'd498;
a_sign0 = 4'd3; a_sign1 = 4'd7; a_sign2 = 4'd8; a_sign3 = 4'd15;
b_sign0 = 4'd4; b_sign1 = 4'd7; b_sign2 = 4'd6; b_sign3 = 4'd14;
@(posedge clk_i);
a_mant0 = 8'd220; a_mant1 = 8'd173; a_mant2 = 8'd42; a_mant3 = 8'd246;
b_mant0 = 8'd140; b_mant1 = 8'd51; b_mant2 = 8'd199; b_mant3 = 8'd211;
a_exp0 = 10'd732; a_exp1 = 10'd467; a_exp2 = 10'd250; a_exp3 = 10'd76;
b_exp0 = 10'd510; b_exp1 = 10'd227; b_exp2 = 10'd561; b_exp3 = 10'd203;
a_sign0 = 4'd12; a_sign1 = 4'd15; a_sign2 = 4'd4; a_sign3 = 4'd5;
b_sign0 = 4'd15; b_sign1 = 4'd4; b_sign2 = 4'd16; b_sign3 = 4'd16;
@(posedge clk_i);
a_mant0 = 8'd27; a_mant1 = 8'd144; a_mant2 = 8'd116; a_mant3 = 8'd10;
b_mant0 = 8'd253; b_mant1 = 8'd206; b_mant2 = 8'd206; b_mant3 = 8'd23;
a_exp0 = 10'd910; a_exp1 = 10'd590; a_exp2 = 10'd172; a_exp3 = 10'd15;
b_exp0 = 10'd847; b_exp1 = 10'd921; b_exp2 = 10'd885; b_exp3 = 10'd150;
a_sign0 = 4'd0; a_sign1 = 4'd3; a_sign2 = 4'd15; a_sign3 = 4'd4;
b_sign0 = 4'd15; b_sign1 = 4'd12; b_sign2 = 4'd7; b_sign3 = 4'd12;
@(posedge clk_i);
shared_exps0 = 8'd147;
shared_exps1 = 8'd117;
a_mant0 = 8'd81; a_mant1 = 8'd32; a_mant2 = 8'd81; a_mant3 = 8'd0;
b_mant0 = 8'd200; b_mant1 = 8'd42; b_mant2 = 8'd39; b_mant3 = 8'd86;
a_exp0 = 10'd775; a_exp1 = 10'd338; a_exp2 = 10'd343; a_exp3 = 10'd760;
b_exp0 = 10'd392; b_exp1 = 10'd622; b_exp2 = 10'd608; b_exp3 = 10'd59;
a_sign0 = 4'd0; a_sign1 = 4'd15; a_sign2 = 4'd0; a_sign3 = 4'd1;
b_sign0 = 4'd13; b_sign1 = 4'd5; b_sign2 = 4'd0; b_sign3 = 4'd14;
@(posedge clk_i);
a_mant0 = 8'd154; a_mant1 = 8'd57; a_mant2 = 8'd149; a_mant3 = 8'd170;
b_mant0 = 8'd233; b_mant1 = 8'd109; b_mant2 = 8'd104; b_mant3 = 8'd2;
a_exp0 = 10'd629; a_exp1 = 10'd989; a_exp2 = 10'd200; a_exp3 = 10'd372;
b_exp0 = 10'd724; b_exp1 = 10'd502; b_exp2 = 10'd76; b_exp3 = 10'd56;
a_sign0 = 4'd0; a_sign1 = 4'd15; a_sign2 = 4'd8; a_sign3 = 4'd13;
b_sign0 = 4'd10; b_sign1 = 4'd16; b_sign2 = 4'd13; b_sign3 = 4'd6;
@(posedge clk_i);
a_mant0 = 8'd26; a_mant1 = 8'd131; a_mant2 = 8'd236; a_mant3 = 8'd223;
b_mant0 = 8'd51; b_mant1 = 8'd40; b_mant2 = 8'd147; b_mant3 = 8'd58;
a_exp0 = 10'd359; a_exp1 = 10'd961; a_exp2 = 10'd632; a_exp3 = 10'd654;
b_exp0 = 10'd240; b_exp1 = 10'd862; b_exp2 = 10'd440; b_exp3 = 10'd736;
a_sign0 = 4'd3; a_sign1 = 4'd11; a_sign2 = 4'd6; a_sign3 = 4'd14;
b_sign0 = 4'd1; b_sign1 = 4'd13; b_sign2 = 4'd8; b_sign3 = 4'd4;
@(posedge clk_i);
a_mant0 = 8'd216; a_mant1 = 8'd213; a_mant2 = 8'd138; a_mant3 = 8'd171;
b_mant0 = 8'd2; b_mant1 = 8'd149; b_mant2 = 8'd248; b_mant3 = 8'd159;
a_exp0 = 10'd143; a_exp1 = 10'd291; a_exp2 = 10'd958; a_exp3 = 10'd647;
b_exp0 = 10'd328; b_exp1 = 10'd575; b_exp2 = 10'd11; b_exp3 = 10'd509;
a_sign0 = 4'd10; a_sign1 = 4'd11; a_sign2 = 4'd11; a_sign3 = 4'd2;
b_sign0 = 4'd16; b_sign1 = 4'd12; b_sign2 = 4'd9; b_sign3 = 4'd7;
@(posedge clk_i);
a_mant0 = 8'd196; a_mant1 = 8'd25; a_mant2 = 8'd23; a_mant3 = 8'd63;
b_mant0 = 8'd216; b_mant1 = 8'd108; b_mant2 = 8'd56; b_mant3 = 8'd180;
a_exp0 = 10'd836; a_exp1 = 10'd876; a_exp2 = 10'd747; a_exp3 = 10'd149;
b_exp0 = 10'd272; b_exp1 = 10'd597; b_exp2 = 10'd450; b_exp3 = 10'd834;
a_sign0 = 4'd0; a_sign1 = 4'd12; a_sign2 = 4'd16; a_sign3 = 4'd14;
b_sign0 = 4'd7; b_sign1 = 4'd7; b_sign2 = 4'd4; b_sign3 = 4'd6;
@(posedge clk_i);
a_mant0 = 8'd73; a_mant1 = 8'd153; a_mant2 = 8'd136; a_mant3 = 8'd195;
b_mant0 = 8'd238; b_mant1 = 8'd98; b_mant2 = 8'd90; b_mant3 = 8'd241;
a_exp0 = 10'd512; a_exp1 = 10'd386; a_exp2 = 10'd925; a_exp3 = 10'd534;
b_exp0 = 10'd876; b_exp1 = 10'd203; b_exp2 = 10'd180; b_exp3 = 10'd989;
a_sign0 = 4'd14; a_sign1 = 4'd14; a_sign2 = 4'd3; a_sign3 = 4'd1;
b_sign0 = 4'd6; b_sign1 = 4'd12; b_sign2 = 4'd9; b_sign3 = 4'd3;
@(posedge clk_i);
a_mant0 = 8'd187; a_mant1 = 8'd169; a_mant2 = 8'd184; a_mant3 = 8'd193;
b_mant0 = 8'd176; b_mant1 = 8'd11; b_mant2 = 8'd67; b_mant3 = 8'd182;
a_exp0 = 10'd495; a_exp1 = 10'd309; a_exp2 = 10'd708; a_exp3 = 10'd773;
b_exp0 = 10'd636; b_exp1 = 10'd42; b_exp2 = 10'd51; b_exp3 = 10'd230;
a_sign0 = 4'd14; a_sign1 = 4'd9; a_sign2 = 4'd14; a_sign3 = 4'd10;
b_sign0 = 4'd2; b_sign1 = 4'd3; b_sign2 = 4'd4; b_sign3 = 4'd16;
@(posedge clk_i);
a_mant0 = 8'd241; a_mant1 = 8'd130; a_mant2 = 8'd170; a_mant3 = 8'd244;
b_mant0 = 8'd208; b_mant1 = 8'd100; b_mant2 = 8'd204; b_mant3 = 8'd233;
a_exp0 = 10'd658; a_exp1 = 10'd908; a_exp2 = 10'd386; a_exp3 = 10'd851;
b_exp0 = 10'd795; b_exp1 = 10'd189; b_exp2 = 10'd897; b_exp3 = 10'd927;
a_sign0 = 4'd4; a_sign1 = 4'd16; a_sign2 = 4'd3; a_sign3 = 4'd6;
b_sign0 = 4'd5; b_sign1 = 4'd6; b_sign2 = 4'd10; b_sign3 = 4'd8;
@(posedge clk_i);
shared_exps0 = 8'd114;
shared_exps1 = 8'd118;
a_mant0 = 8'd15; a_mant1 = 8'd165; a_mant2 = 8'd210; a_mant3 = 8'd59;
b_mant0 = 8'd59; b_mant1 = 8'd111; b_mant2 = 8'd76; b_mant3 = 8'd183;
a_exp0 = 10'd886; a_exp1 = 10'd628; a_exp2 = 10'd848; a_exp3 = 10'd605;
b_exp0 = 10'd800; b_exp1 = 10'd1020; b_exp2 = 10'd729; b_exp3 = 10'd322;
a_sign0 = 4'd4; a_sign1 = 4'd7; a_sign2 = 4'd6; a_sign3 = 4'd13;
b_sign0 = 4'd2; b_sign1 = 4'd12; b_sign2 = 4'd0; b_sign3 = 4'd16;
@(posedge clk_i);
a_mant0 = 8'd210; a_mant1 = 8'd89; a_mant2 = 8'd249; a_mant3 = 8'd12;
b_mant0 = 8'd197; b_mant1 = 8'd61; b_mant2 = 8'd69; b_mant3 = 8'd109;
a_exp0 = 10'd279; a_exp1 = 10'd431; a_exp2 = 10'd918; a_exp3 = 10'd910;
b_exp0 = 10'd461; b_exp1 = 10'd178; b_exp2 = 10'd761; b_exp3 = 10'd945;
a_sign0 = 4'd2; a_sign1 = 4'd4; a_sign2 = 4'd10; a_sign3 = 4'd2;
b_sign0 = 4'd6; b_sign1 = 4'd5; b_sign2 = 4'd4; b_sign3 = 4'd8;
@(posedge clk_i);
a_mant0 = 8'd50; a_mant1 = 8'd165; a_mant2 = 8'd221; a_mant3 = 8'd157;
b_mant0 = 8'd76; b_mant1 = 8'd238; b_mant2 = 8'd170; b_mant3 = 8'd215;
a_exp0 = 10'd569; a_exp1 = 10'd523; a_exp2 = 10'd769; a_exp3 = 10'd18;
b_exp0 = 10'd380; b_exp1 = 10'd356; b_exp2 = 10'd187; b_exp3 = 10'd1;
a_sign0 = 4'd5; a_sign1 = 4'd14; a_sign2 = 4'd10; a_sign3 = 4'd5;
b_sign0 = 4'd7; b_sign1 = 4'd13; b_sign2 = 4'd15; b_sign3 = 4'd4;
@(posedge clk_i);
a_mant0 = 8'd22; a_mant1 = 8'd92; a_mant2 = 8'd156; a_mant3 = 8'd180;
b_mant0 = 8'd42; b_mant1 = 8'd235; b_mant2 = 8'd179; b_mant3 = 8'd179;
a_exp0 = 10'd387; a_exp1 = 10'd449; a_exp2 = 10'd748; a_exp3 = 10'd141;
b_exp0 = 10'd830; b_exp1 = 10'd437; b_exp2 = 10'd142; b_exp3 = 10'd440;
a_sign0 = 4'd8; a_sign1 = 4'd4; a_sign2 = 4'd10; a_sign3 = 4'd8;
b_sign0 = 4'd10; b_sign1 = 4'd16; b_sign2 = 4'd16; b_sign3 = 4'd6;
@(posedge clk_i);
a_mant0 = 8'd88; a_mant1 = 8'd24; a_mant2 = 8'd67; a_mant3 = 8'd253;
b_mant0 = 8'd186; b_mant1 = 8'd129; b_mant2 = 8'd201; b_mant3 = 8'd183;
a_exp0 = 10'd113; a_exp1 = 10'd81; a_exp2 = 10'd479; a_exp3 = 10'd428;
b_exp0 = 10'd497; b_exp1 = 10'd402; b_exp2 = 10'd694; b_exp3 = 10'd776;
a_sign0 = 4'd16; a_sign1 = 4'd15; a_sign2 = 4'd1; a_sign3 = 4'd6;
b_sign0 = 4'd1; b_sign1 = 4'd2; b_sign2 = 4'd8; b_sign3 = 4'd2;
@(posedge clk_i);
a_mant0 = 8'd46; a_mant1 = 8'd148; a_mant2 = 8'd70; a_mant3 = 8'd151;
b_mant0 = 8'd174; b_mant1 = 8'd241; b_mant2 = 8'd171; b_mant3 = 8'd163;
a_exp0 = 10'd679; a_exp1 = 10'd699; a_exp2 = 10'd8; a_exp3 = 10'd562;
b_exp0 = 10'd912; b_exp1 = 10'd167; b_exp2 = 10'd435; b_exp3 = 10'd1019;
a_sign0 = 4'd6; a_sign1 = 4'd16; a_sign2 = 4'd2; a_sign3 = 4'd6;
b_sign0 = 4'd11; b_sign1 = 4'd15; b_sign2 = 4'd6; b_sign3 = 4'd9;
@(posedge clk_i);
a_mant0 = 8'd251; a_mant1 = 8'd106; a_mant2 = 8'd251; a_mant3 = 8'd92;
b_mant0 = 8'd211; b_mant1 = 8'd182; b_mant2 = 8'd160; b_mant3 = 8'd89;
a_exp0 = 10'd155; a_exp1 = 10'd947; a_exp2 = 10'd309; a_exp3 = 10'd370;
b_exp0 = 10'd774; b_exp1 = 10'd269; b_exp2 = 10'd562; b_exp3 = 10'd1018;
a_sign0 = 4'd11; a_sign1 = 4'd13; a_sign2 = 4'd4; a_sign3 = 4'd0;
b_sign0 = 4'd8; b_sign1 = 4'd6; b_sign2 = 4'd7; b_sign3 = 4'd11;
@(posedge clk_i);
a_mant0 = 8'd87; a_mant1 = 8'd239; a_mant2 = 8'd106; a_mant3 = 8'd222;
b_mant0 = 8'd76; b_mant1 = 8'd85; b_mant2 = 8'd255; b_mant3 = 8'd236;
a_exp0 = 10'd154; a_exp1 = 10'd898; a_exp2 = 10'd530; a_exp3 = 10'd556;
b_exp0 = 10'd123; b_exp1 = 10'd626; b_exp2 = 10'd570; b_exp3 = 10'd530;
a_sign0 = 4'd0; a_sign1 = 4'd14; a_sign2 = 4'd3; a_sign3 = 4'd13;
b_sign0 = 4'd6; b_sign1 = 4'd5; b_sign2 = 4'd16; b_sign3 = 4'd14;
@(posedge clk_i);
shared_exps0 = 8'd133;
shared_exps1 = 8'd167;
rstn = 0;
@(posedge clk_i);
rstn = 1;
a_mant0 = 8'd170; a_mant1 = 8'd230; a_mant2 = 8'd118; a_mant3 = 8'd182;
b_mant0 = 8'd218; b_mant1 = 8'd103; b_mant2 = 8'd233; b_mant3 = 8'd106;
a_exp0 = 10'd311; a_exp1 = 10'd759; a_exp2 = 10'd140; a_exp3 = 10'd446;
b_exp0 = 10'd834; b_exp1 = 10'd7; b_exp2 = 10'd957; b_exp3 = 10'd78;
a_sign0 = 4'd1; a_sign1 = 4'd1; a_sign2 = 4'd11; a_sign3 = 4'd12;
b_sign0 = 4'd8; b_sign1 = 4'd10; b_sign2 = 4'd4; b_sign3 = 4'd7;
@(posedge clk_i);
a_mant0 = 8'd183; a_mant1 = 8'd213; a_mant2 = 8'd20; a_mant3 = 8'd15;
b_mant0 = 8'd25; b_mant1 = 8'd222; b_mant2 = 8'd54; b_mant3 = 8'd62;
a_exp0 = 10'd8; a_exp1 = 10'd115; a_exp2 = 10'd723; a_exp3 = 10'd188;
b_exp0 = 10'd653; b_exp1 = 10'd782; b_exp2 = 10'd36; b_exp3 = 10'd590;
a_sign0 = 4'd1; a_sign1 = 4'd13; a_sign2 = 4'd5; a_sign3 = 4'd16;
b_sign0 = 4'd10; b_sign1 = 4'd7; b_sign2 = 4'd16; b_sign3 = 4'd6;
@(posedge clk_i);
a_mant0 = 8'd146; a_mant1 = 8'd135; a_mant2 = 8'd170; a_mant3 = 8'd146;
b_mant0 = 8'd23; b_mant1 = 8'd128; b_mant2 = 8'd165; b_mant3 = 8'd136;
a_exp0 = 10'd29; a_exp1 = 10'd594; a_exp2 = 10'd440; a_exp3 = 10'd582;
b_exp0 = 10'd211; b_exp1 = 10'd614; b_exp2 = 10'd129; b_exp3 = 10'd64;
a_sign0 = 4'd12; a_sign1 = 4'd9; a_sign2 = 4'd2; a_sign3 = 4'd16;
b_sign0 = 4'd12; b_sign1 = 4'd16; b_sign2 = 4'd16; b_sign3 = 4'd3;
@(posedge clk_i);
a_mant0 = 8'd222; a_mant1 = 8'd158; a_mant2 = 8'd15; a_mant3 = 8'd229;
b_mant0 = 8'd161; b_mant1 = 8'd39; b_mant2 = 8'd183; b_mant3 = 8'd8;
a_exp0 = 10'd1006; a_exp1 = 10'd685; a_exp2 = 10'd675; a_exp3 = 10'd537;
b_exp0 = 10'd757; b_exp1 = 10'd549; b_exp2 = 10'd252; b_exp3 = 10'd1000;
a_sign0 = 4'd13; a_sign1 = 4'd7; a_sign2 = 4'd4; a_sign3 = 4'd14;
b_sign0 = 4'd5; b_sign1 = 4'd2; b_sign2 = 4'd10; b_sign3 = 4'd14;
@(posedge clk_i);
a_mant0 = 8'd223; a_mant1 = 8'd12; a_mant2 = 8'd144; a_mant3 = 8'd117;
b_mant0 = 8'd145; b_mant1 = 8'd131; b_mant2 = 8'd174; b_mant3 = 8'd168;
a_exp0 = 10'd899; a_exp1 = 10'd1007; a_exp2 = 10'd89; a_exp3 = 10'd770;
b_exp0 = 10'd536; b_exp1 = 10'd1010; b_exp2 = 10'd196; b_exp3 = 10'd132;
a_sign0 = 4'd9; a_sign1 = 4'd6; a_sign2 = 4'd1; a_sign3 = 4'd6;
b_sign0 = 4'd2; b_sign1 = 4'd6; b_sign2 = 4'd6; b_sign3 = 4'd16;
@(posedge clk_i);
a_mant0 = 8'd15; a_mant1 = 8'd234; a_mant2 = 8'd99; a_mant3 = 8'd27;
b_mant0 = 8'd234; b_mant1 = 8'd48; b_mant2 = 8'd106; b_mant3 = 8'd82;
a_exp0 = 10'd475; a_exp1 = 10'd465; a_exp2 = 10'd773; a_exp3 = 10'd705;
b_exp0 = 10'd402; b_exp1 = 10'd265; b_exp2 = 10'd839; b_exp3 = 10'd895;
a_sign0 = 4'd9; a_sign1 = 4'd9; a_sign2 = 4'd7; a_sign3 = 4'd10;
b_sign0 = 4'd15; b_sign1 = 4'd14; b_sign2 = 4'd15; b_sign3 = 4'd15;
@(posedge clk_i);
a_mant0 = 8'd116; a_mant1 = 8'd207; a_mant2 = 8'd125; a_mant3 = 8'd138;
b_mant0 = 8'd226; b_mant1 = 8'd141; b_mant2 = 8'd173; b_mant3 = 8'd255;
a_exp0 = 10'd909; a_exp1 = 10'd903; a_exp2 = 10'd473; a_exp3 = 10'd520;
b_exp0 = 10'd99; b_exp1 = 10'd52; b_exp2 = 10'd345; b_exp3 = 10'd639;
a_sign0 = 4'd14; a_sign1 = 4'd12; a_sign2 = 4'd3; a_sign3 = 4'd9;
b_sign0 = 4'd1; b_sign1 = 4'd3; b_sign2 = 4'd3; b_sign3 = 4'd15;
@(posedge clk_i);
shared_exps0 = 8'd136;
shared_exps1 = 8'd126;
a_mant0 = 8'd199; a_mant1 = 8'd40; a_mant2 = 8'd39; a_mant3 = 8'd228;
b_mant0 = 8'd134; b_mant1 = 8'd75; b_mant2 = 8'd11; b_mant3 = 8'd253;
a_exp0 = 10'd383; a_exp1 = 10'd290; a_exp2 = 10'd35; a_exp3 = 10'd488;
b_exp0 = 10'd1010; b_exp1 = 10'd437; b_exp2 = 10'd38; b_exp3 = 10'd721;
a_sign0 = 4'd8; a_sign1 = 4'd1; a_sign2 = 4'd3; a_sign3 = 4'd2;
b_sign0 = 4'd9; b_sign1 = 4'd3; b_sign2 = 4'd2; b_sign3 = 4'd16;
@(posedge clk_i);
a_mant0 = 8'd117; a_mant1 = 8'd93; a_mant2 = 8'd179; a_mant3 = 8'd181;
b_mant0 = 8'd21; b_mant1 = 8'd40; b_mant2 = 8'd70; b_mant3 = 8'd71;
a_exp0 = 10'd197; a_exp1 = 10'd21; a_exp2 = 10'd899; a_exp3 = 10'd491;
b_exp0 = 10'd159; b_exp1 = 10'd969; b_exp2 = 10'd368; b_exp3 = 10'd458;
a_sign0 = 4'd14; a_sign1 = 4'd14; a_sign2 = 4'd6; a_sign3 = 4'd9;
b_sign0 = 4'd7; b_sign1 = 4'd11; b_sign2 = 4'd11; b_sign3 = 4'd12;
@(posedge clk_i);
a_mant0 = 8'd87; a_mant1 = 8'd54; a_mant2 = 8'd197; a_mant3 = 8'd221;
b_mant0 = 8'd57; b_mant1 = 8'd127; b_mant2 = 8'd73; b_mant3 = 8'd191;
a_exp0 = 10'd742; a_exp1 = 10'd47; a_exp2 = 10'd199; a_exp3 = 10'd603;
b_exp0 = 10'd896; b_exp1 = 10'd935; b_exp2 = 10'd516; b_exp3 = 10'd442;
a_sign0 = 4'd9; a_sign1 = 4'd12; a_sign2 = 4'd3; a_sign3 = 4'd5;
b_sign0 = 4'd8; b_sign1 = 4'd3; b_sign2 = 4'd3; b_sign3 = 4'd5;
@(posedge clk_i);
a_mant0 = 8'd54; a_mant1 = 8'd143; a_mant2 = 8'd96; a_mant3 = 8'd67;
b_mant0 = 8'd164; b_mant1 = 8'd64; b_mant2 = 8'd197; b_mant3 = 8'd19;
a_exp0 = 10'd780; a_exp1 = 10'd251; a_exp2 = 10'd692; a_exp3 = 10'd872;
b_exp0 = 10'd203; b_exp1 = 10'd470; b_exp2 = 10'd527; b_exp3 = 10'd673;
a_sign0 = 4'd3; a_sign1 = 4'd14; a_sign2 = 4'd8; a_sign3 = 4'd3;
b_sign0 = 4'd3; b_sign1 = 4'd6; b_sign2 = 4'd4; b_sign3 = 4'd5;
@(posedge clk_i);
a_mant0 = 8'd111; a_mant1 = 8'd228; a_mant2 = 8'd165; a_mant3 = 8'd229;
b_mant0 = 8'd9; b_mant1 = 8'd243; b_mant2 = 8'd41; b_mant3 = 8'd228;
a_exp0 = 10'd203; a_exp1 = 10'd210; a_exp2 = 10'd128; a_exp3 = 10'd354;
b_exp0 = 10'd268; b_exp1 = 10'd1001; b_exp2 = 10'd843; b_exp3 = 10'd50;
a_sign0 = 4'd11; a_sign1 = 4'd13; a_sign2 = 4'd10; a_sign3 = 4'd12;
b_sign0 = 4'd11; b_sign1 = 4'd11; b_sign2 = 4'd13; b_sign3 = 4'd8;
@(posedge clk_i);
a_mant0 = 8'd64; a_mant1 = 8'd180; a_mant2 = 8'd121; a_mant3 = 8'd137;
b_mant0 = 8'd81; b_mant1 = 8'd117; b_mant2 = 8'd203; b_mant3 = 8'd178;
a_exp0 = 10'd86; a_exp1 = 10'd47; a_exp2 = 10'd671; a_exp3 = 10'd542;
b_exp0 = 10'd1018; b_exp1 = 10'd546; b_exp2 = 10'd8; b_exp3 = 10'd1003;
a_sign0 = 4'd11; a_sign1 = 4'd8; a_sign2 = 4'd11; a_sign3 = 4'd5;
b_sign0 = 4'd10; b_sign1 = 4'd4; b_sign2 = 4'd13; b_sign3 = 4'd16;
@(posedge clk_i);
a_mant0 = 8'd202; a_mant1 = 8'd0; a_mant2 = 8'd230; a_mant3 = 8'd144;
b_mant0 = 8'd246; b_mant1 = 8'd185; b_mant2 = 8'd249; b_mant3 = 8'd203;
a_exp0 = 10'd78; a_exp1 = 10'd384; a_exp2 = 10'd746; a_exp3 = 10'd920;
b_exp0 = 10'd527; b_exp1 = 10'd583; b_exp2 = 10'd273; b_exp3 = 10'd798;
a_sign0 = 4'd11; a_sign1 = 4'd14; a_sign2 = 4'd2; a_sign3 = 4'd10;
b_sign0 = 4'd15; b_sign1 = 4'd15; b_sign2 = 4'd11; b_sign3 = 4'd4;
@(posedge clk_i);
a_mant0 = 8'd153; a_mant1 = 8'd199; a_mant2 = 8'd65; a_mant3 = 8'd92;
b_mant0 = 8'd134; b_mant1 = 8'd64; b_mant2 = 8'd9; b_mant3 = 8'd98;
a_exp0 = 10'd620; a_exp1 = 10'd403; a_exp2 = 10'd157; a_exp3 = 10'd637;
b_exp0 = 10'd95; b_exp1 = 10'd323; b_exp2 = 10'd742; b_exp3 = 10'd931;
a_sign0 = 4'd3; a_sign1 = 4'd12; a_sign2 = 4'd6; a_sign3 = 4'd8;
b_sign0 = 4'd4; b_sign1 = 4'd11; b_sign2 = 4'd2; b_sign3 = 4'd7;
@(posedge clk_i);
shared_exps0 = 8'd130;
shared_exps1 = 8'd117;
a_mant0 = 8'd216; a_mant1 = 8'd69; a_mant2 = 8'd94; a_mant3 = 8'd70;
b_mant0 = 8'd110; b_mant1 = 8'd48; b_mant2 = 8'd109; b_mant3 = 8'd159;
a_exp0 = 10'd637; a_exp1 = 10'd574; a_exp2 = 10'd61; a_exp3 = 10'd699;
b_exp0 = 10'd735; b_exp1 = 10'd194; b_exp2 = 10'd693; b_exp3 = 10'd239;
a_sign0 = 4'd0; a_sign1 = 4'd16; a_sign2 = 4'd2; a_sign3 = 4'd4;
b_sign0 = 4'd12; b_sign1 = 4'd11; b_sign2 = 4'd9; b_sign3 = 4'd10;
@(posedge clk_i);
a_mant0 = 8'd168; a_mant1 = 8'd19; a_mant2 = 8'd110; a_mant3 = 8'd44;
b_mant0 = 8'd47; b_mant1 = 8'd156; b_mant2 = 8'd85; b_mant3 = 8'd246;
a_exp0 = 10'd732; a_exp1 = 10'd70; a_exp2 = 10'd7; a_exp3 = 10'd715;
b_exp0 = 10'd116; b_exp1 = 10'd990; b_exp2 = 10'd629; b_exp3 = 10'd123;
a_sign0 = 4'd9; a_sign1 = 4'd0; a_sign2 = 4'd15; a_sign3 = 4'd9;
b_sign0 = 4'd7; b_sign1 = 4'd4; b_sign2 = 4'd15; b_sign3 = 4'd4;
@(posedge clk_i);
a_mant0 = 8'd37; a_mant1 = 8'd28; a_mant2 = 8'd152; a_mant3 = 8'd32;
b_mant0 = 8'd158; b_mant1 = 8'd186; b_mant2 = 8'd109; b_mant3 = 8'd175;
a_exp0 = 10'd157; a_exp1 = 10'd628; a_exp2 = 10'd241; a_exp3 = 10'd407;
b_exp0 = 10'd802; b_exp1 = 10'd480; b_exp2 = 10'd1017; b_exp3 = 10'd492;
a_sign0 = 4'd0; a_sign1 = 4'd13; a_sign2 = 4'd16; a_sign3 = 4'd3;
b_sign0 = 4'd9; b_sign1 = 4'd5; b_sign2 = 4'd12; b_sign3 = 4'd7;
@(posedge clk_i);
a_mant0 = 8'd40; a_mant1 = 8'd155; a_mant2 = 8'd13; a_mant3 = 8'd21;
b_mant0 = 8'd240; b_mant1 = 8'd101; b_mant2 = 8'd148; b_mant3 = 8'd125;
a_exp0 = 10'd648; a_exp1 = 10'd939; a_exp2 = 10'd884; a_exp3 = 10'd533;
b_exp0 = 10'd718; b_exp1 = 10'd350; b_exp2 = 10'd801; b_exp3 = 10'd859;
a_sign0 = 4'd5; a_sign1 = 4'd11; a_sign2 = 4'd7; a_sign3 = 4'd2;
b_sign0 = 4'd13; b_sign1 = 4'd14; b_sign2 = 4'd4; b_sign3 = 4'd10;
@(posedge clk_i);
a_mant0 = 8'd213; a_mant1 = 8'd31; a_mant2 = 8'd154; a_mant3 = 8'd56;
b_mant0 = 8'd240; b_mant1 = 8'd7; b_mant2 = 8'd247; b_mant3 = 8'd243;
a_exp0 = 10'd583; a_exp1 = 10'd343; a_exp2 = 10'd1016; a_exp3 = 10'd147;
b_exp0 = 10'd60; b_exp1 = 10'd487; b_exp2 = 10'd659; b_exp3 = 10'd729;
a_sign0 = 4'd4; a_sign1 = 4'd0; a_sign2 = 4'd8; a_sign3 = 4'd11;
b_sign0 = 4'd4; b_sign1 = 4'd7; b_sign2 = 4'd7; b_sign3 = 4'd14;
@(posedge clk_i);
a_mant0 = 8'd189; a_mant1 = 8'd51; a_mant2 = 8'd217; a_mant3 = 8'd125;
b_mant0 = 8'd72; b_mant1 = 8'd110; b_mant2 = 8'd167; b_mant3 = 8'd109;
a_exp0 = 10'd585; a_exp1 = 10'd111; a_exp2 = 10'd852; a_exp3 = 10'd575;
b_exp0 = 10'd874; b_exp1 = 10'd1016; b_exp2 = 10'd382; b_exp3 = 10'd547;
a_sign0 = 4'd13; a_sign1 = 4'd13; a_sign2 = 4'd14; a_sign3 = 4'd12;
b_sign0 = 4'd5; b_sign1 = 4'd1; b_sign2 = 4'd8; b_sign3 = 4'd12;
@(posedge clk_i);
a_mant0 = 8'd159; a_mant1 = 8'd108; a_mant2 = 8'd86; a_mant3 = 8'd98;
b_mant0 = 8'd39; b_mant1 = 8'd136; b_mant2 = 8'd245; b_mant3 = 8'd80;
a_exp0 = 10'd124; a_exp1 = 10'd913; a_exp2 = 10'd422; a_exp3 = 10'd827;
b_exp0 = 10'd753; b_exp1 = 10'd618; b_exp2 = 10'd92; b_exp3 = 10'd627;
a_sign0 = 4'd0; a_sign1 = 4'd1; a_sign2 = 4'd9; a_sign3 = 4'd2;
b_sign0 = 4'd13; b_sign1 = 4'd8; b_sign2 = 4'd10; b_sign3 = 4'd9;
@(posedge clk_i);
a_mant0 = 8'd153; a_mant1 = 8'd237; a_mant2 = 8'd151; a_mant3 = 8'd87;
b_mant0 = 8'd87; b_mant1 = 8'd12; b_mant2 = 8'd68; b_mant3 = 8'd190;
a_exp0 = 10'd201; a_exp1 = 10'd737; a_exp2 = 10'd220; a_exp3 = 10'd769;
b_exp0 = 10'd781; b_exp1 = 10'd797; b_exp2 = 10'd729; b_exp3 = 10'd915;
a_sign0 = 4'd1; a_sign1 = 4'd3; a_sign2 = 4'd1; a_sign3 = 4'd1;
b_sign0 = 4'd0; b_sign1 = 4'd4; b_sign2 = 4'd8; b_sign3 = 4'd5;
@(posedge clk_i);
shared_exps0 = 8'd112;
shared_exps1 = 8'd128;
a_mant0 = 8'd113; a_mant1 = 8'd3; a_mant2 = 8'd116; a_mant3 = 8'd166;
b_mant0 = 8'd78; b_mant1 = 8'd148; b_mant2 = 8'd241; b_mant3 = 8'd150;
a_exp0 = 10'd924; a_exp1 = 10'd189; a_exp2 = 10'd646; a_exp3 = 10'd292;
b_exp0 = 10'd625; b_exp1 = 10'd873; b_exp2 = 10'd63; b_exp3 = 10'd714;
a_sign0 = 4'd10; a_sign1 = 4'd3; a_sign2 = 4'd0; a_sign3 = 4'd12;
b_sign0 = 4'd0; b_sign1 = 4'd10; b_sign2 = 4'd11; b_sign3 = 4'd15;
@(posedge clk_i);
a_mant0 = 8'd194; a_mant1 = 8'd82; a_mant2 = 8'd4; a_mant3 = 8'd253;
b_mant0 = 8'd80; b_mant1 = 8'd214; b_mant2 = 8'd240; b_mant3 = 8'd85;
a_exp0 = 10'd5; a_exp1 = 10'd634; a_exp2 = 10'd499; a_exp3 = 10'd694;
b_exp0 = 10'd1012; b_exp1 = 10'd52; b_exp2 = 10'd597; b_exp3 = 10'd744;
a_sign0 = 4'd0; a_sign1 = 4'd7; a_sign2 = 4'd11; a_sign3 = 4'd16;
b_sign0 = 4'd2; b_sign1 = 4'd12; b_sign2 = 4'd6; b_sign3 = 4'd9;
@(posedge clk_i);
a_mant0 = 8'd105; a_mant1 = 8'd32; a_mant2 = 8'd188; a_mant3 = 8'd14;
b_mant0 = 8'd207; b_mant1 = 8'd167; b_mant2 = 8'd255; b_mant3 = 8'd109;
a_exp0 = 10'd566; a_exp1 = 10'd26; a_exp2 = 10'd584; a_exp3 = 10'd207;
b_exp0 = 10'd792; b_exp1 = 10'd753; b_exp2 = 10'd483; b_exp3 = 10'd922;
a_sign0 = 4'd2; a_sign1 = 4'd14; a_sign2 = 4'd5; a_sign3 = 4'd12;
b_sign0 = 4'd6; b_sign1 = 4'd14; b_sign2 = 4'd14; b_sign3 = 4'd5;
@(posedge clk_i);
a_mant0 = 8'd248; a_mant1 = 8'd233; a_mant2 = 8'd105; a_mant3 = 8'd120;
b_mant0 = 8'd95; b_mant1 = 8'd191; b_mant2 = 8'd46; b_mant3 = 8'd23;
a_exp0 = 10'd961; a_exp1 = 10'd78; a_exp2 = 10'd896; a_exp3 = 10'd759;
b_exp0 = 10'd25; b_exp1 = 10'd582; b_exp2 = 10'd667; b_exp3 = 10'd820;
a_sign0 = 4'd0; a_sign1 = 4'd13; a_sign2 = 4'd4; a_sign3 = 4'd12;
b_sign0 = 4'd9; b_sign1 = 4'd7; b_sign2 = 4'd15; b_sign3 = 4'd5;
@(posedge clk_i);
a_mant0 = 8'd35; a_mant1 = 8'd177; a_mant2 = 8'd134; a_mant3 = 8'd237;
b_mant0 = 8'd124; b_mant1 = 8'd212; b_mant2 = 8'd190; b_mant3 = 8'd170;
a_exp0 = 10'd405; a_exp1 = 10'd314; a_exp2 = 10'd756; a_exp3 = 10'd860;
b_exp0 = 10'd957; b_exp1 = 10'd914; b_exp2 = 10'd686; b_exp3 = 10'd1021;
a_sign0 = 4'd8; a_sign1 = 4'd0; a_sign2 = 4'd13; a_sign3 = 4'd14;
b_sign0 = 4'd10; b_sign1 = 4'd0; b_sign2 = 4'd2; b_sign3 = 4'd0;
@(posedge clk_i);
a_mant0 = 8'd49; a_mant1 = 8'd191; a_mant2 = 8'd79; a_mant3 = 8'd65;
b_mant0 = 8'd144; b_mant1 = 8'd204; b_mant2 = 8'd134; b_mant3 = 8'd188;
a_exp0 = 10'd485; a_exp1 = 10'd537; a_exp2 = 10'd800; a_exp3 = 10'd400;
b_exp0 = 10'd274; b_exp1 = 10'd793; b_exp2 = 10'd110; b_exp3 = 10'd129;
a_sign0 = 4'd1; a_sign1 = 4'd5; a_sign2 = 4'd10; a_sign3 = 4'd13;
b_sign0 = 4'd7; b_sign1 = 4'd15; b_sign2 = 4'd3; b_sign3 = 4'd6;
@(posedge clk_i);
a_mant0 = 8'd27; a_mant1 = 8'd248; a_mant2 = 8'd149; a_mant3 = 8'd71;
b_mant0 = 8'd177; b_mant1 = 8'd183; b_mant2 = 8'd244; b_mant3 = 8'd89;
a_exp0 = 10'd156; a_exp1 = 10'd310; a_exp2 = 10'd943; a_exp3 = 10'd1004;
b_exp0 = 10'd421; b_exp1 = 10'd449; b_exp2 = 10'd976; b_exp3 = 10'd550;
a_sign0 = 4'd16; a_sign1 = 4'd10; a_sign2 = 4'd2; a_sign3 = 4'd5;
b_sign0 = 4'd3; b_sign1 = 4'd6; b_sign2 = 4'd8; b_sign3 = 4'd0;
@(posedge clk_i);
a_mant0 = 8'd164; a_mant1 = 8'd239; a_mant2 = 8'd187; a_mant3 = 8'd101;
b_mant0 = 8'd248; b_mant1 = 8'd44; b_mant2 = 8'd146; b_mant3 = 8'd83;
a_exp0 = 10'd186; a_exp1 = 10'd793; a_exp2 = 10'd926; a_exp3 = 10'd958;
b_exp0 = 10'd451; b_exp1 = 10'd641; b_exp2 = 10'd872; b_exp3 = 10'd310;
a_sign0 = 4'd3; a_sign1 = 4'd14; a_sign2 = 4'd1; a_sign3 = 4'd4;
b_sign0 = 4'd0; b_sign1 = 4'd8; b_sign2 = 4'd14; b_sign3 = 4'd9;
@(posedge clk_i);
shared_exps0 = 8'd124;
shared_exps1 = 8'd101;
rstn = 0;
@(posedge clk_i);
rstn = 1;
a_mant0 = 8'd255; a_mant1 = 8'd158; a_mant2 = 8'd208; a_mant3 = 8'd215;
b_mant0 = 8'd236; b_mant1 = 8'd15; b_mant2 = 8'd158; b_mant3 = 8'd77;
a_exp0 = 10'd623; a_exp1 = 10'd749; a_exp2 = 10'd59; a_exp3 = 10'd997;
b_exp0 = 10'd578; b_exp1 = 10'd214; b_exp2 = 10'd261; b_exp3 = 10'd726;
a_sign0 = 4'd2; a_sign1 = 4'd1; a_sign2 = 4'd7; a_sign3 = 4'd5;
b_sign0 = 4'd1; b_sign1 = 4'd14; b_sign2 = 4'd15; b_sign3 = 4'd4;
@(posedge clk_i);
a_mant0 = 8'd158; a_mant1 = 8'd160; a_mant2 = 8'd75; a_mant3 = 8'd82;
b_mant0 = 8'd243; b_mant1 = 8'd99; b_mant2 = 8'd102; b_mant3 = 8'd142;
a_exp0 = 10'd371; a_exp1 = 10'd128; a_exp2 = 10'd67; a_exp3 = 10'd425;
b_exp0 = 10'd933; b_exp1 = 10'd581; b_exp2 = 10'd940; b_exp3 = 10'd490;
a_sign0 = 4'd12; a_sign1 = 4'd15; a_sign2 = 4'd14; a_sign3 = 4'd9;
b_sign0 = 4'd3; b_sign1 = 4'd11; b_sign2 = 4'd5; b_sign3 = 4'd9;
@(posedge clk_i);
a_mant0 = 8'd83; a_mant1 = 8'd249; a_mant2 = 8'd181; a_mant3 = 8'd184;
b_mant0 = 8'd11; b_mant1 = 8'd50; b_mant2 = 8'd21; b_mant3 = 8'd116;
a_exp0 = 10'd264; a_exp1 = 10'd711; a_exp2 = 10'd392; a_exp3 = 10'd365;
b_exp0 = 10'd457; b_exp1 = 10'd205; b_exp2 = 10'd765; b_exp3 = 10'd724;
a_sign0 = 4'd5; a_sign1 = 4'd9; a_sign2 = 4'd1; a_sign3 = 4'd1;
b_sign0 = 4'd9; b_sign1 = 4'd8; b_sign2 = 4'd2; b_sign3 = 4'd1;
@(posedge clk_i);
a_mant0 = 8'd107; a_mant1 = 8'd114; a_mant2 = 8'd89; a_mant3 = 8'd226;
b_mant0 = 8'd89; b_mant1 = 8'd207; b_mant2 = 8'd118; b_mant3 = 8'd88;
a_exp0 = 10'd445; a_exp1 = 10'd403; a_exp2 = 10'd275; a_exp3 = 10'd234;
b_exp0 = 10'd213; b_exp1 = 10'd380; b_exp2 = 10'd544; b_exp3 = 10'd884;
a_sign0 = 4'd4; a_sign1 = 4'd15; a_sign2 = 4'd6; a_sign3 = 4'd6;
b_sign0 = 4'd14; b_sign1 = 4'd2; b_sign2 = 4'd15; b_sign3 = 4'd8;
@(posedge clk_i);
a_mant0 = 8'd72; a_mant1 = 8'd48; a_mant2 = 8'd33; a_mant3 = 8'd102;
b_mant0 = 8'd229; b_mant1 = 8'd49; b_mant2 = 8'd124; b_mant3 = 8'd117;
a_exp0 = 10'd18; a_exp1 = 10'd812; a_exp2 = 10'd104; a_exp3 = 10'd410;
b_exp0 = 10'd120; b_exp1 = 10'd321; b_exp2 = 10'd111; b_exp3 = 10'd541;
a_sign0 = 4'd15; a_sign1 = 4'd9; a_sign2 = 4'd5; a_sign3 = 4'd0;
b_sign0 = 4'd15; b_sign1 = 4'd1; b_sign2 = 4'd8; b_sign3 = 4'd3;
@(posedge clk_i);
a_mant0 = 8'd115; a_mant1 = 8'd122; a_mant2 = 8'd90; a_mant3 = 8'd107;
b_mant0 = 8'd203; b_mant1 = 8'd202; b_mant2 = 8'd129; b_mant3 = 8'd13;
a_exp0 = 10'd886; a_exp1 = 10'd135; a_exp2 = 10'd626; a_exp3 = 10'd921;
b_exp0 = 10'd315; b_exp1 = 10'd687; b_exp2 = 10'd1016; b_exp3 = 10'd799;
a_sign0 = 4'd0; a_sign1 = 4'd14; a_sign2 = 4'd2; a_sign3 = 4'd13;
b_sign0 = 4'd1; b_sign1 = 4'd3; b_sign2 = 4'd4; b_sign3 = 4'd6;
@(posedge clk_i);
a_mant0 = 8'd159; a_mant1 = 8'd213; a_mant2 = 8'd211; a_mant3 = 8'd241;
b_mant0 = 8'd50; b_mant1 = 8'd114; b_mant2 = 8'd168; b_mant3 = 8'd13;
a_exp0 = 10'd803; a_exp1 = 10'd131; a_exp2 = 10'd824; a_exp3 = 10'd614;
b_exp0 = 10'd848; b_exp1 = 10'd706; b_exp2 = 10'd273; b_exp3 = 10'd430;
a_sign0 = 4'd13; a_sign1 = 4'd3; a_sign2 = 4'd4; a_sign3 = 4'd3;
b_sign0 = 4'd14; b_sign1 = 4'd7; b_sign2 = 4'd4; b_sign3 = 4'd3;
@(posedge clk_i);
shared_exps0 = 8'd103;
shared_exps1 = 8'd147;
a_mant0 = 8'd41; a_mant1 = 8'd97; a_mant2 = 8'd48; a_mant3 = 8'd98;
b_mant0 = 8'd172; b_mant1 = 8'd74; b_mant2 = 8'd0; b_mant3 = 8'd154;
a_exp0 = 10'd610; a_exp1 = 10'd458; a_exp2 = 10'd864; a_exp3 = 10'd285;
b_exp0 = 10'd359; b_exp1 = 10'd321; b_exp2 = 10'd348; b_exp3 = 10'd239;
a_sign0 = 4'd0; a_sign1 = 4'd3; a_sign2 = 4'd7; a_sign3 = 4'd12;
b_sign0 = 4'd10; b_sign1 = 4'd13; b_sign2 = 4'd3; b_sign3 = 4'd9;
@(posedge clk_i);
a_mant0 = 8'd252; a_mant1 = 8'd214; a_mant2 = 8'd199; a_mant3 = 8'd116;
b_mant0 = 8'd162; b_mant1 = 8'd20; b_mant2 = 8'd189; b_mant3 = 8'd195;
a_exp0 = 10'd828; a_exp1 = 10'd302; a_exp2 = 10'd357; a_exp3 = 10'd263;
b_exp0 = 10'd261; b_exp1 = 10'd528; b_exp2 = 10'd622; b_exp3 = 10'd915;
a_sign0 = 4'd0; a_sign1 = 4'd2; a_sign2 = 4'd1; a_sign3 = 4'd13;
b_sign0 = 4'd0; b_sign1 = 4'd5; b_sign2 = 4'd5; b_sign3 = 4'd6;
@(posedge clk_i);
a_mant0 = 8'd116; a_mant1 = 8'd42; a_mant2 = 8'd144; a_mant3 = 8'd191;
b_mant0 = 8'd255; b_mant1 = 8'd173; b_mant2 = 8'd18; b_mant3 = 8'd55;
a_exp0 = 10'd942; a_exp1 = 10'd336; a_exp2 = 10'd929; a_exp3 = 10'd114;
b_exp0 = 10'd359; b_exp1 = 10'd672; b_exp2 = 10'd645; b_exp3 = 10'd899;
a_sign0 = 4'd3; a_sign1 = 4'd6; a_sign2 = 4'd6; a_sign3 = 4'd15;
b_sign0 = 4'd5; b_sign1 = 4'd3; b_sign2 = 4'd12; b_sign3 = 4'd8;
@(posedge clk_i);
a_mant0 = 8'd203; a_mant1 = 8'd94; a_mant2 = 8'd71; a_mant3 = 8'd22;
b_mant0 = 8'd249; b_mant1 = 8'd4; b_mant2 = 8'd42; b_mant3 = 8'd191;
a_exp0 = 10'd606; a_exp1 = 10'd660; a_exp2 = 10'd327; a_exp3 = 10'd176;
b_exp0 = 10'd215; b_exp1 = 10'd856; b_exp2 = 10'd553; b_exp3 = 10'd57;
a_sign0 = 4'd1; a_sign1 = 4'd11; a_sign2 = 4'd7; a_sign3 = 4'd7;
b_sign0 = 4'd12; b_sign1 = 4'd11; b_sign2 = 4'd6; b_sign3 = 4'd7;
@(posedge clk_i);
a_mant0 = 8'd105; a_mant1 = 8'd7; a_mant2 = 8'd251; a_mant3 = 8'd74;
b_mant0 = 8'd94; b_mant1 = 8'd191; b_mant2 = 8'd205; b_mant3 = 8'd208;
a_exp0 = 10'd577; a_exp1 = 10'd777; a_exp2 = 10'd809; a_exp3 = 10'd410;
b_exp0 = 10'd455; b_exp1 = 10'd278; b_exp2 = 10'd150; b_exp3 = 10'd843;
a_sign0 = 4'd3; a_sign1 = 4'd4; a_sign2 = 4'd6; a_sign3 = 4'd11;
b_sign0 = 4'd11; b_sign1 = 4'd16; b_sign2 = 4'd6; b_sign3 = 4'd1;
@(posedge clk_i);
a_mant0 = 8'd216; a_mant1 = 8'd46; a_mant2 = 8'd240; a_mant3 = 8'd163;
b_mant0 = 8'd147; b_mant1 = 8'd175; b_mant2 = 8'd60; b_mant3 = 8'd124;
a_exp0 = 10'd220; a_exp1 = 10'd494; a_exp2 = 10'd5; a_exp3 = 10'd462;
b_exp0 = 10'd197; b_exp1 = 10'd694; b_exp2 = 10'd43; b_exp3 = 10'd925;
a_sign0 = 4'd16; a_sign1 = 4'd8; a_sign2 = 4'd15; a_sign3 = 4'd13;
b_sign0 = 4'd9; b_sign1 = 4'd12; b_sign2 = 4'd1; b_sign3 = 4'd13;
@(posedge clk_i);
a_mant0 = 8'd192; a_mant1 = 8'd24; a_mant2 = 8'd220; a_mant3 = 8'd207;
b_mant0 = 8'd44; b_mant1 = 8'd12; b_mant2 = 8'd37; b_mant3 = 8'd27;
a_exp0 = 10'd604; a_exp1 = 10'd701; a_exp2 = 10'd748; a_exp3 = 10'd721;
b_exp0 = 10'd371; b_exp1 = 10'd344; b_exp2 = 10'd279; b_exp3 = 10'd38;
a_sign0 = 4'd7; a_sign1 = 4'd4; a_sign2 = 4'd2; a_sign3 = 4'd7;
b_sign0 = 4'd16; b_sign1 = 4'd11; b_sign2 = 4'd11; b_sign3 = 4'd10;
@(posedge clk_i);
a_mant0 = 8'd47; a_mant1 = 8'd29; a_mant2 = 8'd88; a_mant3 = 8'd226;
b_mant0 = 8'd31; b_mant1 = 8'd85; b_mant2 = 8'd81; b_mant3 = 8'd166;
a_exp0 = 10'd658; a_exp1 = 10'd302; a_exp2 = 10'd496; a_exp3 = 10'd982;
b_exp0 = 10'd415; b_exp1 = 10'd610; b_exp2 = 10'd562; b_exp3 = 10'd985;
a_sign0 = 4'd10; a_sign1 = 4'd16; a_sign2 = 4'd11; a_sign3 = 4'd16;
b_sign0 = 4'd10; b_sign1 = 4'd3; b_sign2 = 4'd5; b_sign3 = 4'd11;
@(posedge clk_i);
shared_exps0 = 8'd115;
shared_exps1 = 8'd139;
a_mant0 = 8'd238; a_mant1 = 8'd94; a_mant2 = 8'd177; a_mant3 = 8'd8;
b_mant0 = 8'd143; b_mant1 = 8'd42; b_mant2 = 8'd219; b_mant3 = 8'd119;
a_exp0 = 10'd236; a_exp1 = 10'd441; a_exp2 = 10'd647; a_exp3 = 10'd38;
b_exp0 = 10'd437; b_exp1 = 10'd296; b_exp2 = 10'd630; b_exp3 = 10'd345;
a_sign0 = 4'd12; a_sign1 = 4'd2; a_sign2 = 4'd7; a_sign3 = 4'd16;
b_sign0 = 4'd13; b_sign1 = 4'd3; b_sign2 = 4'd10; b_sign3 = 4'd13;
@(posedge clk_i);
a_mant0 = 8'd146; a_mant1 = 8'd197; a_mant2 = 8'd92; a_mant3 = 8'd164;
b_mant0 = 8'd165; b_mant1 = 8'd29; b_mant2 = 8'd109; b_mant3 = 8'd58;
a_exp0 = 10'd201; a_exp1 = 10'd458; a_exp2 = 10'd240; a_exp3 = 10'd600;
b_exp0 = 10'd599; b_exp1 = 10'd257; b_exp2 = 10'd449; b_exp3 = 10'd449;
a_sign0 = 4'd2; a_sign1 = 4'd6; a_sign2 = 4'd11; a_sign3 = 4'd0;
b_sign0 = 4'd9; b_sign1 = 4'd0; b_sign2 = 4'd0; b_sign3 = 4'd9;
@(posedge clk_i);
a_mant0 = 8'd183; a_mant1 = 8'd77; a_mant2 = 8'd227; a_mant3 = 8'd92;
b_mant0 = 8'd164; b_mant1 = 8'd4; b_mant2 = 8'd24; b_mant3 = 8'd142;
a_exp0 = 10'd95; a_exp1 = 10'd238; a_exp2 = 10'd712; a_exp3 = 10'd411;
b_exp0 = 10'd374; b_exp1 = 10'd476; b_exp2 = 10'd660; b_exp3 = 10'd407;
a_sign0 = 4'd1; a_sign1 = 4'd16; a_sign2 = 4'd8; a_sign3 = 4'd4;
b_sign0 = 4'd11; b_sign1 = 4'd11; b_sign2 = 4'd4; b_sign3 = 4'd1;
@(posedge clk_i);
a_mant0 = 8'd139; a_mant1 = 8'd224; a_mant2 = 8'd134; a_mant3 = 8'd6;
b_mant0 = 8'd120; b_mant1 = 8'd86; b_mant2 = 8'd129; b_mant3 = 8'd78;
a_exp0 = 10'd492; a_exp1 = 10'd419; a_exp2 = 10'd60; a_exp3 = 10'd898;
b_exp0 = 10'd968; b_exp1 = 10'd370; b_exp2 = 10'd32; b_exp3 = 10'd421;
a_sign0 = 4'd13; a_sign1 = 4'd6; a_sign2 = 4'd12; a_sign3 = 4'd9;
b_sign0 = 4'd7; b_sign1 = 4'd11; b_sign2 = 4'd4; b_sign3 = 4'd9;
@(posedge clk_i);
a_mant0 = 8'd145; a_mant1 = 8'd251; a_mant2 = 8'd110; a_mant3 = 8'd15;
b_mant0 = 8'd233; b_mant1 = 8'd124; b_mant2 = 8'd78; b_mant3 = 8'd192;
a_exp0 = 10'd891; a_exp1 = 10'd794; a_exp2 = 10'd956; a_exp3 = 10'd232;
b_exp0 = 10'd356; b_exp1 = 10'd746; b_exp2 = 10'd314; b_exp3 = 10'd840;
a_sign0 = 4'd15; a_sign1 = 4'd2; a_sign2 = 4'd15; a_sign3 = 4'd1;
b_sign0 = 4'd16; b_sign1 = 4'd12; b_sign2 = 4'd5; b_sign3 = 4'd6;
@(posedge clk_i);
a_mant0 = 8'd128; a_mant1 = 8'd66; a_mant2 = 8'd182; a_mant3 = 8'd62;
b_mant0 = 8'd237; b_mant1 = 8'd35; b_mant2 = 8'd2; b_mant3 = 8'd193;
a_exp0 = 10'd427; a_exp1 = 10'd228; a_exp2 = 10'd713; a_exp3 = 10'd945;
b_exp0 = 10'd182; b_exp1 = 10'd838; b_exp2 = 10'd890; b_exp3 = 10'd132;
a_sign0 = 4'd2; a_sign1 = 4'd3; a_sign2 = 4'd14; a_sign3 = 4'd16;
b_sign0 = 4'd5; b_sign1 = 4'd13; b_sign2 = 4'd0; b_sign3 = 4'd15;
@(posedge clk_i);
a_mant0 = 8'd39; a_mant1 = 8'd0; a_mant2 = 8'd210; a_mant3 = 8'd239;
b_mant0 = 8'd134; b_mant1 = 8'd24; b_mant2 = 8'd173; b_mant3 = 8'd48;
a_exp0 = 10'd289; a_exp1 = 10'd279; a_exp2 = 10'd636; a_exp3 = 10'd59;
b_exp0 = 10'd277; b_exp1 = 10'd967; b_exp2 = 10'd554; b_exp3 = 10'd779;
a_sign0 = 4'd15; a_sign1 = 4'd9; a_sign2 = 4'd15; a_sign3 = 4'd1;
b_sign0 = 4'd11; b_sign1 = 4'd10; b_sign2 = 4'd4; b_sign3 = 4'd5;
@(posedge clk_i);
a_mant0 = 8'd13; a_mant1 = 8'd200; a_mant2 = 8'd150; a_mant3 = 8'd193;
b_mant0 = 8'd57; b_mant1 = 8'd122; b_mant2 = 8'd240; b_mant3 = 8'd243;
a_exp0 = 10'd549; a_exp1 = 10'd536; a_exp2 = 10'd785; a_exp3 = 10'd943;
b_exp0 = 10'd728; b_exp1 = 10'd299; b_exp2 = 10'd506; b_exp3 = 10'd564;
a_sign0 = 4'd8; a_sign1 = 4'd4; a_sign2 = 4'd13; a_sign3 = 4'd9;
b_sign0 = 4'd4; b_sign1 = 4'd5; b_sign2 = 4'd7; b_sign3 = 4'd2;
@(posedge clk_i);
shared_exps0 = 8'd118;
shared_exps1 = 8'd104;
a_mant0 = 8'd152; a_mant1 = 8'd131; a_mant2 = 8'd123; a_mant3 = 8'd178;
b_mant0 = 8'd3; b_mant1 = 8'd155; b_mant2 = 8'd205; b_mant3 = 8'd172;
a_exp0 = 10'd930; a_exp1 = 10'd742; a_exp2 = 10'd306; a_exp3 = 10'd550;
b_exp0 = 10'd729; b_exp1 = 10'd300; b_exp2 = 10'd828; b_exp3 = 10'd883;
a_sign0 = 4'd14; a_sign1 = 4'd12; a_sign2 = 4'd13; a_sign3 = 4'd6;
b_sign0 = 4'd4; b_sign1 = 4'd15; b_sign2 = 4'd9; b_sign3 = 4'd11;
@(posedge clk_i);
a_mant0 = 8'd63; a_mant1 = 8'd82; a_mant2 = 8'd193; a_mant3 = 8'd219;
b_mant0 = 8'd116; b_mant1 = 8'd228; b_mant2 = 8'd247; b_mant3 = 8'd37;
a_exp0 = 10'd435; a_exp1 = 10'd11; a_exp2 = 10'd907; a_exp3 = 10'd888;
b_exp0 = 10'd466; b_exp1 = 10'd944; b_exp2 = 10'd996; b_exp3 = 10'd1005;
a_sign0 = 4'd7; a_sign1 = 4'd4; a_sign2 = 4'd3; a_sign3 = 4'd6;
b_sign0 = 4'd4; b_sign1 = 4'd5; b_sign2 = 4'd14; b_sign3 = 4'd12;
@(posedge clk_i);
a_mant0 = 8'd247; a_mant1 = 8'd217; a_mant2 = 8'd37; a_mant3 = 8'd51;
b_mant0 = 8'd172; b_mant1 = 8'd128; b_mant2 = 8'd239; b_mant3 = 8'd92;
a_exp0 = 10'd986; a_exp1 = 10'd636; a_exp2 = 10'd831; a_exp3 = 10'd820;
b_exp0 = 10'd973; b_exp1 = 10'd1; b_exp2 = 10'd816; b_exp3 = 10'd634;
a_sign0 = 4'd8; a_sign1 = 4'd8; a_sign2 = 4'd5; a_sign3 = 4'd4;
b_sign0 = 4'd11; b_sign1 = 4'd11; b_sign2 = 4'd9; b_sign3 = 4'd2;
@(posedge clk_i);
a_mant0 = 8'd40; a_mant1 = 8'd16; a_mant2 = 8'd9; a_mant3 = 8'd218;
b_mant0 = 8'd63; b_mant1 = 8'd4; b_mant2 = 8'd105; b_mant3 = 8'd248;
a_exp0 = 10'd928; a_exp1 = 10'd943; a_exp2 = 10'd460; a_exp3 = 10'd432;
b_exp0 = 10'd415; b_exp1 = 10'd882; b_exp2 = 10'd910; b_exp3 = 10'd768;
a_sign0 = 4'd13; a_sign1 = 4'd13; a_sign2 = 4'd6; a_sign3 = 4'd3;
b_sign0 = 4'd11; b_sign1 = 4'd11; b_sign2 = 4'd5; b_sign3 = 4'd15;
@(posedge clk_i);
a_mant0 = 8'd186; a_mant1 = 8'd41; a_mant2 = 8'd153; a_mant3 = 8'd171;
b_mant0 = 8'd110; b_mant1 = 8'd219; b_mant2 = 8'd60; b_mant3 = 8'd182;
a_exp0 = 10'd236; a_exp1 = 10'd715; a_exp2 = 10'd263; a_exp3 = 10'd887;
b_exp0 = 10'd133; b_exp1 = 10'd262; b_exp2 = 10'd163; b_exp3 = 10'd277;
a_sign0 = 4'd15; a_sign1 = 4'd0; a_sign2 = 4'd6; a_sign3 = 4'd11;
b_sign0 = 4'd14; b_sign1 = 4'd11; b_sign2 = 4'd9; b_sign3 = 4'd2;
@(posedge clk_i);
a_mant0 = 8'd21; a_mant1 = 8'd199; a_mant2 = 8'd151; a_mant3 = 8'd199;
b_mant0 = 8'd37; b_mant1 = 8'd56; b_mant2 = 8'd145; b_mant3 = 8'd71;
a_exp0 = 10'd800; a_exp1 = 10'd138; a_exp2 = 10'd744; a_exp3 = 10'd556;
b_exp0 = 10'd420; b_exp1 = 10'd876; b_exp2 = 10'd585; b_exp3 = 10'd797;
a_sign0 = 4'd4; a_sign1 = 4'd5; a_sign2 = 4'd5; a_sign3 = 4'd14;
b_sign0 = 4'd13; b_sign1 = 4'd14; b_sign2 = 4'd13; b_sign3 = 4'd14;
@(posedge clk_i);
a_mant0 = 8'd167; a_mant1 = 8'd175; a_mant2 = 8'd91; a_mant3 = 8'd228;
b_mant0 = 8'd200; b_mant1 = 8'd190; b_mant2 = 8'd171; b_mant3 = 8'd131;
a_exp0 = 10'd578; a_exp1 = 10'd410; a_exp2 = 10'd811; a_exp3 = 10'd551;
b_exp0 = 10'd337; b_exp1 = 10'd775; b_exp2 = 10'd774; b_exp3 = 10'd161;
a_sign0 = 4'd2; a_sign1 = 4'd6; a_sign2 = 4'd1; a_sign3 = 4'd13;
b_sign0 = 4'd6; b_sign1 = 4'd14; b_sign2 = 4'd13; b_sign3 = 4'd0;
@(posedge clk_i);
a_mant0 = 8'd129; a_mant1 = 8'd44; a_mant2 = 8'd235; a_mant3 = 8'd168;
b_mant0 = 8'd189; b_mant1 = 8'd115; b_mant2 = 8'd174; b_mant3 = 8'd143;
a_exp0 = 10'd827; a_exp1 = 10'd899; a_exp2 = 10'd505; a_exp3 = 10'd938;
b_exp0 = 10'd168; b_exp1 = 10'd444; b_exp2 = 10'd410; b_exp3 = 10'd206;
a_sign0 = 4'd14; a_sign1 = 4'd3; a_sign2 = 4'd0; a_sign3 = 4'd2;
b_sign0 = 4'd15; b_sign1 = 4'd2; b_sign2 = 4'd10; b_sign3 = 4'd12;
@(posedge clk_i);
shared_exps0 = 8'd110;
shared_exps1 = 8'd137;
rstn = 0;
@(posedge clk_i);
rstn = 1;
a_mant0 = 8'd10; a_mant1 = 8'd161; a_mant2 = 8'd40; a_mant3 = 8'd234;
b_mant0 = 8'd147; b_mant1 = 8'd102; b_mant2 = 8'd13; b_mant3 = 8'd75;
a_exp0 = 10'd298; a_exp1 = 10'd162; a_exp2 = 10'd90; a_exp3 = 10'd141;
b_exp0 = 10'd574; b_exp1 = 10'd831; b_exp2 = 10'd655; b_exp3 = 10'd442;
a_sign0 = 4'd6; a_sign1 = 4'd1; a_sign2 = 4'd4; a_sign3 = 4'd13;
b_sign0 = 4'd15; b_sign1 = 4'd16; b_sign2 = 4'd10; b_sign3 = 4'd2;
@(posedge clk_i);
a_mant0 = 8'd226; a_mant1 = 8'd77; a_mant2 = 8'd95; a_mant3 = 8'd223;
b_mant0 = 8'd224; b_mant1 = 8'd110; b_mant2 = 8'd70; b_mant3 = 8'd2;
a_exp0 = 10'd733; a_exp1 = 10'd92; a_exp2 = 10'd51; a_exp3 = 10'd67;
b_exp0 = 10'd166; b_exp1 = 10'd153; b_exp2 = 10'd471; b_exp3 = 10'd1013;
a_sign0 = 4'd9; a_sign1 = 4'd13; a_sign2 = 4'd3; a_sign3 = 4'd14;
b_sign0 = 4'd9; b_sign1 = 4'd0; b_sign2 = 4'd1; b_sign3 = 4'd8;
@(posedge clk_i);
a_mant0 = 8'd229; a_mant1 = 8'd112; a_mant2 = 8'd35; a_mant3 = 8'd22;
b_mant0 = 8'd53; b_mant1 = 8'd48; b_mant2 = 8'd150; b_mant3 = 8'd51;
a_exp0 = 10'd568; a_exp1 = 10'd364; a_exp2 = 10'd309; a_exp3 = 10'd182;
b_exp0 = 10'd830; b_exp1 = 10'd965; b_exp2 = 10'd728; b_exp3 = 10'd943;
a_sign0 = 4'd13; a_sign1 = 4'd1; a_sign2 = 4'd5; a_sign3 = 4'd4;
b_sign0 = 4'd2; b_sign1 = 4'd3; b_sign2 = 4'd1; b_sign3 = 4'd13;
@(posedge clk_i);
a_mant0 = 8'd118; a_mant1 = 8'd135; a_mant2 = 8'd51; a_mant3 = 8'd152;
b_mant0 = 8'd102; b_mant1 = 8'd156; b_mant2 = 8'd31; b_mant3 = 8'd48;
a_exp0 = 10'd116; a_exp1 = 10'd833; a_exp2 = 10'd130; a_exp3 = 10'd13;
b_exp0 = 10'd118; b_exp1 = 10'd335; b_exp2 = 10'd573; b_exp3 = 10'd1020;
a_sign0 = 4'd3; a_sign1 = 4'd5; a_sign2 = 4'd11; a_sign3 = 4'd0;
b_sign0 = 4'd15; b_sign1 = 4'd16; b_sign2 = 4'd13; b_sign3 = 4'd0;
@(posedge clk_i);
a_mant0 = 8'd219; a_mant1 = 8'd99; a_mant2 = 8'd98; a_mant3 = 8'd170;
b_mant0 = 8'd158; b_mant1 = 8'd64; b_mant2 = 8'd147; b_mant3 = 8'd216;
a_exp0 = 10'd352; a_exp1 = 10'd30; a_exp2 = 10'd212; a_exp3 = 10'd771;
b_exp0 = 10'd947; b_exp1 = 10'd441; b_exp2 = 10'd879; b_exp3 = 10'd373;
a_sign0 = 4'd9; a_sign1 = 4'd8; a_sign2 = 4'd10; a_sign3 = 4'd15;
b_sign0 = 4'd0; b_sign1 = 4'd6; b_sign2 = 4'd11; b_sign3 = 4'd13;
@(posedge clk_i);
a_mant0 = 8'd114; a_mant1 = 8'd120; a_mant2 = 8'd36; a_mant3 = 8'd115;
b_mant0 = 8'd245; b_mant1 = 8'd36; b_mant2 = 8'd185; b_mant3 = 8'd245;
a_exp0 = 10'd25; a_exp1 = 10'd873; a_exp2 = 10'd302; a_exp3 = 10'd468;
b_exp0 = 10'd68; b_exp1 = 10'd244; b_exp2 = 10'd428; b_exp3 = 10'd211;
a_sign0 = 4'd10; a_sign1 = 4'd6; a_sign2 = 4'd1; a_sign3 = 4'd11;
b_sign0 = 4'd1; b_sign1 = 4'd8; b_sign2 = 4'd5; b_sign3 = 4'd16;
@(posedge clk_i);
a_mant0 = 8'd140; a_mant1 = 8'd32; a_mant2 = 8'd225; a_mant3 = 8'd76;
b_mant0 = 8'd118; b_mant1 = 8'd133; b_mant2 = 8'd234; b_mant3 = 8'd137;
a_exp0 = 10'd298; a_exp1 = 10'd29; a_exp2 = 10'd177; a_exp3 = 10'd215;
b_exp0 = 10'd115; b_exp1 = 10'd891; b_exp2 = 10'd671; b_exp3 = 10'd317;
a_sign0 = 4'd0; a_sign1 = 4'd0; a_sign2 = 4'd5; a_sign3 = 4'd11;
b_sign0 = 4'd4; b_sign1 = 4'd12; b_sign2 = 4'd6; b_sign3 = 4'd10;
@(posedge clk_i);
shared_exps0 = 8'd131;
shared_exps1 = 8'd110;
a_mant0 = 8'd35; a_mant1 = 8'd123; a_mant2 = 8'd139; a_mant3 = 8'd176;
b_mant0 = 8'd60; b_mant1 = 8'd12; b_mant2 = 8'd142; b_mant3 = 8'd224;
a_exp0 = 10'd399; a_exp1 = 10'd53; a_exp2 = 10'd211; a_exp3 = 10'd872;
b_exp0 = 10'd145; b_exp1 = 10'd469; b_exp2 = 10'd378; b_exp3 = 10'd300;
a_sign0 = 4'd8; a_sign1 = 4'd15; a_sign2 = 4'd3; a_sign3 = 4'd16;
b_sign0 = 4'd2; b_sign1 = 4'd13; b_sign2 = 4'd6; b_sign3 = 4'd13;
@(posedge clk_i);
a_mant0 = 8'd254; a_mant1 = 8'd118; a_mant2 = 8'd220; a_mant3 = 8'd42;
b_mant0 = 8'd217; b_mant1 = 8'd108; b_mant2 = 8'd71; b_mant3 = 8'd57;
a_exp0 = 10'd945; a_exp1 = 10'd623; a_exp2 = 10'd742; a_exp3 = 10'd59;
b_exp0 = 10'd424; b_exp1 = 10'd68; b_exp2 = 10'd902; b_exp3 = 10'd421;
a_sign0 = 4'd7; a_sign1 = 4'd13; a_sign2 = 4'd9; a_sign3 = 4'd7;
b_sign0 = 4'd11; b_sign1 = 4'd11; b_sign2 = 4'd10; b_sign3 = 4'd15;
@(posedge clk_i);
a_mant0 = 8'd82; a_mant1 = 8'd61; a_mant2 = 8'd226; a_mant3 = 8'd136;
b_mant0 = 8'd48; b_mant1 = 8'd32; b_mant2 = 8'd142; b_mant3 = 8'd97;
a_exp0 = 10'd706; a_exp1 = 10'd790; a_exp2 = 10'd864; a_exp3 = 10'd141;
b_exp0 = 10'd160; b_exp1 = 10'd479; b_exp2 = 10'd49; b_exp3 = 10'd963;
a_sign0 = 4'd1; a_sign1 = 4'd10; a_sign2 = 4'd13; a_sign3 = 4'd5;
b_sign0 = 4'd12; b_sign1 = 4'd11; b_sign2 = 4'd4; b_sign3 = 4'd12;
@(posedge clk_i);
a_mant0 = 8'd195; a_mant1 = 8'd62; a_mant2 = 8'd210; a_mant3 = 8'd29;
b_mant0 = 8'd48; b_mant1 = 8'd4; b_mant2 = 8'd63; b_mant3 = 8'd40;
a_exp0 = 10'd494; a_exp1 = 10'd813; a_exp2 = 10'd529; a_exp3 = 10'd719;
b_exp0 = 10'd515; b_exp1 = 10'd964; b_exp2 = 10'd934; b_exp3 = 10'd506;
a_sign0 = 4'd3; a_sign1 = 4'd2; a_sign2 = 4'd13; a_sign3 = 4'd13;
b_sign0 = 4'd0; b_sign1 = 4'd1; b_sign2 = 4'd9; b_sign3 = 4'd7;
@(posedge clk_i);
a_mant0 = 8'd9; a_mant1 = 8'd31; a_mant2 = 8'd132; a_mant3 = 8'd199;
b_mant0 = 8'd154; b_mant1 = 8'd243; b_mant2 = 8'd5; b_mant3 = 8'd70;
a_exp0 = 10'd408; a_exp1 = 10'd630; a_exp2 = 10'd194; a_exp3 = 10'd365;
b_exp0 = 10'd592; b_exp1 = 10'd462; b_exp2 = 10'd357; b_exp3 = 10'd859;
a_sign0 = 4'd3; a_sign1 = 4'd12; a_sign2 = 4'd5; a_sign3 = 4'd3;
b_sign0 = 4'd5; b_sign1 = 4'd12; b_sign2 = 4'd16; b_sign3 = 4'd6;
@(posedge clk_i);
a_mant0 = 8'd243; a_mant1 = 8'd205; a_mant2 = 8'd116; a_mant3 = 8'd65;
b_mant0 = 8'd70; b_mant1 = 8'd189; b_mant2 = 8'd202; b_mant3 = 8'd147;
a_exp0 = 10'd492; a_exp1 = 10'd990; a_exp2 = 10'd719; a_exp3 = 10'd971;
b_exp0 = 10'd360; b_exp1 = 10'd217; b_exp2 = 10'd744; b_exp3 = 10'd929;
a_sign0 = 4'd7; a_sign1 = 4'd3; a_sign2 = 4'd5; a_sign3 = 4'd10;
b_sign0 = 4'd10; b_sign1 = 4'd4; b_sign2 = 4'd7; b_sign3 = 4'd2;
@(posedge clk_i);
a_mant0 = 8'd157; a_mant1 = 8'd11; a_mant2 = 8'd198; a_mant3 = 8'd74;
b_mant0 = 8'd149; b_mant1 = 8'd83; b_mant2 = 8'd19; b_mant3 = 8'd77;
a_exp0 = 10'd507; a_exp1 = 10'd780; a_exp2 = 10'd795; a_exp3 = 10'd685;
b_exp0 = 10'd804; b_exp1 = 10'd978; b_exp2 = 10'd845; b_exp3 = 10'd290;
a_sign0 = 4'd9; a_sign1 = 4'd9; a_sign2 = 4'd7; a_sign3 = 4'd11;
b_sign0 = 4'd15; b_sign1 = 4'd13; b_sign2 = 4'd4; b_sign3 = 4'd4;
@(posedge clk_i);
a_mant0 = 8'd43; a_mant1 = 8'd211; a_mant2 = 8'd173; a_mant3 = 8'd49;
b_mant0 = 8'd204; b_mant1 = 8'd177; b_mant2 = 8'd255; b_mant3 = 8'd187;
a_exp0 = 10'd1021; a_exp1 = 10'd239; a_exp2 = 10'd262; a_exp3 = 10'd909;
b_exp0 = 10'd116; b_exp1 = 10'd351; b_exp2 = 10'd283; b_exp3 = 10'd902;
a_sign0 = 4'd15; a_sign1 = 4'd6; a_sign2 = 4'd16; a_sign3 = 4'd1;
b_sign0 = 4'd6; b_sign1 = 4'd11; b_sign2 = 4'd13; b_sign3 = 4'd3;
@(posedge clk_i);
shared_exps0 = 8'd153;
shared_exps1 = 8'd137;
a_mant0 = 8'd211; a_mant1 = 8'd92; a_mant2 = 8'd54; a_mant3 = 8'd35;
b_mant0 = 8'd7; b_mant1 = 8'd151; b_mant2 = 8'd36; b_mant3 = 8'd44;
a_exp0 = 10'd31; a_exp1 = 10'd492; a_exp2 = 10'd898; a_exp3 = 10'd774;
b_exp0 = 10'd335; b_exp1 = 10'd793; b_exp2 = 10'd609; b_exp3 = 10'd69;
a_sign0 = 4'd11; a_sign1 = 4'd3; a_sign2 = 4'd10; a_sign3 = 4'd5;
b_sign0 = 4'd16; b_sign1 = 4'd16; b_sign2 = 4'd3; b_sign3 = 4'd16;
@(posedge clk_i);
a_mant0 = 8'd229; a_mant1 = 8'd249; a_mant2 = 8'd197; a_mant3 = 8'd170;
b_mant0 = 8'd12; b_mant1 = 8'd48; b_mant2 = 8'd232; b_mant3 = 8'd160;
a_exp0 = 10'd152; a_exp1 = 10'd816; a_exp2 = 10'd989; a_exp3 = 10'd561;
b_exp0 = 10'd91; b_exp1 = 10'd456; b_exp2 = 10'd338; b_exp3 = 10'd285;
a_sign0 = 4'd14; a_sign1 = 4'd10; a_sign2 = 4'd10; a_sign3 = 4'd4;
b_sign0 = 4'd3; b_sign1 = 4'd3; b_sign2 = 4'd11; b_sign3 = 4'd13;
@(posedge clk_i);
a_mant0 = 8'd50; a_mant1 = 8'd52; a_mant2 = 8'd1; a_mant3 = 8'd164;
b_mant0 = 8'd62; b_mant1 = 8'd78; b_mant2 = 8'd92; b_mant3 = 8'd244;
a_exp0 = 10'd39; a_exp1 = 10'd95; a_exp2 = 10'd8; a_exp3 = 10'd262;
b_exp0 = 10'd379; b_exp1 = 10'd280; b_exp2 = 10'd50; b_exp3 = 10'd484;
a_sign0 = 4'd15; a_sign1 = 4'd14; a_sign2 = 4'd15; a_sign3 = 4'd7;
b_sign0 = 4'd12; b_sign1 = 4'd6; b_sign2 = 4'd3; b_sign3 = 4'd0;
@(posedge clk_i);
a_mant0 = 8'd232; a_mant1 = 8'd99; a_mant2 = 8'd19; a_mant3 = 8'd192;
b_mant0 = 8'd3; b_mant1 = 8'd182; b_mant2 = 8'd212; b_mant3 = 8'd75;
a_exp0 = 10'd756; a_exp1 = 10'd295; a_exp2 = 10'd206; a_exp3 = 10'd154;
b_exp0 = 10'd303; b_exp1 = 10'd61; b_exp2 = 10'd863; b_exp3 = 10'd615;
a_sign0 = 4'd2; a_sign1 = 4'd6; a_sign2 = 4'd16; a_sign3 = 4'd7;
b_sign0 = 4'd16; b_sign1 = 4'd6; b_sign2 = 4'd15; b_sign3 = 4'd4;
@(posedge clk_i);
a_mant0 = 8'd84; a_mant1 = 8'd177; a_mant2 = 8'd155; a_mant3 = 8'd81;
b_mant0 = 8'd136; b_mant1 = 8'd185; b_mant2 = 8'd249; b_mant3 = 8'd157;
a_exp0 = 10'd179; a_exp1 = 10'd1016; a_exp2 = 10'd287; a_exp3 = 10'd308;
b_exp0 = 10'd241; b_exp1 = 10'd15; b_exp2 = 10'd15; b_exp3 = 10'd713;
a_sign0 = 4'd2; a_sign1 = 4'd10; a_sign2 = 4'd11; a_sign3 = 4'd2;
b_sign0 = 4'd15; b_sign1 = 4'd5; b_sign2 = 4'd3; b_sign3 = 4'd6;
@(posedge clk_i);
a_mant0 = 8'd26; a_mant1 = 8'd2; a_mant2 = 8'd216; a_mant3 = 8'd186;
b_mant0 = 8'd70; b_mant1 = 8'd172; b_mant2 = 8'd196; b_mant3 = 8'd234;
a_exp0 = 10'd655; a_exp1 = 10'd569; a_exp2 = 10'd425; a_exp3 = 10'd597;
b_exp0 = 10'd569; b_exp1 = 10'd500; b_exp2 = 10'd361; b_exp3 = 10'd474;
a_sign0 = 4'd10; a_sign1 = 4'd13; a_sign2 = 4'd6; a_sign3 = 4'd15;
b_sign0 = 4'd2; b_sign1 = 4'd16; b_sign2 = 4'd12; b_sign3 = 4'd4;
@(posedge clk_i);
a_mant0 = 8'd158; a_mant1 = 8'd145; a_mant2 = 8'd140; a_mant3 = 8'd37;
b_mant0 = 8'd162; b_mant1 = 8'd202; b_mant2 = 8'd85; b_mant3 = 8'd135;
a_exp0 = 10'd606; a_exp1 = 10'd680; a_exp2 = 10'd619; a_exp3 = 10'd304;
b_exp0 = 10'd723; b_exp1 = 10'd624; b_exp2 = 10'd290; b_exp3 = 10'd596;
a_sign0 = 4'd10; a_sign1 = 4'd6; a_sign2 = 4'd8; a_sign3 = 4'd1;
b_sign0 = 4'd8; b_sign1 = 4'd3; b_sign2 = 4'd13; b_sign3 = 4'd8;
@(posedge clk_i);
a_mant0 = 8'd120; a_mant1 = 8'd29; a_mant2 = 8'd217; a_mant3 = 8'd76;
b_mant0 = 8'd101; b_mant1 = 8'd177; b_mant2 = 8'd141; b_mant3 = 8'd137;
a_exp0 = 10'd147; a_exp1 = 10'd521; a_exp2 = 10'd290; a_exp3 = 10'd631;
b_exp0 = 10'd610; b_exp1 = 10'd719; b_exp2 = 10'd778; b_exp3 = 10'd27;
a_sign0 = 4'd15; a_sign1 = 4'd2; a_sign2 = 4'd4; a_sign3 = 4'd12;
b_sign0 = 4'd8; b_sign1 = 4'd5; b_sign2 = 4'd8; b_sign3 = 4'd7;
@(posedge clk_i);
shared_exps0 = 8'd120;
shared_exps1 = 8'd123;
a_mant0 = 8'd175; a_mant1 = 8'd91; a_mant2 = 8'd51; a_mant3 = 8'd50;
b_mant0 = 8'd44; b_mant1 = 8'd133; b_mant2 = 8'd221; b_mant3 = 8'd191;
a_exp0 = 10'd197; a_exp1 = 10'd791; a_exp2 = 10'd934; a_exp3 = 10'd676;
b_exp0 = 10'd632; b_exp1 = 10'd813; b_exp2 = 10'd197; b_exp3 = 10'd450;
a_sign0 = 4'd1; a_sign1 = 4'd0; a_sign2 = 4'd0; a_sign3 = 4'd11;
b_sign0 = 4'd6; b_sign1 = 4'd4; b_sign2 = 4'd5; b_sign3 = 4'd12;
@(posedge clk_i);
a_mant0 = 8'd76; a_mant1 = 8'd58; a_mant2 = 8'd16; a_mant3 = 8'd48;
b_mant0 = 8'd8; b_mant1 = 8'd3; b_mant2 = 8'd127; b_mant3 = 8'd201;
a_exp0 = 10'd64; a_exp1 = 10'd680; a_exp2 = 10'd601; a_exp3 = 10'd49;
b_exp0 = 10'd563; b_exp1 = 10'd600; b_exp2 = 10'd206; b_exp3 = 10'd203;
a_sign0 = 4'd5; a_sign1 = 4'd6; a_sign2 = 4'd8; a_sign3 = 4'd11;
b_sign0 = 4'd4; b_sign1 = 4'd3; b_sign2 = 4'd2; b_sign3 = 4'd3;
@(posedge clk_i);
a_mant0 = 8'd19; a_mant1 = 8'd59; a_mant2 = 8'd22; a_mant3 = 8'd218;
b_mant0 = 8'd190; b_mant1 = 8'd163; b_mant2 = 8'd156; b_mant3 = 8'd63;
a_exp0 = 10'd325; a_exp1 = 10'd919; a_exp2 = 10'd507; a_exp3 = 10'd869;
b_exp0 = 10'd550; b_exp1 = 10'd271; b_exp2 = 10'd943; b_exp3 = 10'd176;
a_sign0 = 4'd7; a_sign1 = 4'd7; a_sign2 = 4'd14; a_sign3 = 4'd15;
b_sign0 = 4'd13; b_sign1 = 4'd4; b_sign2 = 4'd15; b_sign3 = 4'd12;
@(posedge clk_i);
a_mant0 = 8'd83; a_mant1 = 8'd106; a_mant2 = 8'd87; a_mant3 = 8'd58;
b_mant0 = 8'd2; b_mant1 = 8'd76; b_mant2 = 8'd191; b_mant3 = 8'd76;
a_exp0 = 10'd582; a_exp1 = 10'd399; a_exp2 = 10'd196; a_exp3 = 10'd584;
b_exp0 = 10'd403; b_exp1 = 10'd323; b_exp2 = 10'd469; b_exp3 = 10'd25;
a_sign0 = 4'd9; a_sign1 = 4'd7; a_sign2 = 4'd4; a_sign3 = 4'd13;
b_sign0 = 4'd2; b_sign1 = 4'd2; b_sign2 = 4'd7; b_sign3 = 4'd7;
@(posedge clk_i);
a_mant0 = 8'd187; a_mant1 = 8'd35; a_mant2 = 8'd101; a_mant3 = 8'd49;
b_mant0 = 8'd209; b_mant1 = 8'd150; b_mant2 = 8'd235; b_mant3 = 8'd116;
a_exp0 = 10'd220; a_exp1 = 10'd26; a_exp2 = 10'd337; a_exp3 = 10'd219;
b_exp0 = 10'd48; b_exp1 = 10'd574; b_exp2 = 10'd64; b_exp3 = 10'd863;
a_sign0 = 4'd14; a_sign1 = 4'd5; a_sign2 = 4'd11; a_sign3 = 4'd4;
b_sign0 = 4'd11; b_sign1 = 4'd9; b_sign2 = 4'd4; b_sign3 = 4'd15;
@(posedge clk_i);
a_mant0 = 8'd83; a_mant1 = 8'd254; a_mant2 = 8'd221; a_mant3 = 8'd252;
b_mant0 = 8'd101; b_mant1 = 8'd67; b_mant2 = 8'd113; b_mant3 = 8'd138;
a_exp0 = 10'd105; a_exp1 = 10'd991; a_exp2 = 10'd748; a_exp3 = 10'd601;
b_exp0 = 10'd84; b_exp1 = 10'd694; b_exp2 = 10'd51; b_exp3 = 10'd52;
a_sign0 = 4'd16; a_sign1 = 4'd2; a_sign2 = 4'd11; a_sign3 = 4'd9;
b_sign0 = 4'd13; b_sign1 = 4'd1; b_sign2 = 4'd2; b_sign3 = 4'd14;
@(posedge clk_i);
a_mant0 = 8'd114; a_mant1 = 8'd178; a_mant2 = 8'd15; a_mant3 = 8'd165;
b_mant0 = 8'd172; b_mant1 = 8'd101; b_mant2 = 8'd125; b_mant3 = 8'd171;
a_exp0 = 10'd927; a_exp1 = 10'd181; a_exp2 = 10'd124; a_exp3 = 10'd376;
b_exp0 = 10'd80; b_exp1 = 10'd297; b_exp2 = 10'd701; b_exp3 = 10'd522;
a_sign0 = 4'd7; a_sign1 = 4'd9; a_sign2 = 4'd3; a_sign3 = 4'd15;
b_sign0 = 4'd7; b_sign1 = 4'd6; b_sign2 = 4'd1; b_sign3 = 4'd16;
@(posedge clk_i);
a_mant0 = 8'd232; a_mant1 = 8'd158; a_mant2 = 8'd17; a_mant3 = 8'd145;
b_mant0 = 8'd119; b_mant1 = 8'd145; b_mant2 = 8'd70; b_mant3 = 8'd253;
a_exp0 = 10'd968; a_exp1 = 10'd603; a_exp2 = 10'd579; a_exp3 = 10'd230;
b_exp0 = 10'd736; b_exp1 = 10'd454; b_exp2 = 10'd729; b_exp3 = 10'd996;
a_sign0 = 4'd12; a_sign1 = 4'd10; a_sign2 = 4'd10; a_sign3 = 4'd13;
b_sign0 = 4'd12; b_sign1 = 4'd4; b_sign2 = 4'd0; b_sign3 = 4'd1;
@(posedge clk_i);
shared_exps0 = 8'd129;
shared_exps1 = 8'd112;
rstn = 0;
@(posedge clk_i);
rstn = 1;
a_mant0 = 8'd77; a_mant1 = 8'd81; a_mant2 = 8'd235; a_mant3 = 8'd33;
b_mant0 = 8'd251; b_mant1 = 8'd1; b_mant2 = 8'd228; b_mant3 = 8'd63;
a_exp0 = 10'd680; a_exp1 = 10'd183; a_exp2 = 10'd80; a_exp3 = 10'd97;
b_exp0 = 10'd809; b_exp1 = 10'd1006; b_exp2 = 10'd444; b_exp3 = 10'd586;
a_sign0 = 4'd3; a_sign1 = 4'd12; a_sign2 = 4'd12; a_sign3 = 4'd9;
b_sign0 = 4'd10; b_sign1 = 4'd2; b_sign2 = 4'd13; b_sign3 = 4'd10;
@(posedge clk_i);
a_mant0 = 8'd2; a_mant1 = 8'd11; a_mant2 = 8'd210; a_mant3 = 8'd180;
b_mant0 = 8'd27; b_mant1 = 8'd239; b_mant2 = 8'd14; b_mant3 = 8'd42;
a_exp0 = 10'd317; a_exp1 = 10'd293; a_exp2 = 10'd301; a_exp3 = 10'd140;
b_exp0 = 10'd665; b_exp1 = 10'd565; b_exp2 = 10'd827; b_exp3 = 10'd748;
a_sign0 = 4'd11; a_sign1 = 4'd1; a_sign2 = 4'd15; a_sign3 = 4'd9;
b_sign0 = 4'd14; b_sign1 = 4'd5; b_sign2 = 4'd10; b_sign3 = 4'd15;
@(posedge clk_i);
a_mant0 = 8'd65; a_mant1 = 8'd17; a_mant2 = 8'd36; a_mant3 = 8'd245;
b_mant0 = 8'd19; b_mant1 = 8'd59; b_mant2 = 8'd177; b_mant3 = 8'd218;
a_exp0 = 10'd719; a_exp1 = 10'd203; a_exp2 = 10'd111; a_exp3 = 10'd388;
b_exp0 = 10'd2; b_exp1 = 10'd59; b_exp2 = 10'd804; b_exp3 = 10'd1022;
a_sign0 = 4'd12; a_sign1 = 4'd2; a_sign2 = 4'd3; a_sign3 = 4'd4;
b_sign0 = 4'd10; b_sign1 = 4'd12; b_sign2 = 4'd16; b_sign3 = 4'd11;
@(posedge clk_i);
a_mant0 = 8'd91; a_mant1 = 8'd210; a_mant2 = 8'd27; a_mant3 = 8'd153;
b_mant0 = 8'd191; b_mant1 = 8'd29; b_mant2 = 8'd249; b_mant3 = 8'd37;
a_exp0 = 10'd687; a_exp1 = 10'd98; a_exp2 = 10'd1011; a_exp3 = 10'd1001;
b_exp0 = 10'd381; b_exp1 = 10'd843; b_exp2 = 10'd530; b_exp3 = 10'd820;
a_sign0 = 4'd1; a_sign1 = 4'd3; a_sign2 = 4'd11; a_sign3 = 4'd8;
b_sign0 = 4'd4; b_sign1 = 4'd2; b_sign2 = 4'd16; b_sign3 = 4'd5;
@(posedge clk_i);
a_mant0 = 8'd117; a_mant1 = 8'd27; a_mant2 = 8'd23; a_mant3 = 8'd61;
b_mant0 = 8'd246; b_mant1 = 8'd164; b_mant2 = 8'd117; b_mant3 = 8'd77;
a_exp0 = 10'd665; a_exp1 = 10'd97; a_exp2 = 10'd807; a_exp3 = 10'd947;
b_exp0 = 10'd469; b_exp1 = 10'd388; b_exp2 = 10'd343; b_exp3 = 10'd852;
a_sign0 = 4'd6; a_sign1 = 4'd10; a_sign2 = 4'd4; a_sign3 = 4'd12;
b_sign0 = 4'd1; b_sign1 = 4'd1; b_sign2 = 4'd11; b_sign3 = 4'd12;
@(posedge clk_i);
a_mant0 = 8'd169; a_mant1 = 8'd107; a_mant2 = 8'd192; a_mant3 = 8'd139;
b_mant0 = 8'd40; b_mant1 = 8'd223; b_mant2 = 8'd74; b_mant3 = 8'd26;
a_exp0 = 10'd729; a_exp1 = 10'd145; a_exp2 = 10'd237; a_exp3 = 10'd696;
b_exp0 = 10'd877; b_exp1 = 10'd745; b_exp2 = 10'd594; b_exp3 = 10'd358;
a_sign0 = 4'd7; a_sign1 = 4'd16; a_sign2 = 4'd9; a_sign3 = 4'd13;
b_sign0 = 4'd13; b_sign1 = 4'd7; b_sign2 = 4'd9; b_sign3 = 4'd2;
@(posedge clk_i);
a_mant0 = 8'd89; a_mant1 = 8'd14; a_mant2 = 8'd114; a_mant3 = 8'd29;
b_mant0 = 8'd52; b_mant1 = 8'd79; b_mant2 = 8'd60; b_mant3 = 8'd179;
a_exp0 = 10'd587; a_exp1 = 10'd978; a_exp2 = 10'd472; a_exp3 = 10'd622;
b_exp0 = 10'd3; b_exp1 = 10'd421; b_exp2 = 10'd305; b_exp3 = 10'd987;
a_sign0 = 4'd15; a_sign1 = 4'd16; a_sign2 = 4'd14; a_sign3 = 4'd8;
b_sign0 = 4'd7; b_sign1 = 4'd3; b_sign2 = 4'd2; b_sign3 = 4'd11;
@(posedge clk_i);
shared_exps0 = 8'd123;
shared_exps1 = 8'd122;
a_mant0 = 8'd38; a_mant1 = 8'd145; a_mant2 = 8'd27; a_mant3 = 8'd165;
b_mant0 = 8'd246; b_mant1 = 8'd154; b_mant2 = 8'd37; b_mant3 = 8'd14;
a_exp0 = 10'd628; a_exp1 = 10'd55; a_exp2 = 10'd421; a_exp3 = 10'd665;
b_exp0 = 10'd596; b_exp1 = 10'd961; b_exp2 = 10'd872; b_exp3 = 10'd462;
a_sign0 = 4'd6; a_sign1 = 4'd10; a_sign2 = 4'd4; a_sign3 = 4'd14;
b_sign0 = 4'd12; b_sign1 = 4'd8; b_sign2 = 4'd13; b_sign3 = 4'd3;
@(posedge clk_i);
a_mant0 = 8'd148; a_mant1 = 8'd254; a_mant2 = 8'd138; a_mant3 = 8'd13;
b_mant0 = 8'd156; b_mant1 = 8'd56; b_mant2 = 8'd36; b_mant3 = 8'd205;
a_exp0 = 10'd693; a_exp1 = 10'd22; a_exp2 = 10'd550; a_exp3 = 10'd296;
b_exp0 = 10'd571; b_exp1 = 10'd537; b_exp2 = 10'd968; b_exp3 = 10'd725;
a_sign0 = 4'd10; a_sign1 = 4'd8; a_sign2 = 4'd14; a_sign3 = 4'd16;
b_sign0 = 4'd15; b_sign1 = 4'd12; b_sign2 = 4'd9; b_sign3 = 4'd16;
@(posedge clk_i);
a_mant0 = 8'd218; a_mant1 = 8'd148; a_mant2 = 8'd129; a_mant3 = 8'd130;
b_mant0 = 8'd225; b_mant1 = 8'd129; b_mant2 = 8'd174; b_mant3 = 8'd118;
a_exp0 = 10'd1022; a_exp1 = 10'd339; a_exp2 = 10'd878; a_exp3 = 10'd942;
b_exp0 = 10'd697; b_exp1 = 10'd83; b_exp2 = 10'd589; b_exp3 = 10'd772;
a_sign0 = 4'd10; a_sign1 = 4'd6; a_sign2 = 4'd3; a_sign3 = 4'd8;
b_sign0 = 4'd9; b_sign1 = 4'd3; b_sign2 = 4'd2; b_sign3 = 4'd10;
@(posedge clk_i);
a_mant0 = 8'd26; a_mant1 = 8'd234; a_mant2 = 8'd169; a_mant3 = 8'd71;
b_mant0 = 8'd253; b_mant1 = 8'd76; b_mant2 = 8'd228; b_mant3 = 8'd189;
a_exp0 = 10'd648; a_exp1 = 10'd153; a_exp2 = 10'd547; a_exp3 = 10'd242;
b_exp0 = 10'd378; b_exp1 = 10'd702; b_exp2 = 10'd948; b_exp3 = 10'd558;
a_sign0 = 4'd6; a_sign1 = 4'd13; a_sign2 = 4'd4; a_sign3 = 4'd4;
b_sign0 = 4'd7; b_sign1 = 4'd4; b_sign2 = 4'd13; b_sign3 = 4'd3;
@(posedge clk_i);
a_mant0 = 8'd139; a_mant1 = 8'd59; a_mant2 = 8'd164; a_mant3 = 8'd4;
b_mant0 = 8'd95; b_mant1 = 8'd170; b_mant2 = 8'd47; b_mant3 = 8'd176;
a_exp0 = 10'd691; a_exp1 = 10'd530; a_exp2 = 10'd646; a_exp3 = 10'd179;
b_exp0 = 10'd246; b_exp1 = 10'd912; b_exp2 = 10'd591; b_exp3 = 10'd588;
a_sign0 = 4'd3; a_sign1 = 4'd3; a_sign2 = 4'd11; a_sign3 = 4'd4;
b_sign0 = 4'd13; b_sign1 = 4'd1; b_sign2 = 4'd11; b_sign3 = 4'd4;
@(posedge clk_i);
a_mant0 = 8'd229; a_mant1 = 8'd234; a_mant2 = 8'd235; a_mant3 = 8'd238;
b_mant0 = 8'd211; b_mant1 = 8'd216; b_mant2 = 8'd132; b_mant3 = 8'd23;
a_exp0 = 10'd316; a_exp1 = 10'd763; a_exp2 = 10'd92; a_exp3 = 10'd122;
b_exp0 = 10'd631; b_exp1 = 10'd751; b_exp2 = 10'd944; b_exp3 = 10'd392;
a_sign0 = 4'd13; a_sign1 = 4'd9; a_sign2 = 4'd13; a_sign3 = 4'd13;
b_sign0 = 4'd2; b_sign1 = 4'd11; b_sign2 = 4'd9; b_sign3 = 4'd4;
@(posedge clk_i);
a_mant0 = 8'd104; a_mant1 = 8'd174; a_mant2 = 8'd112; a_mant3 = 8'd227;
b_mant0 = 8'd66; b_mant1 = 8'd245; b_mant2 = 8'd216; b_mant3 = 8'd241;
a_exp0 = 10'd1011; a_exp1 = 10'd992; a_exp2 = 10'd977; a_exp3 = 10'd564;
b_exp0 = 10'd131; b_exp1 = 10'd768; b_exp2 = 10'd62; b_exp3 = 10'd248;
a_sign0 = 4'd13; a_sign1 = 4'd16; a_sign2 = 4'd8; a_sign3 = 4'd9;
b_sign0 = 4'd10; b_sign1 = 4'd7; b_sign2 = 4'd0; b_sign3 = 4'd13;
@(posedge clk_i);
a_mant0 = 8'd171; a_mant1 = 8'd113; a_mant2 = 8'd87; a_mant3 = 8'd67;
b_mant0 = 8'd128; b_mant1 = 8'd127; b_mant2 = 8'd45; b_mant3 = 8'd144;
a_exp0 = 10'd64; a_exp1 = 10'd834; a_exp2 = 10'd387; a_exp3 = 10'd747;
b_exp0 = 10'd652; b_exp1 = 10'd245; b_exp2 = 10'd335; b_exp3 = 10'd207;
a_sign0 = 4'd4; a_sign1 = 4'd1; a_sign2 = 4'd6; a_sign3 = 4'd12;
b_sign0 = 4'd15; b_sign1 = 4'd4; b_sign2 = 4'd14; b_sign3 = 4'd10;
@(posedge clk_i);
shared_exps0 = 8'd114;
shared_exps1 = 8'd129;
a_mant0 = 8'd45; a_mant1 = 8'd240; a_mant2 = 8'd109; a_mant3 = 8'd140;
b_mant0 = 8'd148; b_mant1 = 8'd82; b_mant2 = 8'd69; b_mant3 = 8'd147;
a_exp0 = 10'd677; a_exp1 = 10'd981; a_exp2 = 10'd9; a_exp3 = 10'd373;
b_exp0 = 10'd897; b_exp1 = 10'd312; b_exp2 = 10'd496; b_exp3 = 10'd499;
a_sign0 = 4'd9; a_sign1 = 4'd11; a_sign2 = 4'd10; a_sign3 = 4'd2;
b_sign0 = 4'd16; b_sign1 = 4'd10; b_sign2 = 4'd1; b_sign3 = 4'd12;
@(posedge clk_i);
a_mant0 = 8'd23; a_mant1 = 8'd193; a_mant2 = 8'd181; a_mant3 = 8'd243;
b_mant0 = 8'd218; b_mant1 = 8'd6; b_mant2 = 8'd169; b_mant3 = 8'd224;
a_exp0 = 10'd797; a_exp1 = 10'd594; a_exp2 = 10'd394; a_exp3 = 10'd661;
b_exp0 = 10'd997; b_exp1 = 10'd60; b_exp2 = 10'd225; b_exp3 = 10'd604;
a_sign0 = 4'd4; a_sign1 = 4'd9; a_sign2 = 4'd9; a_sign3 = 4'd5;
b_sign0 = 4'd9; b_sign1 = 4'd13; b_sign2 = 4'd0; b_sign3 = 4'd11;
@(posedge clk_i);
a_mant0 = 8'd176; a_mant1 = 8'd177; a_mant2 = 8'd226; a_mant3 = 8'd113;
b_mant0 = 8'd162; b_mant1 = 8'd177; b_mant2 = 8'd198; b_mant3 = 8'd39;
a_exp0 = 10'd50; a_exp1 = 10'd127; a_exp2 = 10'd284; a_exp3 = 10'd759;
b_exp0 = 10'd565; b_exp1 = 10'd749; b_exp2 = 10'd260; b_exp3 = 10'd356;
a_sign0 = 4'd9; a_sign1 = 4'd7; a_sign2 = 4'd7; a_sign3 = 4'd7;
b_sign0 = 4'd14; b_sign1 = 4'd14; b_sign2 = 4'd15; b_sign3 = 4'd9;
@(posedge clk_i);
a_mant0 = 8'd75; a_mant1 = 8'd84; a_mant2 = 8'd201; a_mant3 = 8'd33;
b_mant0 = 8'd128; b_mant1 = 8'd190; b_mant2 = 8'd78; b_mant3 = 8'd178;
a_exp0 = 10'd224; a_exp1 = 10'd936; a_exp2 = 10'd166; a_exp3 = 10'd68;
b_exp0 = 10'd166; b_exp1 = 10'd127; b_exp2 = 10'd248; b_exp3 = 10'd238;
a_sign0 = 4'd4; a_sign1 = 4'd11; a_sign2 = 4'd0; a_sign3 = 4'd4;
b_sign0 = 4'd14; b_sign1 = 4'd6; b_sign2 = 4'd1; b_sign3 = 4'd11;
@(posedge clk_i);
a_mant0 = 8'd117; a_mant1 = 8'd79; a_mant2 = 8'd35; a_mant3 = 8'd73;
b_mant0 = 8'd198; b_mant1 = 8'd139; b_mant2 = 8'd132; b_mant3 = 8'd29;
a_exp0 = 10'd741; a_exp1 = 10'd846; a_exp2 = 10'd326; a_exp3 = 10'd153;
b_exp0 = 10'd816; b_exp1 = 10'd81; b_exp2 = 10'd131; b_exp3 = 10'd26;
a_sign0 = 4'd3; a_sign1 = 4'd11; a_sign2 = 4'd0; a_sign3 = 4'd1;
b_sign0 = 4'd12; b_sign1 = 4'd1; b_sign2 = 4'd16; b_sign3 = 4'd5;
@(posedge clk_i);
a_mant0 = 8'd148; a_mant1 = 8'd217; a_mant2 = 8'd209; a_mant3 = 8'd141;
b_mant0 = 8'd149; b_mant1 = 8'd99; b_mant2 = 8'd77; b_mant3 = 8'd168;
a_exp0 = 10'd872; a_exp1 = 10'd103; a_exp2 = 10'd706; a_exp3 = 10'd648;
b_exp0 = 10'd140; b_exp1 = 10'd439; b_exp2 = 10'd90; b_exp3 = 10'd644;
a_sign0 = 4'd15; a_sign1 = 4'd11; a_sign2 = 4'd10; a_sign3 = 4'd8;
b_sign0 = 4'd9; b_sign1 = 4'd11; b_sign2 = 4'd6; b_sign3 = 4'd0;
@(posedge clk_i);
a_mant0 = 8'd59; a_mant1 = 8'd20; a_mant2 = 8'd121; a_mant3 = 8'd195;
b_mant0 = 8'd118; b_mant1 = 8'd24; b_mant2 = 8'd124; b_mant3 = 8'd161;
a_exp0 = 10'd675; a_exp1 = 10'd863; a_exp2 = 10'd868; a_exp3 = 10'd591;
b_exp0 = 10'd891; b_exp1 = 10'd98; b_exp2 = 10'd957; b_exp3 = 10'd859;
a_sign0 = 4'd10; a_sign1 = 4'd6; a_sign2 = 4'd8; a_sign3 = 4'd8;
b_sign0 = 4'd4; b_sign1 = 4'd6; b_sign2 = 4'd12; b_sign3 = 4'd14;
@(posedge clk_i);
a_mant0 = 8'd160; a_mant1 = 8'd134; a_mant2 = 8'd144; a_mant3 = 8'd90;
b_mant0 = 8'd89; b_mant1 = 8'd231; b_mant2 = 8'd254; b_mant3 = 8'd15;
a_exp0 = 10'd624; a_exp1 = 10'd128; a_exp2 = 10'd454; a_exp3 = 10'd441;
b_exp0 = 10'd20; b_exp1 = 10'd138; b_exp2 = 10'd345; b_exp3 = 10'd911;
a_sign0 = 4'd14; a_sign1 = 4'd10; a_sign2 = 4'd1; a_sign3 = 4'd12;
b_sign0 = 4'd11; b_sign1 = 4'd1; b_sign2 = 4'd0; b_sign3 = 4'd10;
@(posedge clk_i);
shared_exps0 = 8'd134;
shared_exps1 = 8'd116;
a_mant0 = 8'd102; a_mant1 = 8'd38; a_mant2 = 8'd245; a_mant3 = 8'd174;
b_mant0 = 8'd82; b_mant1 = 8'd183; b_mant2 = 8'd89; b_mant3 = 8'd178;
a_exp0 = 10'd868; a_exp1 = 10'd734; a_exp2 = 10'd218; a_exp3 = 10'd798;
b_exp0 = 10'd584; b_exp1 = 10'd754; b_exp2 = 10'd279; b_exp3 = 10'd206;
a_sign0 = 4'd8; a_sign1 = 4'd13; a_sign2 = 4'd12; a_sign3 = 4'd0;
b_sign0 = 4'd9; b_sign1 = 4'd16; b_sign2 = 4'd2; b_sign3 = 4'd1;
@(posedge clk_i);
a_mant0 = 8'd190; a_mant1 = 8'd107; a_mant2 = 8'd210; a_mant3 = 8'd194;
b_mant0 = 8'd13; b_mant1 = 8'd211; b_mant2 = 8'd250; b_mant3 = 8'd96;
a_exp0 = 10'd656; a_exp1 = 10'd989; a_exp2 = 10'd248; a_exp3 = 10'd817;
b_exp0 = 10'd9; b_exp1 = 10'd156; b_exp2 = 10'd426; b_exp3 = 10'd844;
a_sign0 = 4'd1; a_sign1 = 4'd10; a_sign2 = 4'd3; a_sign3 = 4'd11;
b_sign0 = 4'd2; b_sign1 = 4'd2; b_sign2 = 4'd5; b_sign3 = 4'd5;
@(posedge clk_i);
a_mant0 = 8'd204; a_mant1 = 8'd56; a_mant2 = 8'd153; a_mant3 = 8'd248;
b_mant0 = 8'd249; b_mant1 = 8'd202; b_mant2 = 8'd98; b_mant3 = 8'd88;
a_exp0 = 10'd581; a_exp1 = 10'd818; a_exp2 = 10'd801; a_exp3 = 10'd23;
b_exp0 = 10'd911; b_exp1 = 10'd812; b_exp2 = 10'd537; b_exp3 = 10'd205;
a_sign0 = 4'd9; a_sign1 = 4'd3; a_sign2 = 4'd11; a_sign3 = 4'd11;
b_sign0 = 4'd15; b_sign1 = 4'd3; b_sign2 = 4'd2; b_sign3 = 4'd7;
@(posedge clk_i);
a_mant0 = 8'd61; a_mant1 = 8'd92; a_mant2 = 8'd25; a_mant3 = 8'd140;
b_mant0 = 8'd141; b_mant1 = 8'd197; b_mant2 = 8'd36; b_mant3 = 8'd52;
a_exp0 = 10'd818; a_exp1 = 10'd322; a_exp2 = 10'd459; a_exp3 = 10'd796;
b_exp0 = 10'd60; b_exp1 = 10'd928; b_exp2 = 10'd862; b_exp3 = 10'd1001;
a_sign0 = 4'd14; a_sign1 = 4'd4; a_sign2 = 4'd5; a_sign3 = 4'd5;
b_sign0 = 4'd9; b_sign1 = 4'd15; b_sign2 = 4'd0; b_sign3 = 4'd2;
@(posedge clk_i);
a_mant0 = 8'd198; a_mant1 = 8'd55; a_mant2 = 8'd63; a_mant3 = 8'd104;
b_mant0 = 8'd179; b_mant1 = 8'd191; b_mant2 = 8'd82; b_mant3 = 8'd54;
a_exp0 = 10'd722; a_exp1 = 10'd788; a_exp2 = 10'd306; a_exp3 = 10'd419;
b_exp0 = 10'd643; b_exp1 = 10'd653; b_exp2 = 10'd243; b_exp3 = 10'd892;
a_sign0 = 4'd8; a_sign1 = 4'd1; a_sign2 = 4'd13; a_sign3 = 4'd3;
b_sign0 = 4'd10; b_sign1 = 4'd10; b_sign2 = 4'd4; b_sign3 = 4'd13;
@(posedge clk_i);
a_mant0 = 8'd27; a_mant1 = 8'd118; a_mant2 = 8'd111; a_mant3 = 8'd113;
b_mant0 = 8'd73; b_mant1 = 8'd180; b_mant2 = 8'd6; b_mant3 = 8'd117;
a_exp0 = 10'd939; a_exp1 = 10'd885; a_exp2 = 10'd13; a_exp3 = 10'd726;
b_exp0 = 10'd154; b_exp1 = 10'd580; b_exp2 = 10'd43; b_exp3 = 10'd822;
a_sign0 = 4'd4; a_sign1 = 4'd13; a_sign2 = 4'd4; a_sign3 = 4'd14;
b_sign0 = 4'd8; b_sign1 = 4'd12; b_sign2 = 4'd10; b_sign3 = 4'd1;
@(posedge clk_i);
a_mant0 = 8'd211; a_mant1 = 8'd150; a_mant2 = 8'd10; a_mant3 = 8'd36;
b_mant0 = 8'd230; b_mant1 = 8'd34; b_mant2 = 8'd30; b_mant3 = 8'd67;
a_exp0 = 10'd146; a_exp1 = 10'd538; a_exp2 = 10'd800; a_exp3 = 10'd163;
b_exp0 = 10'd612; b_exp1 = 10'd809; b_exp2 = 10'd652; b_exp3 = 10'd831;
a_sign0 = 4'd4; a_sign1 = 4'd15; a_sign2 = 4'd2; a_sign3 = 4'd11;
b_sign0 = 4'd4; b_sign1 = 4'd4; b_sign2 = 4'd5; b_sign3 = 4'd5;
@(posedge clk_i);
a_mant0 = 8'd48; a_mant1 = 8'd94; a_mant2 = 8'd240; a_mant3 = 8'd30;
b_mant0 = 8'd61; b_mant1 = 8'd64; b_mant2 = 8'd7; b_mant3 = 8'd203;
a_exp0 = 10'd1009; a_exp1 = 10'd494; a_exp2 = 10'd82; a_exp3 = 10'd1023;
b_exp0 = 10'd32; b_exp1 = 10'd823; b_exp2 = 10'd903; b_exp3 = 10'd807;
a_sign0 = 4'd15; a_sign1 = 4'd4; a_sign2 = 4'd7; a_sign3 = 4'd15;
b_sign0 = 4'd2; b_sign1 = 4'd11; b_sign2 = 4'd1; b_sign3 = 4'd16;
@(posedge clk_i);
shared_exps0 = 8'd128;
shared_exps1 = 8'd139;
rstn = 0;
@(posedge clk_i);
rstn = 1;
a_mant0 = 8'd179; a_mant1 = 8'd112; a_mant2 = 8'd79; a_mant3 = 8'd255;
b_mant0 = 8'd209; b_mant1 = 8'd156; b_mant2 = 8'd38; b_mant3 = 8'd9;
a_exp0 = 10'd464; a_exp1 = 10'd371; a_exp2 = 10'd403; a_exp3 = 10'd857;
b_exp0 = 10'd76; b_exp1 = 10'd585; b_exp2 = 10'd333; b_exp3 = 10'd463;
a_sign0 = 4'd9; a_sign1 = 4'd12; a_sign2 = 4'd10; a_sign3 = 4'd15;
b_sign0 = 4'd6; b_sign1 = 4'd9; b_sign2 = 4'd14; b_sign3 = 4'd1;
@(posedge clk_i);
a_mant0 = 8'd183; a_mant1 = 8'd63; a_mant2 = 8'd222; a_mant3 = 8'd147;
b_mant0 = 8'd13; b_mant1 = 8'd206; b_mant2 = 8'd160; b_mant3 = 8'd207;
a_exp0 = 10'd325; a_exp1 = 10'd621; a_exp2 = 10'd876; a_exp3 = 10'd462;
b_exp0 = 10'd300; b_exp1 = 10'd948; b_exp2 = 10'd977; b_exp3 = 10'd960;
a_sign0 = 4'd15; a_sign1 = 4'd0; a_sign2 = 4'd8; a_sign3 = 4'd0;
b_sign0 = 4'd6; b_sign1 = 4'd3; b_sign2 = 4'd15; b_sign3 = 4'd8;
@(posedge clk_i);
a_mant0 = 8'd24; a_mant1 = 8'd162; a_mant2 = 8'd16; a_mant3 = 8'd148;
b_mant0 = 8'd74; b_mant1 = 8'd134; b_mant2 = 8'd53; b_mant3 = 8'd31;
a_exp0 = 10'd891; a_exp1 = 10'd915; a_exp2 = 10'd879; a_exp3 = 10'd356;
b_exp0 = 10'd820; b_exp1 = 10'd354; b_exp2 = 10'd542; b_exp3 = 10'd2;
a_sign0 = 4'd16; a_sign1 = 4'd4; a_sign2 = 4'd15; a_sign3 = 4'd8;
b_sign0 = 4'd6; b_sign1 = 4'd16; b_sign2 = 4'd2; b_sign3 = 4'd13;
@(posedge clk_i);
a_mant0 = 8'd174; a_mant1 = 8'd157; a_mant2 = 8'd75; a_mant3 = 8'd187;
b_mant0 = 8'd169; b_mant1 = 8'd204; b_mant2 = 8'd226; b_mant3 = 8'd74;
a_exp0 = 10'd917; a_exp1 = 10'd869; a_exp2 = 10'd679; a_exp3 = 10'd257;
b_exp0 = 10'd451; b_exp1 = 10'd320; b_exp2 = 10'd965; b_exp3 = 10'd541;
a_sign0 = 4'd10; a_sign1 = 4'd3; a_sign2 = 4'd1; a_sign3 = 4'd4;
b_sign0 = 4'd8; b_sign1 = 4'd16; b_sign2 = 4'd8; b_sign3 = 4'd9;
@(posedge clk_i);
a_mant0 = 8'd71; a_mant1 = 8'd42; a_mant2 = 8'd20; a_mant3 = 8'd8;
b_mant0 = 8'd173; b_mant1 = 8'd212; b_mant2 = 8'd136; b_mant3 = 8'd62;
a_exp0 = 10'd720; a_exp1 = 10'd806; a_exp2 = 10'd823; a_exp3 = 10'd440;
b_exp0 = 10'd233; b_exp1 = 10'd198; b_exp2 = 10'd747; b_exp3 = 10'd293;
a_sign0 = 4'd5; a_sign1 = 4'd12; a_sign2 = 4'd6; a_sign3 = 4'd1;
b_sign0 = 4'd10; b_sign1 = 4'd15; b_sign2 = 4'd14; b_sign3 = 4'd0;
@(posedge clk_i);
a_mant0 = 8'd131; a_mant1 = 8'd1; a_mant2 = 8'd61; a_mant3 = 8'd205;
b_mant0 = 8'd149; b_mant1 = 8'd191; b_mant2 = 8'd99; b_mant3 = 8'd154;
a_exp0 = 10'd890; a_exp1 = 10'd995; a_exp2 = 10'd161; a_exp3 = 10'd195;
b_exp0 = 10'd662; b_exp1 = 10'd166; b_exp2 = 10'd261; b_exp3 = 10'd248;
a_sign0 = 4'd16; a_sign1 = 4'd10; a_sign2 = 4'd14; a_sign3 = 4'd12;
b_sign0 = 4'd12; b_sign1 = 4'd7; b_sign2 = 4'd12; b_sign3 = 4'd16;
@(posedge clk_i);
a_mant0 = 8'd133; a_mant1 = 8'd144; a_mant2 = 8'd154; a_mant3 = 8'd75;
b_mant0 = 8'd16; b_mant1 = 8'd190; b_mant2 = 8'd195; b_mant3 = 8'd13;
a_exp0 = 10'd322; a_exp1 = 10'd293; a_exp2 = 10'd230; a_exp3 = 10'd596;
b_exp0 = 10'd356; b_exp1 = 10'd393; b_exp2 = 10'd420; b_exp3 = 10'd518;
a_sign0 = 4'd13; a_sign1 = 4'd9; a_sign2 = 4'd13; a_sign3 = 4'd9;
b_sign0 = 4'd4; b_sign1 = 4'd9; b_sign2 = 4'd3; b_sign3 = 4'd1;
@(posedge clk_i);
shared_exps0 = 8'd153;
shared_exps1 = 8'd118;
a_mant0 = 8'd154; a_mant1 = 8'd24; a_mant2 = 8'd112; a_mant3 = 8'd221;
b_mant0 = 8'd47; b_mant1 = 8'd244; b_mant2 = 8'd191; b_mant3 = 8'd234;
a_exp0 = 10'd517; a_exp1 = 10'd395; a_exp2 = 10'd55; a_exp3 = 10'd671;
b_exp0 = 10'd972; b_exp1 = 10'd256; b_exp2 = 10'd376; b_exp3 = 10'd773;
a_sign0 = 4'd1; a_sign1 = 4'd14; a_sign2 = 4'd10; a_sign3 = 4'd11;
b_sign0 = 4'd0; b_sign1 = 4'd5; b_sign2 = 4'd3; b_sign3 = 4'd14;
@(posedge clk_i);
a_mant0 = 8'd220; a_mant1 = 8'd103; a_mant2 = 8'd48; a_mant3 = 8'd198;
b_mant0 = 8'd214; b_mant1 = 8'd18; b_mant2 = 8'd7; b_mant3 = 8'd5;
a_exp0 = 10'd829; a_exp1 = 10'd683; a_exp2 = 10'd719; a_exp3 = 10'd199;
b_exp0 = 10'd110; b_exp1 = 10'd270; b_exp2 = 10'd725; b_exp3 = 10'd550;
a_sign0 = 4'd7; a_sign1 = 4'd10; a_sign2 = 4'd12; a_sign3 = 4'd8;
b_sign0 = 4'd10; b_sign1 = 4'd0; b_sign2 = 4'd4; b_sign3 = 4'd4;
@(posedge clk_i);
a_mant0 = 8'd234; a_mant1 = 8'd111; a_mant2 = 8'd243; a_mant3 = 8'd57;
b_mant0 = 8'd179; b_mant1 = 8'd61; b_mant2 = 8'd168; b_mant3 = 8'd12;
a_exp0 = 10'd409; a_exp1 = 10'd1000; a_exp2 = 10'd549; a_exp3 = 10'd1016;
b_exp0 = 10'd483; b_exp1 = 10'd410; b_exp2 = 10'd348; b_exp3 = 10'd587;
a_sign0 = 4'd9; a_sign1 = 4'd15; a_sign2 = 4'd1; a_sign3 = 4'd3;
b_sign0 = 4'd12; b_sign1 = 4'd3; b_sign2 = 4'd4; b_sign3 = 4'd3;
@(posedge clk_i);
a_mant0 = 8'd58; a_mant1 = 8'd44; a_mant2 = 8'd229; a_mant3 = 8'd176;
b_mant0 = 8'd93; b_mant1 = 8'd153; b_mant2 = 8'd16; b_mant3 = 8'd83;
a_exp0 = 10'd951; a_exp1 = 10'd659; a_exp2 = 10'd816; a_exp3 = 10'd931;
b_exp0 = 10'd311; b_exp1 = 10'd207; b_exp2 = 10'd671; b_exp3 = 10'd444;
a_sign0 = 4'd12; a_sign1 = 4'd14; a_sign2 = 4'd0; a_sign3 = 4'd3;
b_sign0 = 4'd16; b_sign1 = 4'd10; b_sign2 = 4'd14; b_sign3 = 4'd13;
@(posedge clk_i);
a_mant0 = 8'd36; a_mant1 = 8'd113; a_mant2 = 8'd108; a_mant3 = 8'd61;
b_mant0 = 8'd141; b_mant1 = 8'd74; b_mant2 = 8'd172; b_mant3 = 8'd15;
a_exp0 = 10'd191; a_exp1 = 10'd653; a_exp2 = 10'd373; a_exp3 = 10'd997;
b_exp0 = 10'd76; b_exp1 = 10'd122; b_exp2 = 10'd694; b_exp3 = 10'd833;
a_sign0 = 4'd4; a_sign1 = 4'd11; a_sign2 = 4'd13; a_sign3 = 4'd15;
b_sign0 = 4'd11; b_sign1 = 4'd7; b_sign2 = 4'd13; b_sign3 = 4'd6;
@(posedge clk_i);
a_mant0 = 8'd61; a_mant1 = 8'd219; a_mant2 = 8'd238; a_mant3 = 8'd101;
b_mant0 = 8'd124; b_mant1 = 8'd131; b_mant2 = 8'd154; b_mant3 = 8'd186;
a_exp0 = 10'd64; a_exp1 = 10'd476; a_exp2 = 10'd862; a_exp3 = 10'd142;
b_exp0 = 10'd786; b_exp1 = 10'd758; b_exp2 = 10'd222; b_exp3 = 10'd524;
a_sign0 = 4'd4; a_sign1 = 4'd13; a_sign2 = 4'd0; a_sign3 = 4'd10;
b_sign0 = 4'd2; b_sign1 = 4'd3; b_sign2 = 4'd9; b_sign3 = 4'd16;
@(posedge clk_i);
a_mant0 = 8'd215; a_mant1 = 8'd90; a_mant2 = 8'd139; a_mant3 = 8'd183;
b_mant0 = 8'd186; b_mant1 = 8'd140; b_mant2 = 8'd38; b_mant3 = 8'd2;
a_exp0 = 10'd905; a_exp1 = 10'd75; a_exp2 = 10'd904; a_exp3 = 10'd176;
b_exp0 = 10'd936; b_exp1 = 10'd296; b_exp2 = 10'd677; b_exp3 = 10'd346;
a_sign0 = 4'd5; a_sign1 = 4'd0; a_sign2 = 4'd15; a_sign3 = 4'd7;
b_sign0 = 4'd3; b_sign1 = 4'd15; b_sign2 = 4'd0; b_sign3 = 4'd8;
@(posedge clk_i);
a_mant0 = 8'd35; a_mant1 = 8'd232; a_mant2 = 8'd33; a_mant3 = 8'd169;
b_mant0 = 8'd31; b_mant1 = 8'd53; b_mant2 = 8'd16; b_mant3 = 8'd47;
a_exp0 = 10'd271; a_exp1 = 10'd962; a_exp2 = 10'd217; a_exp3 = 10'd477;
b_exp0 = 10'd164; b_exp1 = 10'd749; b_exp2 = 10'd809; b_exp3 = 10'd564;
a_sign0 = 4'd3; a_sign1 = 4'd1; a_sign2 = 4'd14; a_sign3 = 4'd4;
b_sign0 = 4'd15; b_sign1 = 4'd10; b_sign2 = 4'd8; b_sign3 = 4'd16;
@(posedge clk_i);
shared_exps0 = 8'd147;
shared_exps1 = 8'd125;
a_mant0 = 8'd62; a_mant1 = 8'd108; a_mant2 = 8'd153; a_mant3 = 8'd242;
b_mant0 = 8'd12; b_mant1 = 8'd112; b_mant2 = 8'd47; b_mant3 = 8'd93;
a_exp0 = 10'd577; a_exp1 = 10'd103; a_exp2 = 10'd989; a_exp3 = 10'd864;
b_exp0 = 10'd339; b_exp1 = 10'd567; b_exp2 = 10'd1018; b_exp3 = 10'd187;
a_sign0 = 4'd1; a_sign1 = 4'd8; a_sign2 = 4'd4; a_sign3 = 4'd0;
b_sign0 = 4'd3; b_sign1 = 4'd12; b_sign2 = 4'd9; b_sign3 = 4'd16;
@(posedge clk_i);
a_mant0 = 8'd232; a_mant1 = 8'd174; a_mant2 = 8'd93; a_mant3 = 8'd12;
b_mant0 = 8'd30; b_mant1 = 8'd188; b_mant2 = 8'd185; b_mant3 = 8'd69;
a_exp0 = 10'd797; a_exp1 = 10'd818; a_exp2 = 10'd119; a_exp3 = 10'd670;
b_exp0 = 10'd414; b_exp1 = 10'd1023; b_exp2 = 10'd581; b_exp3 = 10'd535;
a_sign0 = 4'd10; a_sign1 = 4'd6; a_sign2 = 4'd9; a_sign3 = 4'd7;
b_sign0 = 4'd13; b_sign1 = 4'd10; b_sign2 = 4'd6; b_sign3 = 4'd5;
@(posedge clk_i);
a_mant0 = 8'd205; a_mant1 = 8'd253; a_mant2 = 8'd37; a_mant3 = 8'd11;
b_mant0 = 8'd32; b_mant1 = 8'd140; b_mant2 = 8'd58; b_mant3 = 8'd90;
a_exp0 = 10'd938; a_exp1 = 10'd96; a_exp2 = 10'd887; a_exp3 = 10'd29;
b_exp0 = 10'd508; b_exp1 = 10'd320; b_exp2 = 10'd18; b_exp3 = 10'd228;
a_sign0 = 4'd10; a_sign1 = 4'd15; a_sign2 = 4'd15; a_sign3 = 4'd6;
b_sign0 = 4'd0; b_sign1 = 4'd16; b_sign2 = 4'd0; b_sign3 = 4'd2;
@(posedge clk_i);
a_mant0 = 8'd206; a_mant1 = 8'd233; a_mant2 = 8'd42; a_mant3 = 8'd127;
b_mant0 = 8'd225; b_mant1 = 8'd170; b_mant2 = 8'd125; b_mant3 = 8'd141;
a_exp0 = 10'd282; a_exp1 = 10'd648; a_exp2 = 10'd547; a_exp3 = 10'd773;
b_exp0 = 10'd301; b_exp1 = 10'd403; b_exp2 = 10'd966; b_exp3 = 10'd59;
a_sign0 = 4'd15; a_sign1 = 4'd7; a_sign2 = 4'd0; a_sign3 = 4'd8;
b_sign0 = 4'd13; b_sign1 = 4'd7; b_sign2 = 4'd8; b_sign3 = 4'd1;
@(posedge clk_i);
a_mant0 = 8'd86; a_mant1 = 8'd205; a_mant2 = 8'd86; a_mant3 = 8'd245;
b_mant0 = 8'd254; b_mant1 = 8'd0; b_mant2 = 8'd32; b_mant3 = 8'd163;
a_exp0 = 10'd549; a_exp1 = 10'd522; a_exp2 = 10'd672; a_exp3 = 10'd589;
b_exp0 = 10'd351; b_exp1 = 10'd465; b_exp2 = 10'd69; b_exp3 = 10'd923;
a_sign0 = 4'd13; a_sign1 = 4'd8; a_sign2 = 4'd4; a_sign3 = 4'd9;
b_sign0 = 4'd0; b_sign1 = 4'd13; b_sign2 = 4'd8; b_sign3 = 4'd15;
@(posedge clk_i);
a_mant0 = 8'd192; a_mant1 = 8'd22; a_mant2 = 8'd164; a_mant3 = 8'd157;
b_mant0 = 8'd80; b_mant1 = 8'd46; b_mant2 = 8'd103; b_mant3 = 8'd132;
a_exp0 = 10'd513; a_exp1 = 10'd481; a_exp2 = 10'd889; a_exp3 = 10'd207;
b_exp0 = 10'd412; b_exp1 = 10'd504; b_exp2 = 10'd71; b_exp3 = 10'd135;
a_sign0 = 4'd1; a_sign1 = 4'd3; a_sign2 = 4'd7; a_sign3 = 4'd2;
b_sign0 = 4'd8; b_sign1 = 4'd8; b_sign2 = 4'd13; b_sign3 = 4'd13;
@(posedge clk_i);
a_mant0 = 8'd250; a_mant1 = 8'd108; a_mant2 = 8'd163; a_mant3 = 8'd95;
b_mant0 = 8'd230; b_mant1 = 8'd205; b_mant2 = 8'd173; b_mant3 = 8'd85;
a_exp0 = 10'd852; a_exp1 = 10'd561; a_exp2 = 10'd711; a_exp3 = 10'd714;
b_exp0 = 10'd569; b_exp1 = 10'd208; b_exp2 = 10'd472; b_exp3 = 10'd530;
a_sign0 = 4'd11; a_sign1 = 4'd15; a_sign2 = 4'd7; a_sign3 = 4'd3;
b_sign0 = 4'd13; b_sign1 = 4'd3; b_sign2 = 4'd11; b_sign3 = 4'd1;
@(posedge clk_i);
a_mant0 = 8'd124; a_mant1 = 8'd8; a_mant2 = 8'd34; a_mant3 = 8'd93;
b_mant0 = 8'd220; b_mant1 = 8'd66; b_mant2 = 8'd149; b_mant3 = 8'd137;
a_exp0 = 10'd312; a_exp1 = 10'd860; a_exp2 = 10'd324; a_exp3 = 10'd207;
b_exp0 = 10'd167; b_exp1 = 10'd72; b_exp2 = 10'd134; b_exp3 = 10'd231;
a_sign0 = 4'd3; a_sign1 = 4'd1; a_sign2 = 4'd16; a_sign3 = 4'd7;
b_sign0 = 4'd8; b_sign1 = 4'd11; b_sign2 = 4'd9; b_sign3 = 4'd2;
@(posedge clk_i);
shared_exps0 = 8'd114;
shared_exps1 = 8'd157;
a_mant0 = 8'd170; a_mant1 = 8'd141; a_mant2 = 8'd183; a_mant3 = 8'd102;
b_mant0 = 8'd11; b_mant1 = 8'd88; b_mant2 = 8'd128; b_mant3 = 8'd188;
a_exp0 = 10'd512; a_exp1 = 10'd670; a_exp2 = 10'd335; a_exp3 = 10'd982;
b_exp0 = 10'd977; b_exp1 = 10'd452; b_exp2 = 10'd593; b_exp3 = 10'd388;
a_sign0 = 4'd10; a_sign1 = 4'd15; a_sign2 = 4'd10; a_sign3 = 4'd6;
b_sign0 = 4'd13; b_sign1 = 4'd1; b_sign2 = 4'd6; b_sign3 = 4'd16;
@(posedge clk_i);
a_mant0 = 8'd40; a_mant1 = 8'd139; a_mant2 = 8'd239; a_mant3 = 8'd201;
b_mant0 = 8'd122; b_mant1 = 8'd236; b_mant2 = 8'd32; b_mant3 = 8'd193;
a_exp0 = 10'd742; a_exp1 = 10'd624; a_exp2 = 10'd873; a_exp3 = 10'd112;
b_exp0 = 10'd946; b_exp1 = 10'd140; b_exp2 = 10'd922; b_exp3 = 10'd589;
a_sign0 = 4'd3; a_sign1 = 4'd12; a_sign2 = 4'd11; a_sign3 = 4'd14;
b_sign0 = 4'd3; b_sign1 = 4'd0; b_sign2 = 4'd5; b_sign3 = 4'd1;
@(posedge clk_i);
a_mant0 = 8'd151; a_mant1 = 8'd68; a_mant2 = 8'd205; a_mant3 = 8'd107;
b_mant0 = 8'd84; b_mant1 = 8'd219; b_mant2 = 8'd180; b_mant3 = 8'd121;
a_exp0 = 10'd777; a_exp1 = 10'd116; a_exp2 = 10'd35; a_exp3 = 10'd579;
b_exp0 = 10'd741; b_exp1 = 10'd238; b_exp2 = 10'd121; b_exp3 = 10'd471;
a_sign0 = 4'd7; a_sign1 = 4'd0; a_sign2 = 4'd2; a_sign3 = 4'd6;
b_sign0 = 4'd16; b_sign1 = 4'd4; b_sign2 = 4'd0; b_sign3 = 4'd11;
@(posedge clk_i);
a_mant0 = 8'd29; a_mant1 = 8'd29; a_mant2 = 8'd29; a_mant3 = 8'd163;
b_mant0 = 8'd49; b_mant1 = 8'd219; b_mant2 = 8'd89; b_mant3 = 8'd130;
a_exp0 = 10'd566; a_exp1 = 10'd741; a_exp2 = 10'd105; a_exp3 = 10'd632;
b_exp0 = 10'd672; b_exp1 = 10'd779; b_exp2 = 10'd536; b_exp3 = 10'd388;
a_sign0 = 4'd5; a_sign1 = 4'd10; a_sign2 = 4'd6; a_sign3 = 4'd3;
b_sign0 = 4'd6; b_sign1 = 4'd8; b_sign2 = 4'd4; b_sign3 = 4'd13;
@(posedge clk_i);
a_mant0 = 8'd240; a_mant1 = 8'd206; a_mant2 = 8'd84; a_mant3 = 8'd250;
b_mant0 = 8'd174; b_mant1 = 8'd157; b_mant2 = 8'd44; b_mant3 = 8'd217;
a_exp0 = 10'd581; a_exp1 = 10'd229; a_exp2 = 10'd696; a_exp3 = 10'd926;
b_exp0 = 10'd161; b_exp1 = 10'd163; b_exp2 = 10'd487; b_exp3 = 10'd796;
a_sign0 = 4'd0; a_sign1 = 4'd9; a_sign2 = 4'd16; a_sign3 = 4'd10;
b_sign0 = 4'd10; b_sign1 = 4'd12; b_sign2 = 4'd7; b_sign3 = 4'd2;
@(posedge clk_i);
a_mant0 = 8'd5; a_mant1 = 8'd224; a_mant2 = 8'd196; a_mant3 = 8'd179;
b_mant0 = 8'd63; b_mant1 = 8'd114; b_mant2 = 8'd144; b_mant3 = 8'd170;
a_exp0 = 10'd779; a_exp1 = 10'd871; a_exp2 = 10'd304; a_exp3 = 10'd532;
b_exp0 = 10'd615; b_exp1 = 10'd480; b_exp2 = 10'd965; b_exp3 = 10'd806;
a_sign0 = 4'd4; a_sign1 = 4'd2; a_sign2 = 4'd11; a_sign3 = 4'd2;
b_sign0 = 4'd3; b_sign1 = 4'd1; b_sign2 = 4'd11; b_sign3 = 4'd7;
@(posedge clk_i);
a_mant0 = 8'd180; a_mant1 = 8'd101; a_mant2 = 8'd209; a_mant3 = 8'd243;
b_mant0 = 8'd126; b_mant1 = 8'd39; b_mant2 = 8'd74; b_mant3 = 8'd116;
a_exp0 = 10'd124; a_exp1 = 10'd116; a_exp2 = 10'd226; a_exp3 = 10'd1009;
b_exp0 = 10'd64; b_exp1 = 10'd714; b_exp2 = 10'd830; b_exp3 = 10'd670;
a_sign0 = 4'd15; a_sign1 = 4'd11; a_sign2 = 4'd9; a_sign3 = 4'd9;
b_sign0 = 4'd14; b_sign1 = 4'd14; b_sign2 = 4'd8; b_sign3 = 4'd16;
@(posedge clk_i);
a_mant0 = 8'd78; a_mant1 = 8'd254; a_mant2 = 8'd40; a_mant3 = 8'd115;
b_mant0 = 8'd168; b_mant1 = 8'd163; b_mant2 = 8'd16; b_mant3 = 8'd23;
a_exp0 = 10'd663; a_exp1 = 10'd477; a_exp2 = 10'd299; a_exp3 = 10'd201;
b_exp0 = 10'd813; b_exp1 = 10'd294; b_exp2 = 10'd392; b_exp3 = 10'd789;
a_sign0 = 4'd2; a_sign1 = 4'd0; a_sign2 = 4'd2; a_sign3 = 4'd5;
b_sign0 = 4'd16; b_sign1 = 4'd2; b_sign2 = 4'd11; b_sign3 = 4'd16;
@(posedge clk_i);
shared_exps0 = 8'd121;
shared_exps1 = 8'd127;
rstn = 0;
@(posedge clk_i);
rstn = 1;
a_mant0 = 8'd126; a_mant1 = 8'd102; a_mant2 = 8'd54; a_mant3 = 8'd122;
b_mant0 = 8'd76; b_mant1 = 8'd167; b_mant2 = 8'd254; b_mant3 = 8'd242;
a_exp0 = 10'd683; a_exp1 = 10'd61; a_exp2 = 10'd92; a_exp3 = 10'd141;
b_exp0 = 10'd391; b_exp1 = 10'd112; b_exp2 = 10'd175; b_exp3 = 10'd765;
a_sign0 = 4'd14; a_sign1 = 4'd6; a_sign2 = 4'd1; a_sign3 = 4'd16;
b_sign0 = 4'd2; b_sign1 = 4'd9; b_sign2 = 4'd6; b_sign3 = 4'd7;
@(posedge clk_i);
a_mant0 = 8'd240; a_mant1 = 8'd106; a_mant2 = 8'd238; a_mant3 = 8'd241;
b_mant0 = 8'd61; b_mant1 = 8'd197; b_mant2 = 8'd37; b_mant3 = 8'd101;
a_exp0 = 10'd403; a_exp1 = 10'd762; a_exp2 = 10'd415; a_exp3 = 10'd276;
b_exp0 = 10'd128; b_exp1 = 10'd676; b_exp2 = 10'd365; b_exp3 = 10'd477;
a_sign0 = 4'd0; a_sign1 = 4'd8; a_sign2 = 4'd8; a_sign3 = 4'd2;
b_sign0 = 4'd5; b_sign1 = 4'd7; b_sign2 = 4'd15; b_sign3 = 4'd13;
@(posedge clk_i);
a_mant0 = 8'd2; a_mant1 = 8'd181; a_mant2 = 8'd56; a_mant3 = 8'd62;
b_mant0 = 8'd241; b_mant1 = 8'd61; b_mant2 = 8'd150; b_mant3 = 8'd211;
a_exp0 = 10'd319; a_exp1 = 10'd25; a_exp2 = 10'd236; a_exp3 = 10'd29;
b_exp0 = 10'd719; b_exp1 = 10'd27; b_exp2 = 10'd16; b_exp3 = 10'd312;
a_sign0 = 4'd12; a_sign1 = 4'd4; a_sign2 = 4'd7; a_sign3 = 4'd3;
b_sign0 = 4'd1; b_sign1 = 4'd0; b_sign2 = 4'd5; b_sign3 = 4'd8;
@(posedge clk_i);
a_mant0 = 8'd172; a_mant1 = 8'd135; a_mant2 = 8'd157; a_mant3 = 8'd183;
b_mant0 = 8'd105; b_mant1 = 8'd213; b_mant2 = 8'd62; b_mant3 = 8'd52;
a_exp0 = 10'd554; a_exp1 = 10'd256; a_exp2 = 10'd174; a_exp3 = 10'd783;
b_exp0 = 10'd507; b_exp1 = 10'd520; b_exp2 = 10'd578; b_exp3 = 10'd446;
a_sign0 = 4'd10; a_sign1 = 4'd9; a_sign2 = 4'd14; a_sign3 = 4'd1;
b_sign0 = 4'd6; b_sign1 = 4'd3; b_sign2 = 4'd4; b_sign3 = 4'd16;
@(posedge clk_i);
a_mant0 = 8'd82; a_mant1 = 8'd241; a_mant2 = 8'd207; a_mant3 = 8'd101;
b_mant0 = 8'd231; b_mant1 = 8'd95; b_mant2 = 8'd148; b_mant3 = 8'd121;
a_exp0 = 10'd903; a_exp1 = 10'd796; a_exp2 = 10'd107; a_exp3 = 10'd736;
b_exp0 = 10'd116; b_exp1 = 10'd965; b_exp2 = 10'd722; b_exp3 = 10'd658;
a_sign0 = 4'd11; a_sign1 = 4'd3; a_sign2 = 4'd8; a_sign3 = 4'd5;
b_sign0 = 4'd16; b_sign1 = 4'd11; b_sign2 = 4'd14; b_sign3 = 4'd10;
@(posedge clk_i);
a_mant0 = 8'd39; a_mant1 = 8'd16; a_mant2 = 8'd91; a_mant3 = 8'd193;
b_mant0 = 8'd255; b_mant1 = 8'd219; b_mant2 = 8'd245; b_mant3 = 8'd81;
a_exp0 = 10'd304; a_exp1 = 10'd724; a_exp2 = 10'd348; a_exp3 = 10'd747;
b_exp0 = 10'd430; b_exp1 = 10'd714; b_exp2 = 10'd223; b_exp3 = 10'd554;
a_sign0 = 4'd3; a_sign1 = 4'd9; a_sign2 = 4'd12; a_sign3 = 4'd11;
b_sign0 = 4'd13; b_sign1 = 4'd7; b_sign2 = 4'd8; b_sign3 = 4'd12;
@(posedge clk_i);
a_mant0 = 8'd216; a_mant1 = 8'd154; a_mant2 = 8'd183; a_mant3 = 8'd85;
b_mant0 = 8'd221; b_mant1 = 8'd187; b_mant2 = 8'd148; b_mant3 = 8'd239;
a_exp0 = 10'd9; a_exp1 = 10'd928; a_exp2 = 10'd827; a_exp3 = 10'd590;
b_exp0 = 10'd333; b_exp1 = 10'd443; b_exp2 = 10'd596; b_exp3 = 10'd626;
a_sign0 = 4'd0; a_sign1 = 4'd12; a_sign2 = 4'd14; a_sign3 = 4'd5;
b_sign0 = 4'd4; b_sign1 = 4'd4; b_sign2 = 4'd0; b_sign3 = 4'd13;
@(posedge clk_i);
shared_exps0 = 8'd121;
shared_exps1 = 8'd139;
a_mant0 = 8'd124; a_mant1 = 8'd225; a_mant2 = 8'd15; a_mant3 = 8'd27;
b_mant0 = 8'd90; b_mant1 = 8'd191; b_mant2 = 8'd106; b_mant3 = 8'd146;
a_exp0 = 10'd981; a_exp1 = 10'd879; a_exp2 = 10'd103; a_exp3 = 10'd974;
b_exp0 = 10'd312; b_exp1 = 10'd114; b_exp2 = 10'd300; b_exp3 = 10'd553;
a_sign0 = 4'd8; a_sign1 = 4'd6; a_sign2 = 4'd6; a_sign3 = 4'd6;
b_sign0 = 4'd12; b_sign1 = 4'd14; b_sign2 = 4'd3; b_sign3 = 4'd0;
@(posedge clk_i);
a_mant0 = 8'd196; a_mant1 = 8'd49; a_mant2 = 8'd228; a_mant3 = 8'd150;
b_mant0 = 8'd105; b_mant1 = 8'd205; b_mant2 = 8'd105; b_mant3 = 8'd207;
a_exp0 = 10'd82; a_exp1 = 10'd396; a_exp2 = 10'd822; a_exp3 = 10'd0;
b_exp0 = 10'd72; b_exp1 = 10'd181; b_exp2 = 10'd173; b_exp3 = 10'd60;
a_sign0 = 4'd10; a_sign1 = 4'd13; a_sign2 = 4'd2; a_sign3 = 4'd9;
b_sign0 = 4'd7; b_sign1 = 4'd5; b_sign2 = 4'd7; b_sign3 = 4'd6;
@(posedge clk_i);
a_mant0 = 8'd99; a_mant1 = 8'd211; a_mant2 = 8'd158; a_mant3 = 8'd232;
b_mant0 = 8'd111; b_mant1 = 8'd57; b_mant2 = 8'd105; b_mant3 = 8'd82;
a_exp0 = 10'd622; a_exp1 = 10'd876; a_exp2 = 10'd940; a_exp3 = 10'd861;
b_exp0 = 10'd499; b_exp1 = 10'd762; b_exp2 = 10'd169; b_exp3 = 10'd451;
a_sign0 = 4'd13; a_sign1 = 4'd16; a_sign2 = 4'd0; a_sign3 = 4'd13;
b_sign0 = 4'd13; b_sign1 = 4'd15; b_sign2 = 4'd15; b_sign3 = 4'd10;
@(posedge clk_i);
a_mant0 = 8'd50; a_mant1 = 8'd103; a_mant2 = 8'd211; a_mant3 = 8'd25;
b_mant0 = 8'd68; b_mant1 = 8'd154; b_mant2 = 8'd248; b_mant3 = 8'd19;
a_exp0 = 10'd832; a_exp1 = 10'd83; a_exp2 = 10'd824; a_exp3 = 10'd451;
b_exp0 = 10'd541; b_exp1 = 10'd615; b_exp2 = 10'd727; b_exp3 = 10'd65;
a_sign0 = 4'd4; a_sign1 = 4'd7; a_sign2 = 4'd4; a_sign3 = 4'd3;
b_sign0 = 4'd13; b_sign1 = 4'd16; b_sign2 = 4'd10; b_sign3 = 4'd3;
@(posedge clk_i);
a_mant0 = 8'd98; a_mant1 = 8'd80; a_mant2 = 8'd88; a_mant3 = 8'd253;
b_mant0 = 8'd108; b_mant1 = 8'd45; b_mant2 = 8'd156; b_mant3 = 8'd210;
a_exp0 = 10'd727; a_exp1 = 10'd316; a_exp2 = 10'd306; a_exp3 = 10'd972;
b_exp0 = 10'd437; b_exp1 = 10'd480; b_exp2 = 10'd457; b_exp3 = 10'd82;
a_sign0 = 4'd0; a_sign1 = 4'd4; a_sign2 = 4'd6; a_sign3 = 4'd3;
b_sign0 = 4'd1; b_sign1 = 4'd2; b_sign2 = 4'd8; b_sign3 = 4'd10;
@(posedge clk_i);
a_mant0 = 8'd246; a_mant1 = 8'd17; a_mant2 = 8'd212; a_mant3 = 8'd120;
b_mant0 = 8'd138; b_mant1 = 8'd80; b_mant2 = 8'd85; b_mant3 = 8'd146;
a_exp0 = 10'd145; a_exp1 = 10'd917; a_exp2 = 10'd750; a_exp3 = 10'd605;
b_exp0 = 10'd622; b_exp1 = 10'd525; b_exp2 = 10'd815; b_exp3 = 10'd497;
a_sign0 = 4'd8; a_sign1 = 4'd1; a_sign2 = 4'd12; a_sign3 = 4'd13;
b_sign0 = 4'd6; b_sign1 = 4'd6; b_sign2 = 4'd6; b_sign3 = 4'd7;
@(posedge clk_i);
a_mant0 = 8'd252; a_mant1 = 8'd53; a_mant2 = 8'd199; a_mant3 = 8'd151;
b_mant0 = 8'd203; b_mant1 = 8'd46; b_mant2 = 8'd71; b_mant3 = 8'd243;
a_exp0 = 10'd159; a_exp1 = 10'd856; a_exp2 = 10'd612; a_exp3 = 10'd479;
b_exp0 = 10'd299; b_exp1 = 10'd79; b_exp2 = 10'd351; b_exp3 = 10'd951;
a_sign0 = 4'd0; a_sign1 = 4'd12; a_sign2 = 4'd9; a_sign3 = 4'd8;
b_sign0 = 4'd13; b_sign1 = 4'd0; b_sign2 = 4'd7; b_sign3 = 4'd9;
@(posedge clk_i);
a_mant0 = 8'd96; a_mant1 = 8'd231; a_mant2 = 8'd215; a_mant3 = 8'd128;
b_mant0 = 8'd2; b_mant1 = 8'd89; b_mant2 = 8'd23; b_mant3 = 8'd100;
a_exp0 = 10'd660; a_exp1 = 10'd821; a_exp2 = 10'd767; a_exp3 = 10'd366;
b_exp0 = 10'd64; b_exp1 = 10'd915; b_exp2 = 10'd311; b_exp3 = 10'd950;
a_sign0 = 4'd5; a_sign1 = 4'd8; a_sign2 = 4'd8; a_sign3 = 4'd5;
b_sign0 = 4'd15; b_sign1 = 4'd8; b_sign2 = 4'd14; b_sign3 = 4'd11;
@(posedge clk_i);
shared_exps0 = 8'd120;
shared_exps1 = 8'd134;
a_mant0 = 8'd196; a_mant1 = 8'd17; a_mant2 = 8'd182; a_mant3 = 8'd191;
b_mant0 = 8'd180; b_mant1 = 8'd149; b_mant2 = 8'd110; b_mant3 = 8'd206;
a_exp0 = 10'd928; a_exp1 = 10'd249; a_exp2 = 10'd901; a_exp3 = 10'd43;
b_exp0 = 10'd905; b_exp1 = 10'd199; b_exp2 = 10'd60; b_exp3 = 10'd37;
a_sign0 = 4'd7; a_sign1 = 4'd1; a_sign2 = 4'd11; a_sign3 = 4'd16;
b_sign0 = 4'd5; b_sign1 = 4'd7; b_sign2 = 4'd13; b_sign3 = 4'd12;
@(posedge clk_i);
a_mant0 = 8'd188; a_mant1 = 8'd60; a_mant2 = 8'd171; a_mant3 = 8'd217;
b_mant0 = 8'd66; b_mant1 = 8'd183; b_mant2 = 8'd72; b_mant3 = 8'd227;
a_exp0 = 10'd294; a_exp1 = 10'd776; a_exp2 = 10'd197; a_exp3 = 10'd490;
b_exp0 = 10'd62; b_exp1 = 10'd695; b_exp2 = 10'd616; b_exp3 = 10'd999;
a_sign0 = 4'd12; a_sign1 = 4'd12; a_sign2 = 4'd13; a_sign3 = 4'd9;
b_sign0 = 4'd2; b_sign1 = 4'd9; b_sign2 = 4'd15; b_sign3 = 4'd7;
@(posedge clk_i);
a_mant0 = 8'd232; a_mant1 = 8'd174; a_mant2 = 8'd122; a_mant3 = 8'd55;
b_mant0 = 8'd144; b_mant1 = 8'd193; b_mant2 = 8'd251; b_mant3 = 8'd131;
a_exp0 = 10'd637; a_exp1 = 10'd806; a_exp2 = 10'd520; a_exp3 = 10'd806;
b_exp0 = 10'd301; b_exp1 = 10'd26; b_exp2 = 10'd461; b_exp3 = 10'd447;
a_sign0 = 4'd1; a_sign1 = 4'd13; a_sign2 = 4'd6; a_sign3 = 4'd13;
b_sign0 = 4'd14; b_sign1 = 4'd13; b_sign2 = 4'd8; b_sign3 = 4'd0;
@(posedge clk_i);
a_mant0 = 8'd181; a_mant1 = 8'd123; a_mant2 = 8'd16; a_mant3 = 8'd120;
b_mant0 = 8'd173; b_mant1 = 8'd196; b_mant2 = 8'd13; b_mant3 = 8'd225;
a_exp0 = 10'd134; a_exp1 = 10'd147; a_exp2 = 10'd533; a_exp3 = 10'd579;
b_exp0 = 10'd720; b_exp1 = 10'd443; b_exp2 = 10'd713; b_exp3 = 10'd388;
a_sign0 = 4'd12; a_sign1 = 4'd11; a_sign2 = 4'd14; a_sign3 = 4'd13;
b_sign0 = 4'd0; b_sign1 = 4'd13; b_sign2 = 4'd10; b_sign3 = 4'd12;
@(posedge clk_i);
a_mant0 = 8'd79; a_mant1 = 8'd185; a_mant2 = 8'd49; a_mant3 = 8'd127;
b_mant0 = 8'd135; b_mant1 = 8'd73; b_mant2 = 8'd231; b_mant3 = 8'd113;
a_exp0 = 10'd697; a_exp1 = 10'd78; a_exp2 = 10'd958; a_exp3 = 10'd760;
b_exp0 = 10'd148; b_exp1 = 10'd827; b_exp2 = 10'd712; b_exp3 = 10'd448;
a_sign0 = 4'd10; a_sign1 = 4'd4; a_sign2 = 4'd5; a_sign3 = 4'd7;
b_sign0 = 4'd3; b_sign1 = 4'd14; b_sign2 = 4'd12; b_sign3 = 4'd15;
@(posedge clk_i);
a_mant0 = 8'd174; a_mant1 = 8'd27; a_mant2 = 8'd115; a_mant3 = 8'd152;
b_mant0 = 8'd227; b_mant1 = 8'd170; b_mant2 = 8'd125; b_mant3 = 8'd100;
a_exp0 = 10'd983; a_exp1 = 10'd902; a_exp2 = 10'd815; a_exp3 = 10'd949;
b_exp0 = 10'd49; b_exp1 = 10'd484; b_exp2 = 10'd641; b_exp3 = 10'd470;
a_sign0 = 4'd9; a_sign1 = 4'd13; a_sign2 = 4'd5; a_sign3 = 4'd15;
b_sign0 = 4'd15; b_sign1 = 4'd11; b_sign2 = 4'd6; b_sign3 = 4'd4;
@(posedge clk_i);
a_mant0 = 8'd7; a_mant1 = 8'd110; a_mant2 = 8'd153; a_mant3 = 8'd146;
b_mant0 = 8'd45; b_mant1 = 8'd48; b_mant2 = 8'd251; b_mant3 = 8'd9;
a_exp0 = 10'd863; a_exp1 = 10'd68; a_exp2 = 10'd291; a_exp3 = 10'd668;
b_exp0 = 10'd281; b_exp1 = 10'd214; b_exp2 = 10'd253; b_exp3 = 10'd896;
a_sign0 = 4'd14; a_sign1 = 4'd8; a_sign2 = 4'd4; a_sign3 = 4'd13;
b_sign0 = 4'd2; b_sign1 = 4'd9; b_sign2 = 4'd13; b_sign3 = 4'd10;
@(posedge clk_i);
a_mant0 = 8'd123; a_mant1 = 8'd153; a_mant2 = 8'd184; a_mant3 = 8'd212;
b_mant0 = 8'd37; b_mant1 = 8'd137; b_mant2 = 8'd16; b_mant3 = 8'd64;
a_exp0 = 10'd808; a_exp1 = 10'd623; a_exp2 = 10'd547; a_exp3 = 10'd723;
b_exp0 = 10'd437; b_exp1 = 10'd519; b_exp2 = 10'd902; b_exp3 = 10'd385;
a_sign0 = 4'd10; a_sign1 = 4'd13; a_sign2 = 4'd6; a_sign3 = 4'd4;
b_sign0 = 4'd10; b_sign1 = 4'd4; b_sign2 = 4'd4; b_sign3 = 4'd10;
@(posedge clk_i);
shared_exps0 = 8'd127;
shared_exps1 = 8'd113;
a_mant0 = 8'd41; a_mant1 = 8'd78; a_mant2 = 8'd171; a_mant3 = 8'd221;
b_mant0 = 8'd17; b_mant1 = 8'd29; b_mant2 = 8'd139; b_mant3 = 8'd137;
a_exp0 = 10'd290; a_exp1 = 10'd876; a_exp2 = 10'd495; a_exp3 = 10'd588;
b_exp0 = 10'd155; b_exp1 = 10'd464; b_exp2 = 10'd13; b_exp3 = 10'd263;
a_sign0 = 4'd0; a_sign1 = 4'd4; a_sign2 = 4'd7; a_sign3 = 4'd0;
b_sign0 = 4'd2; b_sign1 = 4'd9; b_sign2 = 4'd13; b_sign3 = 4'd0;
@(posedge clk_i);
a_mant0 = 8'd143; a_mant1 = 8'd6; a_mant2 = 8'd201; a_mant3 = 8'd87;
b_mant0 = 8'd255; b_mant1 = 8'd20; b_mant2 = 8'd174; b_mant3 = 8'd192;
a_exp0 = 10'd1010; a_exp1 = 10'd176; a_exp2 = 10'd413; a_exp3 = 10'd103;
b_exp0 = 10'd849; b_exp1 = 10'd67; b_exp2 = 10'd891; b_exp3 = 10'd269;
a_sign0 = 4'd11; a_sign1 = 4'd15; a_sign2 = 4'd3; a_sign3 = 4'd1;
b_sign0 = 4'd0; b_sign1 = 4'd0; b_sign2 = 4'd8; b_sign3 = 4'd0;
@(posedge clk_i);
a_mant0 = 8'd236; a_mant1 = 8'd126; a_mant2 = 8'd122; a_mant3 = 8'd211;
b_mant0 = 8'd15; b_mant1 = 8'd191; b_mant2 = 8'd107; b_mant3 = 8'd59;
a_exp0 = 10'd224; a_exp1 = 10'd215; a_exp2 = 10'd846; a_exp3 = 10'd843;
b_exp0 = 10'd210; b_exp1 = 10'd358; b_exp2 = 10'd658; b_exp3 = 10'd909;
a_sign0 = 4'd0; a_sign1 = 4'd0; a_sign2 = 4'd2; a_sign3 = 4'd2;
b_sign0 = 4'd4; b_sign1 = 4'd12; b_sign2 = 4'd12; b_sign3 = 4'd2;
@(posedge clk_i);
a_mant0 = 8'd227; a_mant1 = 8'd64; a_mant2 = 8'd177; a_mant3 = 8'd221;
b_mant0 = 8'd90; b_mant1 = 8'd224; b_mant2 = 8'd82; b_mant3 = 8'd60;
a_exp0 = 10'd302; a_exp1 = 10'd720; a_exp2 = 10'd351; a_exp3 = 10'd300;
b_exp0 = 10'd558; b_exp1 = 10'd785; b_exp2 = 10'd21; b_exp3 = 10'd456;
a_sign0 = 4'd2; a_sign1 = 4'd10; a_sign2 = 4'd1; a_sign3 = 4'd3;
b_sign0 = 4'd14; b_sign1 = 4'd1; b_sign2 = 4'd9; b_sign3 = 4'd7;
@(posedge clk_i);
a_mant0 = 8'd38; a_mant1 = 8'd236; a_mant2 = 8'd255; a_mant3 = 8'd76;
b_mant0 = 8'd62; b_mant1 = 8'd252; b_mant2 = 8'd205; b_mant3 = 8'd113;
a_exp0 = 10'd661; a_exp1 = 10'd633; a_exp2 = 10'd92; a_exp3 = 10'd272;
b_exp0 = 10'd470; b_exp1 = 10'd169; b_exp2 = 10'd585; b_exp3 = 10'd531;
a_sign0 = 4'd0; a_sign1 = 4'd2; a_sign2 = 4'd16; a_sign3 = 4'd11;
b_sign0 = 4'd1; b_sign1 = 4'd12; b_sign2 = 4'd15; b_sign3 = 4'd1;
@(posedge clk_i);
a_mant0 = 8'd113; a_mant1 = 8'd156; a_mant2 = 8'd248; a_mant3 = 8'd154;
b_mant0 = 8'd90; b_mant1 = 8'd138; b_mant2 = 8'd212; b_mant3 = 8'd166;
a_exp0 = 10'd205; a_exp1 = 10'd407; a_exp2 = 10'd825; a_exp3 = 10'd575;
b_exp0 = 10'd714; b_exp1 = 10'd959; b_exp2 = 10'd1010; b_exp3 = 10'd559;
a_sign0 = 4'd13; a_sign1 = 4'd14; a_sign2 = 4'd15; a_sign3 = 4'd8;
b_sign0 = 4'd6; b_sign1 = 4'd3; b_sign2 = 4'd5; b_sign3 = 4'd9;
@(posedge clk_i);
a_mant0 = 8'd232; a_mant1 = 8'd95; a_mant2 = 8'd54; a_mant3 = 8'd167;
b_mant0 = 8'd122; b_mant1 = 8'd25; b_mant2 = 8'd242; b_mant3 = 8'd4;
a_exp0 = 10'd924; a_exp1 = 10'd754; a_exp2 = 10'd726; a_exp3 = 10'd114;
b_exp0 = 10'd164; b_exp1 = 10'd738; b_exp2 = 10'd738; b_exp3 = 10'd714;
a_sign0 = 4'd0; a_sign1 = 4'd4; a_sign2 = 4'd6; a_sign3 = 4'd16;
b_sign0 = 4'd1; b_sign1 = 4'd2; b_sign2 = 4'd15; b_sign3 = 4'd8;
@(posedge clk_i);
a_mant0 = 8'd141; a_mant1 = 8'd158; a_mant2 = 8'd83; a_mant3 = 8'd6;
b_mant0 = 8'd162; b_mant1 = 8'd44; b_mant2 = 8'd152; b_mant3 = 8'd18;
a_exp0 = 10'd373; a_exp1 = 10'd276; a_exp2 = 10'd184; a_exp3 = 10'd784;
b_exp0 = 10'd336; b_exp1 = 10'd247; b_exp2 = 10'd558; b_exp3 = 10'd356;
a_sign0 = 4'd10; a_sign1 = 4'd2; a_sign2 = 4'd0; a_sign3 = 4'd8;
b_sign0 = 4'd6; b_sign1 = 4'd10; b_sign2 = 4'd3; b_sign3 = 4'd12;
@(posedge clk_i);
shared_exps0 = 8'd142;
shared_exps1 = 8'd89;
rstn = 0;
@(posedge clk_i);
rstn = 1;
a_mant0 = 8'd178; a_mant1 = 8'd49; a_mant2 = 8'd139; a_mant3 = 8'd85;
b_mant0 = 8'd165; b_mant1 = 8'd97; b_mant2 = 8'd24; b_mant3 = 8'd181;
a_exp0 = 10'd701; a_exp1 = 10'd742; a_exp2 = 10'd630; a_exp3 = 10'd175;
b_exp0 = 10'd404; b_exp1 = 10'd78; b_exp2 = 10'd141; b_exp3 = 10'd742;
a_sign0 = 4'd9; a_sign1 = 4'd14; a_sign2 = 4'd2; a_sign3 = 4'd7;
b_sign0 = 4'd4; b_sign1 = 4'd14; b_sign2 = 4'd15; b_sign3 = 4'd1;
@(posedge clk_i);
a_mant0 = 8'd242; a_mant1 = 8'd84; a_mant2 = 8'd39; a_mant3 = 8'd39;
b_mant0 = 8'd242; b_mant1 = 8'd83; b_mant2 = 8'd116; b_mant3 = 8'd89;
a_exp0 = 10'd438; a_exp1 = 10'd119; a_exp2 = 10'd192; a_exp3 = 10'd338;
b_exp0 = 10'd453; b_exp1 = 10'd359; b_exp2 = 10'd567; b_exp3 = 10'd97;
a_sign0 = 4'd2; a_sign1 = 4'd4; a_sign2 = 4'd9; a_sign3 = 4'd10;
b_sign0 = 4'd3; b_sign1 = 4'd3; b_sign2 = 4'd3; b_sign3 = 4'd15;
@(posedge clk_i);
a_mant0 = 8'd205; a_mant1 = 8'd34; a_mant2 = 8'd245; a_mant3 = 8'd212;
b_mant0 = 8'd195; b_mant1 = 8'd179; b_mant2 = 8'd74; b_mant3 = 8'd169;
a_exp0 = 10'd669; a_exp1 = 10'd763; a_exp2 = 10'd464; a_exp3 = 10'd761;
b_exp0 = 10'd126; b_exp1 = 10'd159; b_exp2 = 10'd723; b_exp3 = 10'd51;
a_sign0 = 4'd14; a_sign1 = 4'd7; a_sign2 = 4'd0; a_sign3 = 4'd13;
b_sign0 = 4'd9; b_sign1 = 4'd4; b_sign2 = 4'd3; b_sign3 = 4'd15;
@(posedge clk_i);
a_mant0 = 8'd90; a_mant1 = 8'd2; a_mant2 = 8'd178; a_mant3 = 8'd114;
b_mant0 = 8'd7; b_mant1 = 8'd24; b_mant2 = 8'd22; b_mant3 = 8'd65;
a_exp0 = 10'd901; a_exp1 = 10'd342; a_exp2 = 10'd170; a_exp3 = 10'd917;
b_exp0 = 10'd43; b_exp1 = 10'd936; b_exp2 = 10'd112; b_exp3 = 10'd871;
a_sign0 = 4'd8; a_sign1 = 4'd2; a_sign2 = 4'd5; a_sign3 = 4'd0;
b_sign0 = 4'd16; b_sign1 = 4'd4; b_sign2 = 4'd6; b_sign3 = 4'd16;
@(posedge clk_i);
a_mant0 = 8'd131; a_mant1 = 8'd29; a_mant2 = 8'd216; a_mant3 = 8'd222;
b_mant0 = 8'd174; b_mant1 = 8'd49; b_mant2 = 8'd98; b_mant3 = 8'd27;
a_exp0 = 10'd996; a_exp1 = 10'd651; a_exp2 = 10'd782; a_exp3 = 10'd265;
b_exp0 = 10'd417; b_exp1 = 10'd294; b_exp2 = 10'd512; b_exp3 = 10'd188;
a_sign0 = 4'd2; a_sign1 = 4'd11; a_sign2 = 4'd11; a_sign3 = 4'd1;
b_sign0 = 4'd2; b_sign1 = 4'd14; b_sign2 = 4'd3; b_sign3 = 4'd13;
@(posedge clk_i);
a_mant0 = 8'd21; a_mant1 = 8'd184; a_mant2 = 8'd59; a_mant3 = 8'd245;
b_mant0 = 8'd164; b_mant1 = 8'd111; b_mant2 = 8'd90; b_mant3 = 8'd226;
a_exp0 = 10'd862; a_exp1 = 10'd282; a_exp2 = 10'd1006; a_exp3 = 10'd884;
b_exp0 = 10'd47; b_exp1 = 10'd825; b_exp2 = 10'd798; b_exp3 = 10'd321;
a_sign0 = 4'd14; a_sign1 = 4'd6; a_sign2 = 4'd15; a_sign3 = 4'd10;
b_sign0 = 4'd4; b_sign1 = 4'd13; b_sign2 = 4'd14; b_sign3 = 4'd1;
@(posedge clk_i);
a_mant0 = 8'd103; a_mant1 = 8'd253; a_mant2 = 8'd205; a_mant3 = 8'd230;
b_mant0 = 8'd83; b_mant1 = 8'd35; b_mant2 = 8'd248; b_mant3 = 8'd205;
a_exp0 = 10'd331; a_exp1 = 10'd899; a_exp2 = 10'd906; a_exp3 = 10'd194;
b_exp0 = 10'd561; b_exp1 = 10'd183; b_exp2 = 10'd226; b_exp3 = 10'd636;
a_sign0 = 4'd3; a_sign1 = 4'd5; a_sign2 = 4'd3; a_sign3 = 4'd4;
b_sign0 = 4'd0; b_sign1 = 4'd9; b_sign2 = 4'd8; b_sign3 = 4'd10;
@(posedge clk_i);
shared_exps0 = 8'd134;
shared_exps1 = 8'd121;
a_mant0 = 8'd42; a_mant1 = 8'd128; a_mant2 = 8'd196; a_mant3 = 8'd94;
b_mant0 = 8'd239; b_mant1 = 8'd97; b_mant2 = 8'd72; b_mant3 = 8'd204;
a_exp0 = 10'd895; a_exp1 = 10'd113; a_exp2 = 10'd386; a_exp3 = 10'd71;
b_exp0 = 10'd961; b_exp1 = 10'd849; b_exp2 = 10'd566; b_exp3 = 10'd50;
a_sign0 = 4'd9; a_sign1 = 4'd10; a_sign2 = 4'd8; a_sign3 = 4'd12;
b_sign0 = 4'd8; b_sign1 = 4'd12; b_sign2 = 4'd13; b_sign3 = 4'd13;
@(posedge clk_i);
a_mant0 = 8'd129; a_mant1 = 8'd72; a_mant2 = 8'd15; a_mant3 = 8'd67;
b_mant0 = 8'd62; b_mant1 = 8'd87; b_mant2 = 8'd121; b_mant3 = 8'd255;
a_exp0 = 10'd191; a_exp1 = 10'd174; a_exp2 = 10'd5; a_exp3 = 10'd698;
b_exp0 = 10'd675; b_exp1 = 10'd530; b_exp2 = 10'd425; b_exp3 = 10'd229;
a_sign0 = 4'd15; a_sign1 = 4'd12; a_sign2 = 4'd7; a_sign3 = 4'd7;
b_sign0 = 4'd14; b_sign1 = 4'd14; b_sign2 = 4'd3; b_sign3 = 4'd9;
@(posedge clk_i);
a_mant0 = 8'd170; a_mant1 = 8'd232; a_mant2 = 8'd193; a_mant3 = 8'd162;
b_mant0 = 8'd85; b_mant1 = 8'd86; b_mant2 = 8'd176; b_mant3 = 8'd209;
a_exp0 = 10'd806; a_exp1 = 10'd18; a_exp2 = 10'd241; a_exp3 = 10'd834;
b_exp0 = 10'd47; b_exp1 = 10'd181; b_exp2 = 10'd40; b_exp3 = 10'd190;
a_sign0 = 4'd6; a_sign1 = 4'd1; a_sign2 = 4'd10; a_sign3 = 4'd0;
b_sign0 = 4'd7; b_sign1 = 4'd15; b_sign2 = 4'd11; b_sign3 = 4'd15;
@(posedge clk_i);
a_mant0 = 8'd147; a_mant1 = 8'd202; a_mant2 = 8'd87; a_mant3 = 8'd58;
b_mant0 = 8'd237; b_mant1 = 8'd78; b_mant2 = 8'd36; b_mant3 = 8'd214;
a_exp0 = 10'd563; a_exp1 = 10'd532; a_exp2 = 10'd397; a_exp3 = 10'd719;
b_exp0 = 10'd964; b_exp1 = 10'd414; b_exp2 = 10'd342; b_exp3 = 10'd821;
a_sign0 = 4'd4; a_sign1 = 4'd16; a_sign2 = 4'd13; a_sign3 = 4'd13;
b_sign0 = 4'd8; b_sign1 = 4'd7; b_sign2 = 4'd10; b_sign3 = 4'd16;
@(posedge clk_i);
a_mant0 = 8'd211; a_mant1 = 8'd251; a_mant2 = 8'd85; a_mant3 = 8'd174;
b_mant0 = 8'd72; b_mant1 = 8'd206; b_mant2 = 8'd115; b_mant3 = 8'd5;
a_exp0 = 10'd113; a_exp1 = 10'd557; a_exp2 = 10'd37; a_exp3 = 10'd845;
b_exp0 = 10'd657; b_exp1 = 10'd597; b_exp2 = 10'd856; b_exp3 = 10'd434;
a_sign0 = 4'd0; a_sign1 = 4'd9; a_sign2 = 4'd10; a_sign3 = 4'd14;
b_sign0 = 4'd4; b_sign1 = 4'd16; b_sign2 = 4'd14; b_sign3 = 4'd4;
@(posedge clk_i);
a_mant0 = 8'd203; a_mant1 = 8'd31; a_mant2 = 8'd131; a_mant3 = 8'd130;
b_mant0 = 8'd170; b_mant1 = 8'd190; b_mant2 = 8'd248; b_mant3 = 8'd224;
a_exp0 = 10'd976; a_exp1 = 10'd604; a_exp2 = 10'd146; a_exp3 = 10'd238;
b_exp0 = 10'd547; b_exp1 = 10'd943; b_exp2 = 10'd345; b_exp3 = 10'd399;
a_sign0 = 4'd15; a_sign1 = 4'd13; a_sign2 = 4'd15; a_sign3 = 4'd6;
b_sign0 = 4'd15; b_sign1 = 4'd13; b_sign2 = 4'd0; b_sign3 = 4'd4;
@(posedge clk_i);
a_mant0 = 8'd131; a_mant1 = 8'd177; a_mant2 = 8'd118; a_mant3 = 8'd244;
b_mant0 = 8'd163; b_mant1 = 8'd235; b_mant2 = 8'd200; b_mant3 = 8'd179;
a_exp0 = 10'd743; a_exp1 = 10'd432; a_exp2 = 10'd81; a_exp3 = 10'd228;
b_exp0 = 10'd411; b_exp1 = 10'd175; b_exp2 = 10'd666; b_exp3 = 10'd844;
a_sign0 = 4'd4; a_sign1 = 4'd7; a_sign2 = 4'd15; a_sign3 = 4'd16;
b_sign0 = 4'd1; b_sign1 = 4'd10; b_sign2 = 4'd5; b_sign3 = 4'd14;
@(posedge clk_i);
a_mant0 = 8'd232; a_mant1 = 8'd66; a_mant2 = 8'd43; a_mant3 = 8'd145;
b_mant0 = 8'd189; b_mant1 = 8'd227; b_mant2 = 8'd234; b_mant3 = 8'd172;
a_exp0 = 10'd608; a_exp1 = 10'd835; a_exp2 = 10'd502; a_exp3 = 10'd434;
b_exp0 = 10'd210; b_exp1 = 10'd712; b_exp2 = 10'd681; b_exp3 = 10'd871;
a_sign0 = 4'd3; a_sign1 = 4'd3; a_sign2 = 4'd6; a_sign3 = 4'd11;
b_sign0 = 4'd12; b_sign1 = 4'd14; b_sign2 = 4'd10; b_sign3 = 4'd9;
@(posedge clk_i);
shared_exps0 = 8'd135;
shared_exps1 = 8'd103;
a_mant0 = 8'd37; a_mant1 = 8'd8; a_mant2 = 8'd117; a_mant3 = 8'd126;
b_mant0 = 8'd169; b_mant1 = 8'd26; b_mant2 = 8'd211; b_mant3 = 8'd228;
a_exp0 = 10'd243; a_exp1 = 10'd141; a_exp2 = 10'd546; a_exp3 = 10'd653;
b_exp0 = 10'd354; b_exp1 = 10'd1011; b_exp2 = 10'd299; b_exp3 = 10'd551;
a_sign0 = 4'd4; a_sign1 = 4'd13; a_sign2 = 4'd3; a_sign3 = 4'd6;
b_sign0 = 4'd14; b_sign1 = 4'd12; b_sign2 = 4'd9; b_sign3 = 4'd13;
@(posedge clk_i);
a_mant0 = 8'd193; a_mant1 = 8'd164; a_mant2 = 8'd128; a_mant3 = 8'd238;
b_mant0 = 8'd128; b_mant1 = 8'd133; b_mant2 = 8'd98; b_mant3 = 8'd158;
a_exp0 = 10'd924; a_exp1 = 10'd711; a_exp2 = 10'd640; a_exp3 = 10'd761;
b_exp0 = 10'd577; b_exp1 = 10'd710; b_exp2 = 10'd886; b_exp3 = 10'd951;
a_sign0 = 4'd15; a_sign1 = 4'd14; a_sign2 = 4'd6; a_sign3 = 4'd13;
b_sign0 = 4'd1; b_sign1 = 4'd7; b_sign2 = 4'd4; b_sign3 = 4'd6;
@(posedge clk_i);
a_mant0 = 8'd100; a_mant1 = 8'd88; a_mant2 = 8'd53; a_mant3 = 8'd109;
b_mant0 = 8'd219; b_mant1 = 8'd181; b_mant2 = 8'd123; b_mant3 = 8'd71;
a_exp0 = 10'd676; a_exp1 = 10'd550; a_exp2 = 10'd457; a_exp3 = 10'd564;
b_exp0 = 10'd1016; b_exp1 = 10'd576; b_exp2 = 10'd505; b_exp3 = 10'd680;
a_sign0 = 4'd8; a_sign1 = 4'd16; a_sign2 = 4'd16; a_sign3 = 4'd5;
b_sign0 = 4'd6; b_sign1 = 4'd2; b_sign2 = 4'd13; b_sign3 = 4'd6;
@(posedge clk_i);
a_mant0 = 8'd133; a_mant1 = 8'd60; a_mant2 = 8'd118; a_mant3 = 8'd171;
b_mant0 = 8'd126; b_mant1 = 8'd98; b_mant2 = 8'd18; b_mant3 = 8'd157;
a_exp0 = 10'd698; a_exp1 = 10'd357; a_exp2 = 10'd974; a_exp3 = 10'd771;
b_exp0 = 10'd602; b_exp1 = 10'd667; b_exp2 = 10'd38; b_exp3 = 10'd482;
a_sign0 = 4'd3; a_sign1 = 4'd5; a_sign2 = 4'd3; a_sign3 = 4'd5;
b_sign0 = 4'd0; b_sign1 = 4'd10; b_sign2 = 4'd10; b_sign3 = 4'd11;
@(posedge clk_i);
a_mant0 = 8'd224; a_mant1 = 8'd36; a_mant2 = 8'd8; a_mant3 = 8'd138;
b_mant0 = 8'd163; b_mant1 = 8'd217; b_mant2 = 8'd58; b_mant3 = 8'd128;
a_exp0 = 10'd773; a_exp1 = 10'd193; a_exp2 = 10'd554; a_exp3 = 10'd78;
b_exp0 = 10'd345; b_exp1 = 10'd324; b_exp2 = 10'd571; b_exp3 = 10'd82;
a_sign0 = 4'd9; a_sign1 = 4'd3; a_sign2 = 4'd7; a_sign3 = 4'd11;
b_sign0 = 4'd16; b_sign1 = 4'd3; b_sign2 = 4'd3; b_sign3 = 4'd13;
@(posedge clk_i);
a_mant0 = 8'd125; a_mant1 = 8'd112; a_mant2 = 8'd95; a_mant3 = 8'd71;
b_mant0 = 8'd63; b_mant1 = 8'd200; b_mant2 = 8'd33; b_mant3 = 8'd182;
a_exp0 = 10'd770; a_exp1 = 10'd728; a_exp2 = 10'd784; a_exp3 = 10'd601;
b_exp0 = 10'd583; b_exp1 = 10'd122; b_exp2 = 10'd1; b_exp3 = 10'd9;
a_sign0 = 4'd6; a_sign1 = 4'd16; a_sign2 = 4'd12; a_sign3 = 4'd8;
b_sign0 = 4'd5; b_sign1 = 4'd5; b_sign2 = 4'd0; b_sign3 = 4'd2;
@(posedge clk_i);
a_mant0 = 8'd62; a_mant1 = 8'd43; a_mant2 = 8'd70; a_mant3 = 8'd138;
b_mant0 = 8'd113; b_mant1 = 8'd112; b_mant2 = 8'd226; b_mant3 = 8'd117;
a_exp0 = 10'd187; a_exp1 = 10'd75; a_exp2 = 10'd445; a_exp3 = 10'd998;
b_exp0 = 10'd551; b_exp1 = 10'd593; b_exp2 = 10'd991; b_exp3 = 10'd862;
a_sign0 = 4'd16; a_sign1 = 4'd3; a_sign2 = 4'd14; a_sign3 = 4'd8;
b_sign0 = 4'd11; b_sign1 = 4'd3; b_sign2 = 4'd1; b_sign3 = 4'd8;
@(posedge clk_i);
a_mant0 = 8'd172; a_mant1 = 8'd175; a_mant2 = 8'd190; a_mant3 = 8'd90;
b_mant0 = 8'd171; b_mant1 = 8'd216; b_mant2 = 8'd142; b_mant3 = 8'd16;
a_exp0 = 10'd57; a_exp1 = 10'd585; a_exp2 = 10'd492; a_exp3 = 10'd878;
b_exp0 = 10'd83; b_exp1 = 10'd620; b_exp2 = 10'd178; b_exp3 = 10'd778;
a_sign0 = 4'd15; a_sign1 = 4'd0; a_sign2 = 4'd6; a_sign3 = 4'd13;
b_sign0 = 4'd3; b_sign1 = 4'd3; b_sign2 = 4'd5; b_sign3 = 4'd3;
@(posedge clk_i);
shared_exps0 = 8'd103;
shared_exps1 = 8'd124;
a_mant0 = 8'd135; a_mant1 = 8'd29; a_mant2 = 8'd232; a_mant3 = 8'd205;
b_mant0 = 8'd70; b_mant1 = 8'd31; b_mant2 = 8'd4; b_mant3 = 8'd183;
a_exp0 = 10'd457; a_exp1 = 10'd902; a_exp2 = 10'd668; a_exp3 = 10'd140;
b_exp0 = 10'd716; b_exp1 = 10'd310; b_exp2 = 10'd697; b_exp3 = 10'd1016;
a_sign0 = 4'd12; a_sign1 = 4'd11; a_sign2 = 4'd5; a_sign3 = 4'd2;
b_sign0 = 4'd7; b_sign1 = 4'd9; b_sign2 = 4'd16; b_sign3 = 4'd9;
@(posedge clk_i);
a_mant0 = 8'd101; a_mant1 = 8'd107; a_mant2 = 8'd3; a_mant3 = 8'd166;
b_mant0 = 8'd167; b_mant1 = 8'd99; b_mant2 = 8'd53; b_mant3 = 8'd56;
a_exp0 = 10'd419; a_exp1 = 10'd619; a_exp2 = 10'd426; a_exp3 = 10'd21;
b_exp0 = 10'd216; b_exp1 = 10'd289; b_exp2 = 10'd30; b_exp3 = 10'd561;
a_sign0 = 4'd16; a_sign1 = 4'd16; a_sign2 = 4'd5; a_sign3 = 4'd0;
b_sign0 = 4'd6; b_sign1 = 4'd9; b_sign2 = 4'd0; b_sign3 = 4'd6;
@(posedge clk_i);
a_mant0 = 8'd249; a_mant1 = 8'd83; a_mant2 = 8'd46; a_mant3 = 8'd148;
b_mant0 = 8'd156; b_mant1 = 8'd129; b_mant2 = 8'd16; b_mant3 = 8'd239;
a_exp0 = 10'd771; a_exp1 = 10'd675; a_exp2 = 10'd939; a_exp3 = 10'd160;
b_exp0 = 10'd876; b_exp1 = 10'd342; b_exp2 = 10'd471; b_exp3 = 10'd838;
a_sign0 = 4'd8; a_sign1 = 4'd1; a_sign2 = 4'd2; a_sign3 = 4'd14;
b_sign0 = 4'd15; b_sign1 = 4'd1; b_sign2 = 4'd13; b_sign3 = 4'd3;
@(posedge clk_i);
a_mant0 = 8'd238; a_mant1 = 8'd16; a_mant2 = 8'd41; a_mant3 = 8'd75;
b_mant0 = 8'd88; b_mant1 = 8'd36; b_mant2 = 8'd231; b_mant3 = 8'd134;
a_exp0 = 10'd986; a_exp1 = 10'd323; a_exp2 = 10'd680; a_exp3 = 10'd25;
b_exp0 = 10'd1009; b_exp1 = 10'd760; b_exp2 = 10'd4; b_exp3 = 10'd834;
a_sign0 = 4'd0; a_sign1 = 4'd2; a_sign2 = 4'd4; a_sign3 = 4'd12;
b_sign0 = 4'd4; b_sign1 = 4'd2; b_sign2 = 4'd2; b_sign3 = 4'd9;
@(posedge clk_i);
a_mant0 = 8'd104; a_mant1 = 8'd64; a_mant2 = 8'd240; a_mant3 = 8'd169;
b_mant0 = 8'd2; b_mant1 = 8'd44; b_mant2 = 8'd180; b_mant3 = 8'd170;
a_exp0 = 10'd692; a_exp1 = 10'd549; a_exp2 = 10'd833; a_exp3 = 10'd941;
b_exp0 = 10'd842; b_exp1 = 10'd920; b_exp2 = 10'd933; b_exp3 = 10'd39;
a_sign0 = 4'd1; a_sign1 = 4'd7; a_sign2 = 4'd2; a_sign3 = 4'd8;
b_sign0 = 4'd7; b_sign1 = 4'd9; b_sign2 = 4'd2; b_sign3 = 4'd15;
@(posedge clk_i);
a_mant0 = 8'd135; a_mant1 = 8'd97; a_mant2 = 8'd249; a_mant3 = 8'd214;
b_mant0 = 8'd188; b_mant1 = 8'd245; b_mant2 = 8'd19; b_mant3 = 8'd249;
a_exp0 = 10'd522; a_exp1 = 10'd4; a_exp2 = 10'd333; a_exp3 = 10'd819;
b_exp0 = 10'd889; b_exp1 = 10'd527; b_exp2 = 10'd85; b_exp3 = 10'd246;
a_sign0 = 4'd6; a_sign1 = 4'd8; a_sign2 = 4'd14; a_sign3 = 4'd16;
b_sign0 = 4'd12; b_sign1 = 4'd0; b_sign2 = 4'd15; b_sign3 = 4'd7;
@(posedge clk_i);
a_mant0 = 8'd186; a_mant1 = 8'd190; a_mant2 = 8'd50; a_mant3 = 8'd30;
b_mant0 = 8'd100; b_mant1 = 8'd129; b_mant2 = 8'd233; b_mant3 = 8'd138;
a_exp0 = 10'd524; a_exp1 = 10'd90; a_exp2 = 10'd781; a_exp3 = 10'd265;
b_exp0 = 10'd366; b_exp1 = 10'd19; b_exp2 = 10'd431; b_exp3 = 10'd833;
a_sign0 = 4'd10; a_sign1 = 4'd5; a_sign2 = 4'd2; a_sign3 = 4'd8;
b_sign0 = 4'd3; b_sign1 = 4'd11; b_sign2 = 4'd11; b_sign3 = 4'd0;
@(posedge clk_i);
a_mant0 = 8'd165; a_mant1 = 8'd7; a_mant2 = 8'd128; a_mant3 = 8'd9;
b_mant0 = 8'd157; b_mant1 = 8'd178; b_mant2 = 8'd213; b_mant3 = 8'd9;
a_exp0 = 10'd105; a_exp1 = 10'd629; a_exp2 = 10'd69; a_exp3 = 10'd316;
b_exp0 = 10'd587; b_exp1 = 10'd996; b_exp2 = 10'd770; b_exp3 = 10'd131;
a_sign0 = 4'd11; a_sign1 = 4'd10; a_sign2 = 4'd13; a_sign3 = 4'd4;
b_sign0 = 4'd15; b_sign1 = 4'd0; b_sign2 = 4'd9; b_sign3 = 4'd9;
@(posedge clk_i);
shared_exps0 = 8'd124;
shared_exps1 = 8'd131;
rstn = 0;
@(posedge clk_i);
rstn = 1;
a_mant0 = 8'd12; a_mant1 = 8'd48; a_mant2 = 8'd41; a_mant3 = 8'd21;
b_mant0 = 8'd221; b_mant1 = 8'd188; b_mant2 = 8'd226; b_mant3 = 8'd22;
a_exp0 = 10'd724; a_exp1 = 10'd709; a_exp2 = 10'd861; a_exp3 = 10'd221;
b_exp0 = 10'd417; b_exp1 = 10'd784; b_exp2 = 10'd489; b_exp3 = 10'd1013;
a_sign0 = 4'd3; a_sign1 = 4'd0; a_sign2 = 4'd10; a_sign3 = 4'd0;
b_sign0 = 4'd10; b_sign1 = 4'd4; b_sign2 = 4'd14; b_sign3 = 4'd15;
@(posedge clk_i);
a_mant0 = 8'd242; a_mant1 = 8'd41; a_mant2 = 8'd232; a_mant3 = 8'd170;
b_mant0 = 8'd250; b_mant1 = 8'd53; b_mant2 = 8'd47; b_mant3 = 8'd60;
a_exp0 = 10'd198; a_exp1 = 10'd589; a_exp2 = 10'd772; a_exp3 = 10'd540;
b_exp0 = 10'd619; b_exp1 = 10'd874; b_exp2 = 10'd228; b_exp3 = 10'd942;
a_sign0 = 4'd1; a_sign1 = 4'd0; a_sign2 = 4'd16; a_sign3 = 4'd13;
b_sign0 = 4'd7; b_sign1 = 4'd7; b_sign2 = 4'd9; b_sign3 = 4'd2;
@(posedge clk_i);
a_mant0 = 8'd238; a_mant1 = 8'd95; a_mant2 = 8'd166; a_mant3 = 8'd63;
b_mant0 = 8'd152; b_mant1 = 8'd189; b_mant2 = 8'd173; b_mant3 = 8'd78;
a_exp0 = 10'd15; a_exp1 = 10'd232; a_exp2 = 10'd66; a_exp3 = 10'd531;
b_exp0 = 10'd308; b_exp1 = 10'd475; b_exp2 = 10'd730; b_exp3 = 10'd524;
a_sign0 = 4'd0; a_sign1 = 4'd12; a_sign2 = 4'd15; a_sign3 = 4'd11;
b_sign0 = 4'd2; b_sign1 = 4'd5; b_sign2 = 4'd10; b_sign3 = 4'd15;
@(posedge clk_i);
a_mant0 = 8'd186; a_mant1 = 8'd187; a_mant2 = 8'd250; a_mant3 = 8'd14;
b_mant0 = 8'd160; b_mant1 = 8'd73; b_mant2 = 8'd244; b_mant3 = 8'd74;
a_exp0 = 10'd235; a_exp1 = 10'd151; a_exp2 = 10'd867; a_exp3 = 10'd552;
b_exp0 = 10'd814; b_exp1 = 10'd625; b_exp2 = 10'd1009; b_exp3 = 10'd433;
a_sign0 = 4'd7; a_sign1 = 4'd3; a_sign2 = 4'd13; a_sign3 = 4'd10;
b_sign0 = 4'd14; b_sign1 = 4'd6; b_sign2 = 4'd6; b_sign3 = 4'd10;
@(posedge clk_i);
a_mant0 = 8'd32; a_mant1 = 8'd203; a_mant2 = 8'd118; a_mant3 = 8'd144;
b_mant0 = 8'd34; b_mant1 = 8'd147; b_mant2 = 8'd159; b_mant3 = 8'd120;
a_exp0 = 10'd23; a_exp1 = 10'd248; a_exp2 = 10'd722; a_exp3 = 10'd893;
b_exp0 = 10'd586; b_exp1 = 10'd650; b_exp2 = 10'd596; b_exp3 = 10'd552;
a_sign0 = 4'd13; a_sign1 = 4'd6; a_sign2 = 4'd16; a_sign3 = 4'd3;
b_sign0 = 4'd4; b_sign1 = 4'd4; b_sign2 = 4'd2; b_sign3 = 4'd1;
@(posedge clk_i);
a_mant0 = 8'd164; a_mant1 = 8'd27; a_mant2 = 8'd124; a_mant3 = 8'd25;
b_mant0 = 8'd20; b_mant1 = 8'd99; b_mant2 = 8'd151; b_mant3 = 8'd175;
a_exp0 = 10'd959; a_exp1 = 10'd191; a_exp2 = 10'd5; a_exp3 = 10'd183;
b_exp0 = 10'd424; b_exp1 = 10'd316; b_exp2 = 10'd164; b_exp3 = 10'd366;
a_sign0 = 4'd1; a_sign1 = 4'd11; a_sign2 = 4'd1; a_sign3 = 4'd15;
b_sign0 = 4'd6; b_sign1 = 4'd0; b_sign2 = 4'd10; b_sign3 = 4'd9;
@(posedge clk_i);
a_mant0 = 8'd113; a_mant1 = 8'd240; a_mant2 = 8'd212; a_mant3 = 8'd222;
b_mant0 = 8'd248; b_mant1 = 8'd186; b_mant2 = 8'd225; b_mant3 = 8'd188;
a_exp0 = 10'd62; a_exp1 = 10'd766; a_exp2 = 10'd476; a_exp3 = 10'd645;
b_exp0 = 10'd122; b_exp1 = 10'd337; b_exp2 = 10'd249; b_exp3 = 10'd124;
a_sign0 = 4'd11; a_sign1 = 4'd8; a_sign2 = 4'd12; a_sign3 = 4'd8;
b_sign0 = 4'd7; b_sign1 = 4'd4; b_sign2 = 4'd12; b_sign3 = 4'd2;
@(posedge clk_i);
shared_exps0 = 8'd111;
shared_exps1 = 8'd118;
a_mant0 = 8'd60; a_mant1 = 8'd218; a_mant2 = 8'd157; a_mant3 = 8'd64;
b_mant0 = 8'd149; b_mant1 = 8'd34; b_mant2 = 8'd81; b_mant3 = 8'd168;
a_exp0 = 10'd30; a_exp1 = 10'd631; a_exp2 = 10'd153; a_exp3 = 10'd29;
b_exp0 = 10'd663; b_exp1 = 10'd29; b_exp2 = 10'd638; b_exp3 = 10'd504;
a_sign0 = 4'd8; a_sign1 = 4'd5; a_sign2 = 4'd16; a_sign3 = 4'd8;
b_sign0 = 4'd13; b_sign1 = 4'd12; b_sign2 = 4'd4; b_sign3 = 4'd8;
@(posedge clk_i);
a_mant0 = 8'd168; a_mant1 = 8'd64; a_mant2 = 8'd53; a_mant3 = 8'd220;
b_mant0 = 8'd83; b_mant1 = 8'd241; b_mant2 = 8'd54; b_mant3 = 8'd214;
a_exp0 = 10'd700; a_exp1 = 10'd410; a_exp2 = 10'd82; a_exp3 = 10'd129;
b_exp0 = 10'd883; b_exp1 = 10'd485; b_exp2 = 10'd804; b_exp3 = 10'd995;
a_sign0 = 4'd3; a_sign1 = 4'd11; a_sign2 = 4'd3; a_sign3 = 4'd11;
b_sign0 = 4'd5; b_sign1 = 4'd7; b_sign2 = 4'd14; b_sign3 = 4'd8;
@(posedge clk_i);
a_mant0 = 8'd115; a_mant1 = 8'd247; a_mant2 = 8'd11; a_mant3 = 8'd76;
b_mant0 = 8'd167; b_mant1 = 8'd36; b_mant2 = 8'd212; b_mant3 = 8'd72;
a_exp0 = 10'd169; a_exp1 = 10'd490; a_exp2 = 10'd251; a_exp3 = 10'd207;
b_exp0 = 10'd80; b_exp1 = 10'd1015; b_exp2 = 10'd287; b_exp3 = 10'd457;
a_sign0 = 4'd1; a_sign1 = 4'd12; a_sign2 = 4'd13; a_sign3 = 4'd10;
b_sign0 = 4'd10; b_sign1 = 4'd12; b_sign2 = 4'd5; b_sign3 = 4'd3;
@(posedge clk_i);
a_mant0 = 8'd172; a_mant1 = 8'd215; a_mant2 = 8'd224; a_mant3 = 8'd45;
b_mant0 = 8'd146; b_mant1 = 8'd123; b_mant2 = 8'd201; b_mant3 = 8'd186;
a_exp0 = 10'd917; a_exp1 = 10'd876; a_exp2 = 10'd755; a_exp3 = 10'd197;
b_exp0 = 10'd311; b_exp1 = 10'd237; b_exp2 = 10'd472; b_exp3 = 10'd81;
a_sign0 = 4'd16; a_sign1 = 4'd16; a_sign2 = 4'd14; a_sign3 = 4'd13;
b_sign0 = 4'd16; b_sign1 = 4'd14; b_sign2 = 4'd4; b_sign3 = 4'd0;
@(posedge clk_i);
a_mant0 = 8'd16; a_mant1 = 8'd56; a_mant2 = 8'd173; a_mant3 = 8'd114;
b_mant0 = 8'd77; b_mant1 = 8'd88; b_mant2 = 8'd195; b_mant3 = 8'd69;
a_exp0 = 10'd993; a_exp1 = 10'd622; a_exp2 = 10'd708; a_exp3 = 10'd4;
b_exp0 = 10'd603; b_exp1 = 10'd911; b_exp2 = 10'd108; b_exp3 = 10'd317;
a_sign0 = 4'd15; a_sign1 = 4'd11; a_sign2 = 4'd13; a_sign3 = 4'd0;
b_sign0 = 4'd6; b_sign1 = 4'd2; b_sign2 = 4'd8; b_sign3 = 4'd1;
@(posedge clk_i);
a_mant0 = 8'd168; a_mant1 = 8'd133; a_mant2 = 8'd24; a_mant3 = 8'd44;
b_mant0 = 8'd173; b_mant1 = 8'd43; b_mant2 = 8'd166; b_mant3 = 8'd17;
a_exp0 = 10'd168; a_exp1 = 10'd625; a_exp2 = 10'd665; a_exp3 = 10'd937;
b_exp0 = 10'd246; b_exp1 = 10'd529; b_exp2 = 10'd454; b_exp3 = 10'd711;
a_sign0 = 4'd5; a_sign1 = 4'd1; a_sign2 = 4'd14; a_sign3 = 4'd7;
b_sign0 = 4'd14; b_sign1 = 4'd5; b_sign2 = 4'd7; b_sign3 = 4'd15;
@(posedge clk_i);
a_mant0 = 8'd85; a_mant1 = 8'd75; a_mant2 = 8'd166; a_mant3 = 8'd174;
b_mant0 = 8'd47; b_mant1 = 8'd143; b_mant2 = 8'd110; b_mant3 = 8'd131;
a_exp0 = 10'd389; a_exp1 = 10'd459; a_exp2 = 10'd58; a_exp3 = 10'd34;
b_exp0 = 10'd869; b_exp1 = 10'd22; b_exp2 = 10'd625; b_exp3 = 10'd177;
a_sign0 = 4'd11; a_sign1 = 4'd15; a_sign2 = 4'd1; a_sign3 = 4'd16;
b_sign0 = 4'd2; b_sign1 = 4'd12; b_sign2 = 4'd15; b_sign3 = 4'd9;
@(posedge clk_i);
a_mant0 = 8'd222; a_mant1 = 8'd166; a_mant2 = 8'd19; a_mant3 = 8'd214;
b_mant0 = 8'd1; b_mant1 = 8'd205; b_mant2 = 8'd12; b_mant3 = 8'd10;
a_exp0 = 10'd836; a_exp1 = 10'd947; a_exp2 = 10'd529; a_exp3 = 10'd604;
b_exp0 = 10'd362; b_exp1 = 10'd625; b_exp2 = 10'd193; b_exp3 = 10'd889;
a_sign0 = 4'd8; a_sign1 = 4'd8; a_sign2 = 4'd5; a_sign3 = 4'd10;
b_sign0 = 4'd8; b_sign1 = 4'd10; b_sign2 = 4'd13; b_sign3 = 4'd6;
@(posedge clk_i);
shared_exps0 = 8'd107;
shared_exps1 = 8'd144;
a_mant0 = 8'd67; a_mant1 = 8'd247; a_mant2 = 8'd242; a_mant3 = 8'd64;
b_mant0 = 8'd221; b_mant1 = 8'd169; b_mant2 = 8'd39; b_mant3 = 8'd79;
a_exp0 = 10'd996; a_exp1 = 10'd328; a_exp2 = 10'd960; a_exp3 = 10'd1020;
b_exp0 = 10'd501; b_exp1 = 10'd160; b_exp2 = 10'd936; b_exp3 = 10'd968;
a_sign0 = 4'd13; a_sign1 = 4'd11; a_sign2 = 4'd2; a_sign3 = 4'd11;
b_sign0 = 4'd5; b_sign1 = 4'd2; b_sign2 = 4'd16; b_sign3 = 4'd11;
@(posedge clk_i);
a_mant0 = 8'd30; a_mant1 = 8'd122; a_mant2 = 8'd150; a_mant3 = 8'd202;
b_mant0 = 8'd139; b_mant1 = 8'd82; b_mant2 = 8'd107; b_mant3 = 8'd65;
a_exp0 = 10'd705; a_exp1 = 10'd943; a_exp2 = 10'd408; a_exp3 = 10'd865;
b_exp0 = 10'd68; b_exp1 = 10'd1007; b_exp2 = 10'd755; b_exp3 = 10'd257;
a_sign0 = 4'd8; a_sign1 = 4'd8; a_sign2 = 4'd7; a_sign3 = 4'd14;
b_sign0 = 4'd12; b_sign1 = 4'd2; b_sign2 = 4'd13; b_sign3 = 4'd9;
@(posedge clk_i);
a_mant0 = 8'd25; a_mant1 = 8'd76; a_mant2 = 8'd80; a_mant3 = 8'd17;
b_mant0 = 8'd24; b_mant1 = 8'd22; b_mant2 = 8'd90; b_mant3 = 8'd58;
a_exp0 = 10'd175; a_exp1 = 10'd917; a_exp2 = 10'd783; a_exp3 = 10'd829;
b_exp0 = 10'd249; b_exp1 = 10'd807; b_exp2 = 10'd888; b_exp3 = 10'd570;
a_sign0 = 4'd13; a_sign1 = 4'd0; a_sign2 = 4'd8; a_sign3 = 4'd10;
b_sign0 = 4'd4; b_sign1 = 4'd11; b_sign2 = 4'd4; b_sign3 = 4'd12;
@(posedge clk_i);
a_mant0 = 8'd79; a_mant1 = 8'd118; a_mant2 = 8'd98; a_mant3 = 8'd220;
b_mant0 = 8'd100; b_mant1 = 8'd241; b_mant2 = 8'd111; b_mant3 = 8'd220;
a_exp0 = 10'd187; a_exp1 = 10'd843; a_exp2 = 10'd322; a_exp3 = 10'd211;
b_exp0 = 10'd526; b_exp1 = 10'd842; b_exp2 = 10'd521; b_exp3 = 10'd464;
a_sign0 = 4'd5; a_sign1 = 4'd1; a_sign2 = 4'd13; a_sign3 = 4'd1;
b_sign0 = 4'd7; b_sign1 = 4'd15; b_sign2 = 4'd13; b_sign3 = 4'd0;
@(posedge clk_i);
a_mant0 = 8'd106; a_mant1 = 8'd250; a_mant2 = 8'd73; a_mant3 = 8'd18;
b_mant0 = 8'd148; b_mant1 = 8'd47; b_mant2 = 8'd154; b_mant3 = 8'd16;
a_exp0 = 10'd788; a_exp1 = 10'd296; a_exp2 = 10'd277; a_exp3 = 10'd265;
b_exp0 = 10'd351; b_exp1 = 10'd245; b_exp2 = 10'd899; b_exp3 = 10'd407;
a_sign0 = 4'd2; a_sign1 = 4'd7; a_sign2 = 4'd14; a_sign3 = 4'd8;
b_sign0 = 4'd9; b_sign1 = 4'd12; b_sign2 = 4'd10; b_sign3 = 4'd11;
@(posedge clk_i);
a_mant0 = 8'd212; a_mant1 = 8'd7; a_mant2 = 8'd19; a_mant3 = 8'd193;
b_mant0 = 8'd239; b_mant1 = 8'd133; b_mant2 = 8'd147; b_mant3 = 8'd192;
a_exp0 = 10'd722; a_exp1 = 10'd868; a_exp2 = 10'd648; a_exp3 = 10'd437;
b_exp0 = 10'd356; b_exp1 = 10'd992; b_exp2 = 10'd590; b_exp3 = 10'd58;
a_sign0 = 4'd3; a_sign1 = 4'd5; a_sign2 = 4'd16; a_sign3 = 4'd15;
b_sign0 = 4'd14; b_sign1 = 4'd11; b_sign2 = 4'd11; b_sign3 = 4'd2;
@(posedge clk_i);
a_mant0 = 8'd47; a_mant1 = 8'd18; a_mant2 = 8'd146; a_mant3 = 8'd255;
b_mant0 = 8'd167; b_mant1 = 8'd71; b_mant2 = 8'd139; b_mant3 = 8'd152;
a_exp0 = 10'd1020; a_exp1 = 10'd55; a_exp2 = 10'd791; a_exp3 = 10'd865;
b_exp0 = 10'd1004; b_exp1 = 10'd134; b_exp2 = 10'd286; b_exp3 = 10'd132;
a_sign0 = 4'd15; a_sign1 = 4'd11; a_sign2 = 4'd1; a_sign3 = 4'd7;
b_sign0 = 4'd15; b_sign1 = 4'd10; b_sign2 = 4'd16; b_sign3 = 4'd14;
@(posedge clk_i);
a_mant0 = 8'd239; a_mant1 = 8'd55; a_mant2 = 8'd222; a_mant3 = 8'd21;
b_mant0 = 8'd63; b_mant1 = 8'd43; b_mant2 = 8'd232; b_mant3 = 8'd235;
a_exp0 = 10'd605; a_exp1 = 10'd888; a_exp2 = 10'd202; a_exp3 = 10'd72;
b_exp0 = 10'd330; b_exp1 = 10'd651; b_exp2 = 10'd224; b_exp3 = 10'd625;
a_sign0 = 4'd12; a_sign1 = 4'd16; a_sign2 = 4'd7; a_sign3 = 4'd6;
b_sign0 = 4'd9; b_sign1 = 4'd2; b_sign2 = 4'd12; b_sign3 = 4'd9;
@(posedge clk_i);
shared_exps0 = 8'd121;
shared_exps1 = 8'd125;
a_mant0 = 8'd227; a_mant1 = 8'd208; a_mant2 = 8'd235; a_mant3 = 8'd142;
b_mant0 = 8'd246; b_mant1 = 8'd44; b_mant2 = 8'd191; b_mant3 = 8'd136;
a_exp0 = 10'd0; a_exp1 = 10'd174; a_exp2 = 10'd8; a_exp3 = 10'd603;
b_exp0 = 10'd236; b_exp1 = 10'd140; b_exp2 = 10'd13; b_exp3 = 10'd83;
a_sign0 = 4'd16; a_sign1 = 4'd0; a_sign2 = 4'd5; a_sign3 = 4'd3;
b_sign0 = 4'd5; b_sign1 = 4'd4; b_sign2 = 4'd4; b_sign3 = 4'd14;
@(posedge clk_i);
a_mant0 = 8'd60; a_mant1 = 8'd216; a_mant2 = 8'd81; a_mant3 = 8'd183;
b_mant0 = 8'd182; b_mant1 = 8'd98; b_mant2 = 8'd141; b_mant3 = 8'd107;
a_exp0 = 10'd485; a_exp1 = 10'd168; a_exp2 = 10'd344; a_exp3 = 10'd60;
b_exp0 = 10'd773; b_exp1 = 10'd945; b_exp2 = 10'd598; b_exp3 = 10'd441;
a_sign0 = 4'd8; a_sign1 = 4'd15; a_sign2 = 4'd1; a_sign3 = 4'd2;
b_sign0 = 4'd16; b_sign1 = 4'd9; b_sign2 = 4'd6; b_sign3 = 4'd13;
@(posedge clk_i);
a_mant0 = 8'd138; a_mant1 = 8'd190; a_mant2 = 8'd35; a_mant3 = 8'd97;
b_mant0 = 8'd70; b_mant1 = 8'd230; b_mant2 = 8'd216; b_mant3 = 8'd172;
a_exp0 = 10'd828; a_exp1 = 10'd852; a_exp2 = 10'd1009; a_exp3 = 10'd791;
b_exp0 = 10'd588; b_exp1 = 10'd889; b_exp2 = 10'd390; b_exp3 = 10'd1023;
a_sign0 = 4'd14; a_sign1 = 4'd13; a_sign2 = 4'd8; a_sign3 = 4'd9;
b_sign0 = 4'd6; b_sign1 = 4'd11; b_sign2 = 4'd15; b_sign3 = 4'd11;
@(posedge clk_i);
a_mant0 = 8'd136; a_mant1 = 8'd33; a_mant2 = 8'd129; a_mant3 = 8'd29;
b_mant0 = 8'd58; b_mant1 = 8'd196; b_mant2 = 8'd174; b_mant3 = 8'd138;
a_exp0 = 10'd910; a_exp1 = 10'd421; a_exp2 = 10'd617; a_exp3 = 10'd327;
b_exp0 = 10'd1002; b_exp1 = 10'd88; b_exp2 = 10'd225; b_exp3 = 10'd466;
a_sign0 = 4'd8; a_sign1 = 4'd11; a_sign2 = 4'd11; a_sign3 = 4'd10;
b_sign0 = 4'd0; b_sign1 = 4'd1; b_sign2 = 4'd9; b_sign3 = 4'd3;
@(posedge clk_i);
a_mant0 = 8'd18; a_mant1 = 8'd140; a_mant2 = 8'd65; a_mant3 = 8'd76;
b_mant0 = 8'd2; b_mant1 = 8'd192; b_mant2 = 8'd193; b_mant3 = 8'd212;
a_exp0 = 10'd709; a_exp1 = 10'd368; a_exp2 = 10'd811; a_exp3 = 10'd608;
b_exp0 = 10'd503; b_exp1 = 10'd371; b_exp2 = 10'd362; b_exp3 = 10'd175;
a_sign0 = 4'd15; a_sign1 = 4'd4; a_sign2 = 4'd16; a_sign3 = 4'd7;
b_sign0 = 4'd12; b_sign1 = 4'd11; b_sign2 = 4'd10; b_sign3 = 4'd2;
@(posedge clk_i);
a_mant0 = 8'd90; a_mant1 = 8'd90; a_mant2 = 8'd148; a_mant3 = 8'd51;
b_mant0 = 8'd84; b_mant1 = 8'd133; b_mant2 = 8'd72; b_mant3 = 8'd196;
a_exp0 = 10'd358; a_exp1 = 10'd728; a_exp2 = 10'd537; a_exp3 = 10'd208;
b_exp0 = 10'd617; b_exp1 = 10'd122; b_exp2 = 10'd749; b_exp3 = 10'd219;
a_sign0 = 4'd2; a_sign1 = 4'd9; a_sign2 = 4'd6; a_sign3 = 4'd14;
b_sign0 = 4'd6; b_sign1 = 4'd13; b_sign2 = 4'd8; b_sign3 = 4'd9;
@(posedge clk_i);
a_mant0 = 8'd46; a_mant1 = 8'd217; a_mant2 = 8'd101; a_mant3 = 8'd231;
b_mant0 = 8'd247; b_mant1 = 8'd126; b_mant2 = 8'd70; b_mant3 = 8'd48;
a_exp0 = 10'd148; a_exp1 = 10'd6; a_exp2 = 10'd905; a_exp3 = 10'd210;
b_exp0 = 10'd130; b_exp1 = 10'd1015; b_exp2 = 10'd841; b_exp3 = 10'd364;
a_sign0 = 4'd7; a_sign1 = 4'd9; a_sign2 = 4'd16; a_sign3 = 4'd5;
b_sign0 = 4'd12; b_sign1 = 4'd16; b_sign2 = 4'd7; b_sign3 = 4'd12;
@(posedge clk_i);
a_mant0 = 8'd125; a_mant1 = 8'd1; a_mant2 = 8'd198; a_mant3 = 8'd38;
b_mant0 = 8'd119; b_mant1 = 8'd63; b_mant2 = 8'd46; b_mant3 = 8'd209;
a_exp0 = 10'd226; a_exp1 = 10'd404; a_exp2 = 10'd700; a_exp3 = 10'd297;
b_exp0 = 10'd389; b_exp1 = 10'd393; b_exp2 = 10'd363; b_exp3 = 10'd750;
a_sign0 = 4'd13; a_sign1 = 4'd11; a_sign2 = 4'd15; a_sign3 = 4'd5;
b_sign0 = 4'd3; b_sign1 = 4'd9; b_sign2 = 4'd15; b_sign3 = 4'd12;
@(posedge clk_i);
shared_exps0 = 8'd139;
shared_exps1 = 8'd143;
rstn = 0;
@(posedge clk_i);
rstn = 1;
a_mant0 = 8'd17; a_mant1 = 8'd84; a_mant2 = 8'd230; a_mant3 = 8'd149;
b_mant0 = 8'd80; b_mant1 = 8'd246; b_mant2 = 8'd114; b_mant3 = 8'd196;
a_exp0 = 10'd988; a_exp1 = 10'd173; a_exp2 = 10'd576; a_exp3 = 10'd517;
b_exp0 = 10'd361; b_exp1 = 10'd214; b_exp2 = 10'd227; b_exp3 = 10'd639;
a_sign0 = 4'd1; a_sign1 = 4'd2; a_sign2 = 4'd4; a_sign3 = 4'd16;
b_sign0 = 4'd1; b_sign1 = 4'd8; b_sign2 = 4'd0; b_sign3 = 4'd4;
@(posedge clk_i);
a_mant0 = 8'd197; a_mant1 = 8'd192; a_mant2 = 8'd215; a_mant3 = 8'd217;
b_mant0 = 8'd71; b_mant1 = 8'd137; b_mant2 = 8'd110; b_mant3 = 8'd180;
a_exp0 = 10'd765; a_exp1 = 10'd308; a_exp2 = 10'd193; a_exp3 = 10'd673;
b_exp0 = 10'd573; b_exp1 = 10'd655; b_exp2 = 10'd104; b_exp3 = 10'd880;
a_sign0 = 4'd14; a_sign1 = 4'd9; a_sign2 = 4'd6; a_sign3 = 4'd16;
b_sign0 = 4'd8; b_sign1 = 4'd10; b_sign2 = 4'd9; b_sign3 = 4'd11;
@(posedge clk_i);
a_mant0 = 8'd45; a_mant1 = 8'd240; a_mant2 = 8'd218; a_mant3 = 8'd206;
b_mant0 = 8'd194; b_mant1 = 8'd235; b_mant2 = 8'd152; b_mant3 = 8'd178;
a_exp0 = 10'd986; a_exp1 = 10'd213; a_exp2 = 10'd975; a_exp3 = 10'd149;
b_exp0 = 10'd149; b_exp1 = 10'd709; b_exp2 = 10'd955; b_exp3 = 10'd415;
a_sign0 = 4'd13; a_sign1 = 4'd2; a_sign2 = 4'd4; a_sign3 = 4'd2;
b_sign0 = 4'd7; b_sign1 = 4'd4; b_sign2 = 4'd10; b_sign3 = 4'd4;
@(posedge clk_i);
a_mant0 = 8'd221; a_mant1 = 8'd8; a_mant2 = 8'd129; a_mant3 = 8'd66;
b_mant0 = 8'd135; b_mant1 = 8'd97; b_mant2 = 8'd43; b_mant3 = 8'd150;
a_exp0 = 10'd800; a_exp1 = 10'd826; a_exp2 = 10'd455; a_exp3 = 10'd530;
b_exp0 = 10'd727; b_exp1 = 10'd399; b_exp2 = 10'd218; b_exp3 = 10'd823;
a_sign0 = 4'd8; a_sign1 = 4'd3; a_sign2 = 4'd13; a_sign3 = 4'd7;
b_sign0 = 4'd6; b_sign1 = 4'd3; b_sign2 = 4'd13; b_sign3 = 4'd16;
@(posedge clk_i);
a_mant0 = 8'd160; a_mant1 = 8'd185; a_mant2 = 8'd138; a_mant3 = 8'd165;
b_mant0 = 8'd9; b_mant1 = 8'd35; b_mant2 = 8'd210; b_mant3 = 8'd202;
a_exp0 = 10'd35; a_exp1 = 10'd294; a_exp2 = 10'd499; a_exp3 = 10'd506;
b_exp0 = 10'd618; b_exp1 = 10'd469; b_exp2 = 10'd62; b_exp3 = 10'd484;
a_sign0 = 4'd5; a_sign1 = 4'd6; a_sign2 = 4'd12; a_sign3 = 4'd1;
b_sign0 = 4'd9; b_sign1 = 4'd11; b_sign2 = 4'd8; b_sign3 = 4'd13;
@(posedge clk_i);
a_mant0 = 8'd203; a_mant1 = 8'd124; a_mant2 = 8'd202; a_mant3 = 8'd91;
b_mant0 = 8'd47; b_mant1 = 8'd11; b_mant2 = 8'd16; b_mant3 = 8'd45;
a_exp0 = 10'd572; a_exp1 = 10'd614; a_exp2 = 10'd434; a_exp3 = 10'd452;
b_exp0 = 10'd959; b_exp1 = 10'd118; b_exp2 = 10'd222; b_exp3 = 10'd308;
a_sign0 = 4'd16; a_sign1 = 4'd6; a_sign2 = 4'd6; a_sign3 = 4'd2;
b_sign0 = 4'd9; b_sign1 = 4'd12; b_sign2 = 4'd8; b_sign3 = 4'd13;
@(posedge clk_i);
a_mant0 = 8'd78; a_mant1 = 8'd99; a_mant2 = 8'd222; a_mant3 = 8'd34;
b_mant0 = 8'd63; b_mant1 = 8'd77; b_mant2 = 8'd13; b_mant3 = 8'd92;
a_exp0 = 10'd502; a_exp1 = 10'd813; a_exp2 = 10'd378; a_exp3 = 10'd226;
b_exp0 = 10'd554; b_exp1 = 10'd963; b_exp2 = 10'd816; b_exp3 = 10'd433;
a_sign0 = 4'd13; a_sign1 = 4'd11; a_sign2 = 4'd16; a_sign3 = 4'd14;
b_sign0 = 4'd1; b_sign1 = 4'd15; b_sign2 = 4'd7; b_sign3 = 4'd0;
@(posedge clk_i);
shared_exps0 = 8'd154;
shared_exps1 = 8'd125;
a_mant0 = 8'd237; a_mant1 = 8'd196; a_mant2 = 8'd133; a_mant3 = 8'd25;
b_mant0 = 8'd82; b_mant1 = 8'd173; b_mant2 = 8'd2; b_mant3 = 8'd244;
a_exp0 = 10'd190; a_exp1 = 10'd121; a_exp2 = 10'd204; a_exp3 = 10'd101;
b_exp0 = 10'd756; b_exp1 = 10'd408; b_exp2 = 10'd552; b_exp3 = 10'd949;
a_sign0 = 4'd6; a_sign1 = 4'd7; a_sign2 = 4'd8; a_sign3 = 4'd13;
b_sign0 = 4'd4; b_sign1 = 4'd0; b_sign2 = 4'd5; b_sign3 = 4'd1;
@(posedge clk_i);
a_mant0 = 8'd9; a_mant1 = 8'd26; a_mant2 = 8'd251; a_mant3 = 8'd200;
b_mant0 = 8'd154; b_mant1 = 8'd144; b_mant2 = 8'd119; b_mant3 = 8'd16;
a_exp0 = 10'd846; a_exp1 = 10'd855; a_exp2 = 10'd48; a_exp3 = 10'd536;
b_exp0 = 10'd929; b_exp1 = 10'd295; b_exp2 = 10'd821; b_exp3 = 10'd694;
a_sign0 = 4'd8; a_sign1 = 4'd12; a_sign2 = 4'd9; a_sign3 = 4'd11;
b_sign0 = 4'd3; b_sign1 = 4'd9; b_sign2 = 4'd13; b_sign3 = 4'd13;
@(posedge clk_i);
a_mant0 = 8'd235; a_mant1 = 8'd237; a_mant2 = 8'd77; a_mant3 = 8'd244;
b_mant0 = 8'd30; b_mant1 = 8'd69; b_mant2 = 8'd63; b_mant3 = 8'd242;
a_exp0 = 10'd497; a_exp1 = 10'd64; a_exp2 = 10'd425; a_exp3 = 10'd320;
b_exp0 = 10'd869; b_exp1 = 10'd185; b_exp2 = 10'd142; b_exp3 = 10'd617;
a_sign0 = 4'd15; a_sign1 = 4'd16; a_sign2 = 4'd9; a_sign3 = 4'd8;
b_sign0 = 4'd12; b_sign1 = 4'd8; b_sign2 = 4'd13; b_sign3 = 4'd10;
@(posedge clk_i);
a_mant0 = 8'd138; a_mant1 = 8'd35; a_mant2 = 8'd219; a_mant3 = 8'd4;
b_mant0 = 8'd245; b_mant1 = 8'd125; b_mant2 = 8'd37; b_mant3 = 8'd110;
a_exp0 = 10'd878; a_exp1 = 10'd382; a_exp2 = 10'd699; a_exp3 = 10'd373;
b_exp0 = 10'd263; b_exp1 = 10'd52; b_exp2 = 10'd132; b_exp3 = 10'd32;
a_sign0 = 4'd8; a_sign1 = 4'd7; a_sign2 = 4'd3; a_sign3 = 4'd0;
b_sign0 = 4'd1; b_sign1 = 4'd16; b_sign2 = 4'd3; b_sign3 = 4'd7;
@(posedge clk_i);
a_mant0 = 8'd169; a_mant1 = 8'd124; a_mant2 = 8'd41; a_mant3 = 8'd141;
b_mant0 = 8'd235; b_mant1 = 8'd213; b_mant2 = 8'd189; b_mant3 = 8'd249;
a_exp0 = 10'd468; a_exp1 = 10'd506; a_exp2 = 10'd970; a_exp3 = 10'd667;
b_exp0 = 10'd509; b_exp1 = 10'd575; b_exp2 = 10'd586; b_exp3 = 10'd511;
a_sign0 = 4'd14; a_sign1 = 4'd3; a_sign2 = 4'd12; a_sign3 = 4'd1;
b_sign0 = 4'd8; b_sign1 = 4'd1; b_sign2 = 4'd12; b_sign3 = 4'd7;
@(posedge clk_i);
a_mant0 = 8'd142; a_mant1 = 8'd69; a_mant2 = 8'd66; a_mant3 = 8'd162;
b_mant0 = 8'd118; b_mant1 = 8'd28; b_mant2 = 8'd244; b_mant3 = 8'd86;
a_exp0 = 10'd340; a_exp1 = 10'd430; a_exp2 = 10'd179; a_exp3 = 10'd898;
b_exp0 = 10'd668; b_exp1 = 10'd271; b_exp2 = 10'd913; b_exp3 = 10'd983;
a_sign0 = 4'd1; a_sign1 = 4'd16; a_sign2 = 4'd7; a_sign3 = 4'd2;
b_sign0 = 4'd3; b_sign1 = 4'd13; b_sign2 = 4'd0; b_sign3 = 4'd0;
@(posedge clk_i);
a_mant0 = 8'd134; a_mant1 = 8'd217; a_mant2 = 8'd2; a_mant3 = 8'd247;
b_mant0 = 8'd174; b_mant1 = 8'd75; b_mant2 = 8'd218; b_mant3 = 8'd194;
a_exp0 = 10'd761; a_exp1 = 10'd1002; a_exp2 = 10'd164; a_exp3 = 10'd797;
b_exp0 = 10'd649; b_exp1 = 10'd450; b_exp2 = 10'd945; b_exp3 = 10'd588;
a_sign0 = 4'd13; a_sign1 = 4'd3; a_sign2 = 4'd2; a_sign3 = 4'd5;
b_sign0 = 4'd7; b_sign1 = 4'd8; b_sign2 = 4'd2; b_sign3 = 4'd8;
@(posedge clk_i);
a_mant0 = 8'd26; a_mant1 = 8'd68; a_mant2 = 8'd63; a_mant3 = 8'd18;
b_mant0 = 8'd113; b_mant1 = 8'd17; b_mant2 = 8'd38; b_mant3 = 8'd42;
a_exp0 = 10'd573; a_exp1 = 10'd152; a_exp2 = 10'd686; a_exp3 = 10'd305;
b_exp0 = 10'd987; b_exp1 = 10'd617; b_exp2 = 10'd483; b_exp3 = 10'd11;
a_sign0 = 4'd15; a_sign1 = 4'd9; a_sign2 = 4'd6; a_sign3 = 4'd0;
b_sign0 = 4'd13; b_sign1 = 4'd0; b_sign2 = 4'd11; b_sign3 = 4'd4;
@(posedge clk_i);
shared_exps0 = 8'd129;
shared_exps1 = 8'd131;
a_mant0 = 8'd100; a_mant1 = 8'd174; a_mant2 = 8'd134; a_mant3 = 8'd245;
b_mant0 = 8'd65; b_mant1 = 8'd239; b_mant2 = 8'd70; b_mant3 = 8'd112;
a_exp0 = 10'd490; a_exp1 = 10'd396; a_exp2 = 10'd526; a_exp3 = 10'd136;
b_exp0 = 10'd315; b_exp1 = 10'd106; b_exp2 = 10'd378; b_exp3 = 10'd42;
a_sign0 = 4'd14; a_sign1 = 4'd14; a_sign2 = 4'd1; a_sign3 = 4'd6;
b_sign0 = 4'd4; b_sign1 = 4'd12; b_sign2 = 4'd7; b_sign3 = 4'd0;
@(posedge clk_i);
a_mant0 = 8'd2; a_mant1 = 8'd133; a_mant2 = 8'd249; a_mant3 = 8'd108;
b_mant0 = 8'd133; b_mant1 = 8'd44; b_mant2 = 8'd212; b_mant3 = 8'd252;
a_exp0 = 10'd78; a_exp1 = 10'd168; a_exp2 = 10'd1008; a_exp3 = 10'd219;
b_exp0 = 10'd230; b_exp1 = 10'd912; b_exp2 = 10'd3; b_exp3 = 10'd73;
a_sign0 = 4'd9; a_sign1 = 4'd10; a_sign2 = 4'd2; a_sign3 = 4'd9;
b_sign0 = 4'd1; b_sign1 = 4'd8; b_sign2 = 4'd12; b_sign3 = 4'd14;
@(posedge clk_i);
a_mant0 = 8'd51; a_mant1 = 8'd87; a_mant2 = 8'd90; a_mant3 = 8'd103;
b_mant0 = 8'd55; b_mant1 = 8'd29; b_mant2 = 8'd88; b_mant3 = 8'd195;
a_exp0 = 10'd955; a_exp1 = 10'd541; a_exp2 = 10'd454; a_exp3 = 10'd99;
b_exp0 = 10'd655; b_exp1 = 10'd865; b_exp2 = 10'd979; b_exp3 = 10'd857;
a_sign0 = 4'd16; a_sign1 = 4'd15; a_sign2 = 4'd5; a_sign3 = 4'd6;
b_sign0 = 4'd10; b_sign1 = 4'd9; b_sign2 = 4'd2; b_sign3 = 4'd12;
@(posedge clk_i);
a_mant0 = 8'd242; a_mant1 = 8'd120; a_mant2 = 8'd175; a_mant3 = 8'd215;
b_mant0 = 8'd25; b_mant1 = 8'd46; b_mant2 = 8'd208; b_mant3 = 8'd137;
a_exp0 = 10'd218; a_exp1 = 10'd617; a_exp2 = 10'd146; a_exp3 = 10'd511;
b_exp0 = 10'd251; b_exp1 = 10'd436; b_exp2 = 10'd83; b_exp3 = 10'd837;
a_sign0 = 4'd14; a_sign1 = 4'd9; a_sign2 = 4'd6; a_sign3 = 4'd14;
b_sign0 = 4'd9; b_sign1 = 4'd7; b_sign2 = 4'd4; b_sign3 = 4'd3;
@(posedge clk_i);
a_mant0 = 8'd117; a_mant1 = 8'd242; a_mant2 = 8'd0; a_mant3 = 8'd55;
b_mant0 = 8'd207; b_mant1 = 8'd248; b_mant2 = 8'd120; b_mant3 = 8'd247;
a_exp0 = 10'd210; a_exp1 = 10'd840; a_exp2 = 10'd426; a_exp3 = 10'd444;
b_exp0 = 10'd774; b_exp1 = 10'd844; b_exp2 = 10'd594; b_exp3 = 10'd1007;
a_sign0 = 4'd0; a_sign1 = 4'd9; a_sign2 = 4'd5; a_sign3 = 4'd5;
b_sign0 = 4'd4; b_sign1 = 4'd12; b_sign2 = 4'd8; b_sign3 = 4'd4;
@(posedge clk_i);
a_mant0 = 8'd199; a_mant1 = 8'd16; a_mant2 = 8'd82; a_mant3 = 8'd205;
b_mant0 = 8'd183; b_mant1 = 8'd209; b_mant2 = 8'd254; b_mant3 = 8'd91;
a_exp0 = 10'd2; a_exp1 = 10'd756; a_exp2 = 10'd415; a_exp3 = 10'd800;
b_exp0 = 10'd777; b_exp1 = 10'd54; b_exp2 = 10'd34; b_exp3 = 10'd552;
a_sign0 = 4'd6; a_sign1 = 4'd7; a_sign2 = 4'd9; a_sign3 = 4'd3;
b_sign0 = 4'd16; b_sign1 = 4'd1; b_sign2 = 4'd0; b_sign3 = 4'd0;
@(posedge clk_i);
a_mant0 = 8'd101; a_mant1 = 8'd223; a_mant2 = 8'd61; a_mant3 = 8'd92;
b_mant0 = 8'd149; b_mant1 = 8'd73; b_mant2 = 8'd192; b_mant3 = 8'd77;
a_exp0 = 10'd987; a_exp1 = 10'd603; a_exp2 = 10'd23; a_exp3 = 10'd921;
b_exp0 = 10'd212; b_exp1 = 10'd465; b_exp2 = 10'd451; b_exp3 = 10'd202;
a_sign0 = 4'd11; a_sign1 = 4'd10; a_sign2 = 4'd2; a_sign3 = 4'd10;
b_sign0 = 4'd14; b_sign1 = 4'd15; b_sign2 = 4'd14; b_sign3 = 4'd6;
@(posedge clk_i);
a_mant0 = 8'd42; a_mant1 = 8'd102; a_mant2 = 8'd7; a_mant3 = 8'd189;
b_mant0 = 8'd176; b_mant1 = 8'd220; b_mant2 = 8'd191; b_mant3 = 8'd24;
a_exp0 = 10'd513; a_exp1 = 10'd491; a_exp2 = 10'd246; a_exp3 = 10'd600;
b_exp0 = 10'd730; b_exp1 = 10'd572; b_exp2 = 10'd164; b_exp3 = 10'd183;
a_sign0 = 4'd4; a_sign1 = 4'd7; a_sign2 = 4'd10; a_sign3 = 4'd12;
b_sign0 = 4'd9; b_sign1 = 4'd12; b_sign2 = 4'd10; b_sign3 = 4'd13;
@(posedge clk_i);
shared_exps0 = 8'd144;
shared_exps1 = 8'd128;
a_mant0 = 8'd173; a_mant1 = 8'd159; a_mant2 = 8'd39; a_mant3 = 8'd204;
b_mant0 = 8'd172; b_mant1 = 8'd61; b_mant2 = 8'd122; b_mant3 = 8'd236;
a_exp0 = 10'd92; a_exp1 = 10'd645; a_exp2 = 10'd630; a_exp3 = 10'd62;
b_exp0 = 10'd480; b_exp1 = 10'd966; b_exp2 = 10'd239; b_exp3 = 10'd825;
a_sign0 = 4'd10; a_sign1 = 4'd5; a_sign2 = 4'd7; a_sign3 = 4'd1;
b_sign0 = 4'd16; b_sign1 = 4'd3; b_sign2 = 4'd6; b_sign3 = 4'd2;
@(posedge clk_i);
a_mant0 = 8'd83; a_mant1 = 8'd50; a_mant2 = 8'd146; a_mant3 = 8'd74;
b_mant0 = 8'd74; b_mant1 = 8'd38; b_mant2 = 8'd75; b_mant3 = 8'd183;
a_exp0 = 10'd104; a_exp1 = 10'd769; a_exp2 = 10'd1010; a_exp3 = 10'd590;
b_exp0 = 10'd811; b_exp1 = 10'd425; b_exp2 = 10'd539; b_exp3 = 10'd187;
a_sign0 = 4'd3; a_sign1 = 4'd15; a_sign2 = 4'd3; a_sign3 = 4'd1;
b_sign0 = 4'd4; b_sign1 = 4'd1; b_sign2 = 4'd12; b_sign3 = 4'd4;
@(posedge clk_i);
a_mant0 = 8'd68; a_mant1 = 8'd146; a_mant2 = 8'd47; a_mant3 = 8'd209;
b_mant0 = 8'd196; b_mant1 = 8'd114; b_mant2 = 8'd238; b_mant3 = 8'd86;
a_exp0 = 10'd146; a_exp1 = 10'd967; a_exp2 = 10'd860; a_exp3 = 10'd688;
b_exp0 = 10'd875; b_exp1 = 10'd956; b_exp2 = 10'd970; b_exp3 = 10'd272;
a_sign0 = 4'd0; a_sign1 = 4'd6; a_sign2 = 4'd4; a_sign3 = 4'd5;
b_sign0 = 4'd7; b_sign1 = 4'd4; b_sign2 = 4'd1; b_sign3 = 4'd2;
@(posedge clk_i);
a_mant0 = 8'd209; a_mant1 = 8'd71; a_mant2 = 8'd206; a_mant3 = 8'd96;
b_mant0 = 8'd129; b_mant1 = 8'd10; b_mant2 = 8'd83; b_mant3 = 8'd141;
a_exp0 = 10'd0; a_exp1 = 10'd562; a_exp2 = 10'd502; a_exp3 = 10'd329;
b_exp0 = 10'd715; b_exp1 = 10'd27; b_exp2 = 10'd249; b_exp3 = 10'd846;
a_sign0 = 4'd16; a_sign1 = 4'd3; a_sign2 = 4'd3; a_sign3 = 4'd0;
b_sign0 = 4'd3; b_sign1 = 4'd8; b_sign2 = 4'd8; b_sign3 = 4'd13;
@(posedge clk_i);
a_mant0 = 8'd201; a_mant1 = 8'd211; a_mant2 = 8'd39; a_mant3 = 8'd162;
b_mant0 = 8'd248; b_mant1 = 8'd234; b_mant2 = 8'd159; b_mant3 = 8'd176;
a_exp0 = 10'd581; a_exp1 = 10'd459; a_exp2 = 10'd72; a_exp3 = 10'd454;
b_exp0 = 10'd345; b_exp1 = 10'd1006; b_exp2 = 10'd50; b_exp3 = 10'd277;
a_sign0 = 4'd14; a_sign1 = 4'd8; a_sign2 = 4'd13; a_sign3 = 4'd1;
b_sign0 = 4'd14; b_sign1 = 4'd1; b_sign2 = 4'd15; b_sign3 = 4'd15;
@(posedge clk_i);
a_mant0 = 8'd99; a_mant1 = 8'd119; a_mant2 = 8'd90; a_mant3 = 8'd160;
b_mant0 = 8'd139; b_mant1 = 8'd5; b_mant2 = 8'd32; b_mant3 = 8'd229;
a_exp0 = 10'd462; a_exp1 = 10'd0; a_exp2 = 10'd758; a_exp3 = 10'd147;
b_exp0 = 10'd949; b_exp1 = 10'd886; b_exp2 = 10'd411; b_exp3 = 10'd556;
a_sign0 = 4'd15; a_sign1 = 4'd10; a_sign2 = 4'd15; a_sign3 = 4'd12;
b_sign0 = 4'd3; b_sign1 = 4'd3; b_sign2 = 4'd1; b_sign3 = 4'd7;
@(posedge clk_i);
a_mant0 = 8'd77; a_mant1 = 8'd17; a_mant2 = 8'd149; a_mant3 = 8'd206;
b_mant0 = 8'd67; b_mant1 = 8'd192; b_mant2 = 8'd195; b_mant3 = 8'd206;
a_exp0 = 10'd534; a_exp1 = 10'd268; a_exp2 = 10'd548; a_exp3 = 10'd953;
b_exp0 = 10'd323; b_exp1 = 10'd506; b_exp2 = 10'd706; b_exp3 = 10'd808;
a_sign0 = 4'd12; a_sign1 = 4'd14; a_sign2 = 4'd12; a_sign3 = 4'd5;
b_sign0 = 4'd13; b_sign1 = 4'd12; b_sign2 = 4'd13; b_sign3 = 4'd12;
@(posedge clk_i);
a_mant0 = 8'd204; a_mant1 = 8'd203; a_mant2 = 8'd69; a_mant3 = 8'd0;
b_mant0 = 8'd1; b_mant1 = 8'd21; b_mant2 = 8'd33; b_mant3 = 8'd199;
a_exp0 = 10'd142; a_exp1 = 10'd852; a_exp2 = 10'd711; a_exp3 = 10'd910;
b_exp0 = 10'd140; b_exp1 = 10'd370; b_exp2 = 10'd930; b_exp3 = 10'd854;
a_sign0 = 4'd4; a_sign1 = 4'd15; a_sign2 = 4'd0; a_sign3 = 4'd15;
b_sign0 = 4'd1; b_sign1 = 4'd5; b_sign2 = 4'd0; b_sign3 = 4'd0;
@(posedge clk_i);
shared_exps0 = 8'd131;
shared_exps1 = 8'd137;
rstn = 0;
@(posedge clk_i);
rstn = 1;
a_mant0 = 8'd101; a_mant1 = 8'd118; a_mant2 = 8'd120; a_mant3 = 8'd111;
b_mant0 = 8'd17; b_mant1 = 8'd198; b_mant2 = 8'd0; b_mant3 = 8'd222;
a_exp0 = 10'd672; a_exp1 = 10'd849; a_exp2 = 10'd378; a_exp3 = 10'd960;
b_exp0 = 10'd959; b_exp1 = 10'd145; b_exp2 = 10'd161; b_exp3 = 10'd250;
a_sign0 = 4'd2; a_sign1 = 4'd11; a_sign2 = 4'd11; a_sign3 = 4'd4;
b_sign0 = 4'd4; b_sign1 = 4'd3; b_sign2 = 4'd0; b_sign3 = 4'd11;
@(posedge clk_i);
a_mant0 = 8'd85; a_mant1 = 8'd240; a_mant2 = 8'd113; a_mant3 = 8'd201;
b_mant0 = 8'd68; b_mant1 = 8'd173; b_mant2 = 8'd238; b_mant3 = 8'd29;
a_exp0 = 10'd890; a_exp1 = 10'd844; a_exp2 = 10'd650; a_exp3 = 10'd449;
b_exp0 = 10'd691; b_exp1 = 10'd511; b_exp2 = 10'd837; b_exp3 = 10'd742;
a_sign0 = 4'd6; a_sign1 = 4'd2; a_sign2 = 4'd16; a_sign3 = 4'd2;
b_sign0 = 4'd1; b_sign1 = 4'd12; b_sign2 = 4'd15; b_sign3 = 4'd2;
@(posedge clk_i);
a_mant0 = 8'd16; a_mant1 = 8'd145; a_mant2 = 8'd61; a_mant3 = 8'd70;
b_mant0 = 8'd24; b_mant1 = 8'd157; b_mant2 = 8'd53; b_mant3 = 8'd114;
a_exp0 = 10'd19; a_exp1 = 10'd883; a_exp2 = 10'd675; a_exp3 = 10'd18;
b_exp0 = 10'd46; b_exp1 = 10'd688; b_exp2 = 10'd408; b_exp3 = 10'd37;
a_sign0 = 4'd15; a_sign1 = 4'd10; a_sign2 = 4'd11; a_sign3 = 4'd16;
b_sign0 = 4'd13; b_sign1 = 4'd10; b_sign2 = 4'd11; b_sign3 = 4'd1;
@(posedge clk_i);
a_mant0 = 8'd193; a_mant1 = 8'd216; a_mant2 = 8'd114; a_mant3 = 8'd67;
b_mant0 = 8'd228; b_mant1 = 8'd168; b_mant2 = 8'd121; b_mant3 = 8'd228;
a_exp0 = 10'd744; a_exp1 = 10'd303; a_exp2 = 10'd647; a_exp3 = 10'd981;
b_exp0 = 10'd38; b_exp1 = 10'd203; b_exp2 = 10'd111; b_exp3 = 10'd732;
a_sign0 = 4'd2; a_sign1 = 4'd1; a_sign2 = 4'd0; a_sign3 = 4'd6;
b_sign0 = 4'd15; b_sign1 = 4'd5; b_sign2 = 4'd9; b_sign3 = 4'd14;
@(posedge clk_i);
a_mant0 = 8'd198; a_mant1 = 8'd202; a_mant2 = 8'd247; a_mant3 = 8'd221;
b_mant0 = 8'd93; b_mant1 = 8'd219; b_mant2 = 8'd178; b_mant3 = 8'd168;
a_exp0 = 10'd612; a_exp1 = 10'd908; a_exp2 = 10'd877; a_exp3 = 10'd254;
b_exp0 = 10'd504; b_exp1 = 10'd492; b_exp2 = 10'd20; b_exp3 = 10'd959;
a_sign0 = 4'd15; a_sign1 = 4'd11; a_sign2 = 4'd13; a_sign3 = 4'd15;
b_sign0 = 4'd12; b_sign1 = 4'd9; b_sign2 = 4'd0; b_sign3 = 4'd4;
@(posedge clk_i);
a_mant0 = 8'd161; a_mant1 = 8'd74; a_mant2 = 8'd224; a_mant3 = 8'd222;
b_mant0 = 8'd221; b_mant1 = 8'd47; b_mant2 = 8'd131; b_mant3 = 8'd224;
a_exp0 = 10'd852; a_exp1 = 10'd115; a_exp2 = 10'd626; a_exp3 = 10'd57;
b_exp0 = 10'd235; b_exp1 = 10'd224; b_exp2 = 10'd129; b_exp3 = 10'd150;
a_sign0 = 4'd12; a_sign1 = 4'd15; a_sign2 = 4'd16; a_sign3 = 4'd2;
b_sign0 = 4'd5; b_sign1 = 4'd11; b_sign2 = 4'd8; b_sign3 = 4'd7;
@(posedge clk_i);
a_mant0 = 8'd16; a_mant1 = 8'd222; a_mant2 = 8'd208; a_mant3 = 8'd210;
b_mant0 = 8'd92; b_mant1 = 8'd63; b_mant2 = 8'd95; b_mant3 = 8'd161;
a_exp0 = 10'd85; a_exp1 = 10'd812; a_exp2 = 10'd759; a_exp3 = 10'd1019;
b_exp0 = 10'd557; b_exp1 = 10'd974; b_exp2 = 10'd294; b_exp3 = 10'd804;
a_sign0 = 4'd2; a_sign1 = 4'd5; a_sign2 = 4'd2; a_sign3 = 4'd9;
b_sign0 = 4'd9; b_sign1 = 4'd16; b_sign2 = 4'd5; b_sign3 = 4'd8;
@(posedge clk_i);
shared_exps0 = 8'd134;
shared_exps1 = 8'd132;
a_mant0 = 8'd100; a_mant1 = 8'd19; a_mant2 = 8'd78; a_mant3 = 8'd255;
b_mant0 = 8'd252; b_mant1 = 8'd14; b_mant2 = 8'd153; b_mant3 = 8'd58;
a_exp0 = 10'd808; a_exp1 = 10'd955; a_exp2 = 10'd997; a_exp3 = 10'd809;
b_exp0 = 10'd62; b_exp1 = 10'd340; b_exp2 = 10'd1002; b_exp3 = 10'd969;
a_sign0 = 4'd4; a_sign1 = 4'd5; a_sign2 = 4'd0; a_sign3 = 4'd13;
b_sign0 = 4'd15; b_sign1 = 4'd3; b_sign2 = 4'd12; b_sign3 = 4'd5;
@(posedge clk_i);
a_mant0 = 8'd236; a_mant1 = 8'd101; a_mant2 = 8'd55; a_mant3 = 8'd80;
b_mant0 = 8'd32; b_mant1 = 8'd203; b_mant2 = 8'd251; b_mant3 = 8'd58;
a_exp0 = 10'd344; a_exp1 = 10'd526; a_exp2 = 10'd1006; a_exp3 = 10'd886;
b_exp0 = 10'd629; b_exp1 = 10'd537; b_exp2 = 10'd305; b_exp3 = 10'd252;
a_sign0 = 4'd3; a_sign1 = 4'd16; a_sign2 = 4'd4; a_sign3 = 4'd4;
b_sign0 = 4'd13; b_sign1 = 4'd16; b_sign2 = 4'd3; b_sign3 = 4'd1;
@(posedge clk_i);
a_mant0 = 8'd189; a_mant1 = 8'd39; a_mant2 = 8'd222; a_mant3 = 8'd32;
b_mant0 = 8'd247; b_mant1 = 8'd114; b_mant2 = 8'd73; b_mant3 = 8'd176;
a_exp0 = 10'd276; a_exp1 = 10'd754; a_exp2 = 10'd396; a_exp3 = 10'd1022;
b_exp0 = 10'd474; b_exp1 = 10'd415; b_exp2 = 10'd184; b_exp3 = 10'd45;
a_sign0 = 4'd4; a_sign1 = 4'd1; a_sign2 = 4'd16; a_sign3 = 4'd8;
b_sign0 = 4'd1; b_sign1 = 4'd15; b_sign2 = 4'd6; b_sign3 = 4'd4;
@(posedge clk_i);
a_mant0 = 8'd126; a_mant1 = 8'd225; a_mant2 = 8'd229; a_mant3 = 8'd31;
b_mant0 = 8'd61; b_mant1 = 8'd173; b_mant2 = 8'd238; b_mant3 = 8'd78;
a_exp0 = 10'd235; a_exp1 = 10'd110; a_exp2 = 10'd1010; a_exp3 = 10'd250;
b_exp0 = 10'd244; b_exp1 = 10'd658; b_exp2 = 10'd646; b_exp3 = 10'd374;
a_sign0 = 4'd3; a_sign1 = 4'd9; a_sign2 = 4'd0; a_sign3 = 4'd10;
b_sign0 = 4'd10; b_sign1 = 4'd14; b_sign2 = 4'd1; b_sign3 = 4'd7;
@(posedge clk_i);
a_mant0 = 8'd219; a_mant1 = 8'd251; a_mant2 = 8'd23; a_mant3 = 8'd8;
b_mant0 = 8'd50; b_mant1 = 8'd85; b_mant2 = 8'd171; b_mant3 = 8'd6;
a_exp0 = 10'd993; a_exp1 = 10'd448; a_exp2 = 10'd70; a_exp3 = 10'd431;
b_exp0 = 10'd636; b_exp1 = 10'd949; b_exp2 = 10'd639; b_exp3 = 10'd240;
a_sign0 = 4'd4; a_sign1 = 4'd2; a_sign2 = 4'd0; a_sign3 = 4'd13;
b_sign0 = 4'd11; b_sign1 = 4'd5; b_sign2 = 4'd8; b_sign3 = 4'd8;
@(posedge clk_i);
a_mant0 = 8'd17; a_mant1 = 8'd255; a_mant2 = 8'd181; a_mant3 = 8'd177;
b_mant0 = 8'd3; b_mant1 = 8'd20; b_mant2 = 8'd158; b_mant3 = 8'd5;
a_exp0 = 10'd926; a_exp1 = 10'd865; a_exp2 = 10'd911; a_exp3 = 10'd289;
b_exp0 = 10'd235; b_exp1 = 10'd994; b_exp2 = 10'd396; b_exp3 = 10'd875;
a_sign0 = 4'd3; a_sign1 = 4'd1; a_sign2 = 4'd4; a_sign3 = 4'd9;
b_sign0 = 4'd15; b_sign1 = 4'd16; b_sign2 = 4'd14; b_sign3 = 4'd3;
@(posedge clk_i);
a_mant0 = 8'd16; a_mant1 = 8'd152; a_mant2 = 8'd190; a_mant3 = 8'd32;
b_mant0 = 8'd54; b_mant1 = 8'd78; b_mant2 = 8'd125; b_mant3 = 8'd90;
a_exp0 = 10'd1; a_exp1 = 10'd359; a_exp2 = 10'd213; a_exp3 = 10'd796;
b_exp0 = 10'd486; b_exp1 = 10'd1022; b_exp2 = 10'd293; b_exp3 = 10'd675;
a_sign0 = 4'd12; a_sign1 = 4'd8; a_sign2 = 4'd12; a_sign3 = 4'd11;
b_sign0 = 4'd10; b_sign1 = 4'd14; b_sign2 = 4'd15; b_sign3 = 4'd6;
@(posedge clk_i);
a_mant0 = 8'd72; a_mant1 = 8'd148; a_mant2 = 8'd188; a_mant3 = 8'd211;
b_mant0 = 8'd192; b_mant1 = 8'd199; b_mant2 = 8'd250; b_mant3 = 8'd20;
a_exp0 = 10'd264; a_exp1 = 10'd4; a_exp2 = 10'd824; a_exp3 = 10'd529;
b_exp0 = 10'd259; b_exp1 = 10'd937; b_exp2 = 10'd923; b_exp3 = 10'd393;
a_sign0 = 4'd2; a_sign1 = 4'd0; a_sign2 = 4'd7; a_sign3 = 4'd8;
b_sign0 = 4'd14; b_sign1 = 4'd11; b_sign2 = 4'd8; b_sign3 = 4'd12;
@(posedge clk_i);
shared_exps0 = 8'd120;
shared_exps1 = 8'd155;
a_mant0 = 8'd215; a_mant1 = 8'd216; a_mant2 = 8'd179; a_mant3 = 8'd134;
b_mant0 = 8'd97; b_mant1 = 8'd185; b_mant2 = 8'd9; b_mant3 = 8'd24;
a_exp0 = 10'd40; a_exp1 = 10'd454; a_exp2 = 10'd722; a_exp3 = 10'd414;
b_exp0 = 10'd129; b_exp1 = 10'd82; b_exp2 = 10'd535; b_exp3 = 10'd521;
a_sign0 = 4'd16; a_sign1 = 4'd6; a_sign2 = 4'd15; a_sign3 = 4'd12;
b_sign0 = 4'd3; b_sign1 = 4'd2; b_sign2 = 4'd16; b_sign3 = 4'd14;
@(posedge clk_i);
a_mant0 = 8'd93; a_mant1 = 8'd67; a_mant2 = 8'd88; a_mant3 = 8'd33;
b_mant0 = 8'd105; b_mant1 = 8'd237; b_mant2 = 8'd50; b_mant3 = 8'd178;
a_exp0 = 10'd575; a_exp1 = 10'd615; a_exp2 = 10'd658; a_exp3 = 10'd683;
b_exp0 = 10'd430; b_exp1 = 10'd195; b_exp2 = 10'd758; b_exp3 = 10'd286;
a_sign0 = 4'd0; a_sign1 = 4'd10; a_sign2 = 4'd11; a_sign3 = 4'd11;
b_sign0 = 4'd3; b_sign1 = 4'd6; b_sign2 = 4'd14; b_sign3 = 4'd11;
@(posedge clk_i);
a_mant0 = 8'd102; a_mant1 = 8'd168; a_mant2 = 8'd167; a_mant3 = 8'd85;
b_mant0 = 8'd99; b_mant1 = 8'd145; b_mant2 = 8'd189; b_mant3 = 8'd107;
a_exp0 = 10'd901; a_exp1 = 10'd973; a_exp2 = 10'd318; a_exp3 = 10'd280;
b_exp0 = 10'd293; b_exp1 = 10'd573; b_exp2 = 10'd945; b_exp3 = 10'd818;
a_sign0 = 4'd15; a_sign1 = 4'd10; a_sign2 = 4'd7; a_sign3 = 4'd16;
b_sign0 = 4'd3; b_sign1 = 4'd1; b_sign2 = 4'd1; b_sign3 = 4'd6;
@(posedge clk_i);
a_mant0 = 8'd185; a_mant1 = 8'd225; a_mant2 = 8'd241; a_mant3 = 8'd221;
b_mant0 = 8'd201; b_mant1 = 8'd216; b_mant2 = 8'd27; b_mant3 = 8'd184;
a_exp0 = 10'd742; a_exp1 = 10'd517; a_exp2 = 10'd779; a_exp3 = 10'd423;
b_exp0 = 10'd585; b_exp1 = 10'd864; b_exp2 = 10'd874; b_exp3 = 10'd311;
a_sign0 = 4'd9; a_sign1 = 4'd0; a_sign2 = 4'd14; a_sign3 = 4'd3;
b_sign0 = 4'd16; b_sign1 = 4'd9; b_sign2 = 4'd2; b_sign3 = 4'd4;
@(posedge clk_i);
a_mant0 = 8'd97; a_mant1 = 8'd244; a_mant2 = 8'd106; a_mant3 = 8'd131;
b_mant0 = 8'd46; b_mant1 = 8'd154; b_mant2 = 8'd162; b_mant3 = 8'd143;
a_exp0 = 10'd901; a_exp1 = 10'd499; a_exp2 = 10'd792; a_exp3 = 10'd54;
b_exp0 = 10'd478; b_exp1 = 10'd768; b_exp2 = 10'd824; b_exp3 = 10'd590;
a_sign0 = 4'd11; a_sign1 = 4'd8; a_sign2 = 4'd7; a_sign3 = 4'd6;
b_sign0 = 4'd13; b_sign1 = 4'd12; b_sign2 = 4'd3; b_sign3 = 4'd14;
@(posedge clk_i);
a_mant0 = 8'd73; a_mant1 = 8'd232; a_mant2 = 8'd93; a_mant3 = 8'd192;
b_mant0 = 8'd165; b_mant1 = 8'd225; b_mant2 = 8'd155; b_mant3 = 8'd11;
a_exp0 = 10'd317; a_exp1 = 10'd99; a_exp2 = 10'd215; a_exp3 = 10'd606;
b_exp0 = 10'd918; b_exp1 = 10'd240; b_exp2 = 10'd157; b_exp3 = 10'd297;
a_sign0 = 4'd15; a_sign1 = 4'd3; a_sign2 = 4'd4; a_sign3 = 4'd16;
b_sign0 = 4'd14; b_sign1 = 4'd16; b_sign2 = 4'd3; b_sign3 = 4'd7;
@(posedge clk_i);
a_mant0 = 8'd158; a_mant1 = 8'd107; a_mant2 = 8'd180; a_mant3 = 8'd217;
b_mant0 = 8'd218; b_mant1 = 8'd231; b_mant2 = 8'd8; b_mant3 = 8'd240;
a_exp0 = 10'd521; a_exp1 = 10'd111; a_exp2 = 10'd244; a_exp3 = 10'd527;
b_exp0 = 10'd193; b_exp1 = 10'd709; b_exp2 = 10'd154; b_exp3 = 10'd375;
a_sign0 = 4'd7; a_sign1 = 4'd13; a_sign2 = 4'd12; a_sign3 = 4'd12;
b_sign0 = 4'd4; b_sign1 = 4'd16; b_sign2 = 4'd9; b_sign3 = 4'd16;
@(posedge clk_i);
a_mant0 = 8'd178; a_mant1 = 8'd171; a_mant2 = 8'd45; a_mant3 = 8'd165;
b_mant0 = 8'd21; b_mant1 = 8'd201; b_mant2 = 8'd56; b_mant3 = 8'd30;
a_exp0 = 10'd701; a_exp1 = 10'd86; a_exp2 = 10'd528; a_exp3 = 10'd549;
b_exp0 = 10'd979; b_exp1 = 10'd1014; b_exp2 = 10'd801; b_exp3 = 10'd895;
a_sign0 = 4'd11; a_sign1 = 4'd7; a_sign2 = 4'd9; a_sign3 = 4'd11;
b_sign0 = 4'd0; b_sign1 = 4'd2; b_sign2 = 4'd0; b_sign3 = 4'd6;
@(posedge clk_i);
shared_exps0 = 8'd108;
shared_exps1 = 8'd82;
a_mant0 = 8'd72; a_mant1 = 8'd9; a_mant2 = 8'd171; a_mant3 = 8'd152;
b_mant0 = 8'd185; b_mant1 = 8'd232; b_mant2 = 8'd196; b_mant3 = 8'd235;
a_exp0 = 10'd589; a_exp1 = 10'd109; a_exp2 = 10'd830; a_exp3 = 10'd806;
b_exp0 = 10'd308; b_exp1 = 10'd173; b_exp2 = 10'd550; b_exp3 = 10'd452;
a_sign0 = 4'd9; a_sign1 = 4'd5; a_sign2 = 4'd9; a_sign3 = 4'd5;
b_sign0 = 4'd13; b_sign1 = 4'd0; b_sign2 = 4'd10; b_sign3 = 4'd10;
@(posedge clk_i);
a_mant0 = 8'd164; a_mant1 = 8'd216; a_mant2 = 8'd139; a_mant3 = 8'd0;
b_mant0 = 8'd99; b_mant1 = 8'd162; b_mant2 = 8'd45; b_mant3 = 8'd159;
a_exp0 = 10'd694; a_exp1 = 10'd504; a_exp2 = 10'd838; a_exp3 = 10'd390;
b_exp0 = 10'd379; b_exp1 = 10'd982; b_exp2 = 10'd507; b_exp3 = 10'd459;
a_sign0 = 4'd9; a_sign1 = 4'd4; a_sign2 = 4'd11; a_sign3 = 4'd5;
b_sign0 = 4'd14; b_sign1 = 4'd11; b_sign2 = 4'd16; b_sign3 = 4'd1;
@(posedge clk_i);
a_mant0 = 8'd142; a_mant1 = 8'd42; a_mant2 = 8'd230; a_mant3 = 8'd197;
b_mant0 = 8'd16; b_mant1 = 8'd213; b_mant2 = 8'd28; b_mant3 = 8'd86;
a_exp0 = 10'd137; a_exp1 = 10'd959; a_exp2 = 10'd846; a_exp3 = 10'd628;
b_exp0 = 10'd667; b_exp1 = 10'd853; b_exp2 = 10'd443; b_exp3 = 10'd678;
a_sign0 = 4'd5; a_sign1 = 4'd0; a_sign2 = 4'd7; a_sign3 = 4'd1;
b_sign0 = 4'd3; b_sign1 = 4'd8; b_sign2 = 4'd8; b_sign3 = 4'd7;
@(posedge clk_i);
a_mant0 = 8'd201; a_mant1 = 8'd86; a_mant2 = 8'd102; a_mant3 = 8'd206;
b_mant0 = 8'd158; b_mant1 = 8'd170; b_mant2 = 8'd119; b_mant3 = 8'd225;
a_exp0 = 10'd681; a_exp1 = 10'd39; a_exp2 = 10'd240; a_exp3 = 10'd996;
b_exp0 = 10'd469; b_exp1 = 10'd527; b_exp2 = 10'd870; b_exp3 = 10'd512;
a_sign0 = 4'd16; a_sign1 = 4'd15; a_sign2 = 4'd6; a_sign3 = 4'd12;
b_sign0 = 4'd7; b_sign1 = 4'd11; b_sign2 = 4'd4; b_sign3 = 4'd12;
@(posedge clk_i);
a_mant0 = 8'd202; a_mant1 = 8'd1; a_mant2 = 8'd161; a_mant3 = 8'd239;
b_mant0 = 8'd183; b_mant1 = 8'd119; b_mant2 = 8'd129; b_mant3 = 8'd51;
a_exp0 = 10'd953; a_exp1 = 10'd492; a_exp2 = 10'd743; a_exp3 = 10'd744;
b_exp0 = 10'd402; b_exp1 = 10'd34; b_exp2 = 10'd197; b_exp3 = 10'd707;
a_sign0 = 4'd14; a_sign1 = 4'd10; a_sign2 = 4'd8; a_sign3 = 4'd0;
b_sign0 = 4'd4; b_sign1 = 4'd0; b_sign2 = 4'd3; b_sign3 = 4'd2;
@(posedge clk_i);
a_mant0 = 8'd222; a_mant1 = 8'd136; a_mant2 = 8'd109; a_mant3 = 8'd88;
b_mant0 = 8'd93; b_mant1 = 8'd161; b_mant2 = 8'd249; b_mant3 = 8'd104;
a_exp0 = 10'd317; a_exp1 = 10'd998; a_exp2 = 10'd136; a_exp3 = 10'd33;
b_exp0 = 10'd702; b_exp1 = 10'd710; b_exp2 = 10'd229; b_exp3 = 10'd386;
a_sign0 = 4'd15; a_sign1 = 4'd13; a_sign2 = 4'd14; a_sign3 = 4'd12;
b_sign0 = 4'd3; b_sign1 = 4'd15; b_sign2 = 4'd0; b_sign3 = 4'd13;
@(posedge clk_i);
a_mant0 = 8'd179; a_mant1 = 8'd94; a_mant2 = 8'd69; a_mant3 = 8'd105;
b_mant0 = 8'd186; b_mant1 = 8'd219; b_mant2 = 8'd10; b_mant3 = 8'd252;
a_exp0 = 10'd101; a_exp1 = 10'd482; a_exp2 = 10'd208; a_exp3 = 10'd834;
b_exp0 = 10'd418; b_exp1 = 10'd34; b_exp2 = 10'd116; b_exp3 = 10'd570;
a_sign0 = 4'd12; a_sign1 = 4'd6; a_sign2 = 4'd4; a_sign3 = 4'd12;
b_sign0 = 4'd7; b_sign1 = 4'd15; b_sign2 = 4'd5; b_sign3 = 4'd13;
@(posedge clk_i);
a_mant0 = 8'd129; a_mant1 = 8'd249; a_mant2 = 8'd30; a_mant3 = 8'd96;
b_mant0 = 8'd151; b_mant1 = 8'd133; b_mant2 = 8'd45; b_mant3 = 8'd228;
a_exp0 = 10'd590; a_exp1 = 10'd785; a_exp2 = 10'd614; a_exp3 = 10'd526;
b_exp0 = 10'd276; b_exp1 = 10'd1003; b_exp2 = 10'd397; b_exp3 = 10'd317;
a_sign0 = 4'd9; a_sign1 = 4'd12; a_sign2 = 4'd4; a_sign3 = 4'd5;
b_sign0 = 4'd11; b_sign1 = 4'd4; b_sign2 = 4'd7; b_sign3 = 4'd16;
@(posedge clk_i);
shared_exps0 = 8'd127;
shared_exps1 = 8'd119;
rstn = 0;
@(posedge clk_i);
rstn = 1;
a_mant0 = 8'd63; a_mant1 = 8'd125; a_mant2 = 8'd121; a_mant3 = 8'd102;
b_mant0 = 8'd218; b_mant1 = 8'd101; b_mant2 = 8'd119; b_mant3 = 8'd38;
a_exp0 = 10'd385; a_exp1 = 10'd373; a_exp2 = 10'd121; a_exp3 = 10'd426;
b_exp0 = 10'd406; b_exp1 = 10'd272; b_exp2 = 10'd882; b_exp3 = 10'd233;
a_sign0 = 4'd11; a_sign1 = 4'd13; a_sign2 = 4'd16; a_sign3 = 4'd7;
b_sign0 = 4'd7; b_sign1 = 4'd3; b_sign2 = 4'd5; b_sign3 = 4'd12;
@(posedge clk_i);
a_mant0 = 8'd181; a_mant1 = 8'd7; a_mant2 = 8'd176; a_mant3 = 8'd90;
b_mant0 = 8'd61; b_mant1 = 8'd164; b_mant2 = 8'd179; b_mant3 = 8'd169;
a_exp0 = 10'd885; a_exp1 = 10'd446; a_exp2 = 10'd54; a_exp3 = 10'd670;
b_exp0 = 10'd375; b_exp1 = 10'd80; b_exp2 = 10'd832; b_exp3 = 10'd645;
a_sign0 = 4'd0; a_sign1 = 4'd10; a_sign2 = 4'd12; a_sign3 = 4'd2;
b_sign0 = 4'd2; b_sign1 = 4'd3; b_sign2 = 4'd13; b_sign3 = 4'd4;
@(posedge clk_i);
a_mant0 = 8'd187; a_mant1 = 8'd159; a_mant2 = 8'd114; a_mant3 = 8'd0;
b_mant0 = 8'd167; b_mant1 = 8'd153; b_mant2 = 8'd129; b_mant3 = 8'd248;
a_exp0 = 10'd481; a_exp1 = 10'd943; a_exp2 = 10'd341; a_exp3 = 10'd825;
b_exp0 = 10'd1; b_exp1 = 10'd962; b_exp2 = 10'd560; b_exp3 = 10'd938;
a_sign0 = 4'd13; a_sign1 = 4'd1; a_sign2 = 4'd6; a_sign3 = 4'd6;
b_sign0 = 4'd10; b_sign1 = 4'd13; b_sign2 = 4'd14; b_sign3 = 4'd10;
@(posedge clk_i);
a_mant0 = 8'd122; a_mant1 = 8'd95; a_mant2 = 8'd94; a_mant3 = 8'd34;
b_mant0 = 8'd142; b_mant1 = 8'd64; b_mant2 = 8'd236; b_mant3 = 8'd177;
a_exp0 = 10'd87; a_exp1 = 10'd48; a_exp2 = 10'd825; a_exp3 = 10'd878;
b_exp0 = 10'd431; b_exp1 = 10'd440; b_exp2 = 10'd453; b_exp3 = 10'd426;
a_sign0 = 4'd0; a_sign1 = 4'd12; a_sign2 = 4'd2; a_sign3 = 4'd9;
b_sign0 = 4'd16; b_sign1 = 4'd12; b_sign2 = 4'd8; b_sign3 = 4'd4;
@(posedge clk_i);
a_mant0 = 8'd188; a_mant1 = 8'd45; a_mant2 = 8'd86; a_mant3 = 8'd197;
b_mant0 = 8'd204; b_mant1 = 8'd190; b_mant2 = 8'd59; b_mant3 = 8'd38;
a_exp0 = 10'd976; a_exp1 = 10'd845; a_exp2 = 10'd950; a_exp3 = 10'd645;
b_exp0 = 10'd84; b_exp1 = 10'd851; b_exp2 = 10'd509; b_exp3 = 10'd323;
a_sign0 = 4'd11; a_sign1 = 4'd5; a_sign2 = 4'd1; a_sign3 = 4'd15;
b_sign0 = 4'd12; b_sign1 = 4'd8; b_sign2 = 4'd13; b_sign3 = 4'd12;
@(posedge clk_i);
a_mant0 = 8'd147; a_mant1 = 8'd234; a_mant2 = 8'd235; a_mant3 = 8'd11;
b_mant0 = 8'd223; b_mant1 = 8'd194; b_mant2 = 8'd20; b_mant3 = 8'd158;
a_exp0 = 10'd560; a_exp1 = 10'd334; a_exp2 = 10'd240; a_exp3 = 10'd287;
b_exp0 = 10'd704; b_exp1 = 10'd413; b_exp2 = 10'd391; b_exp3 = 10'd356;
a_sign0 = 4'd7; a_sign1 = 4'd15; a_sign2 = 4'd5; a_sign3 = 4'd5;
b_sign0 = 4'd12; b_sign1 = 4'd7; b_sign2 = 4'd16; b_sign3 = 4'd8;
@(posedge clk_i);
a_mant0 = 8'd198; a_mant1 = 8'd4; a_mant2 = 8'd141; a_mant3 = 8'd119;
b_mant0 = 8'd155; b_mant1 = 8'd38; b_mant2 = 8'd135; b_mant3 = 8'd45;
a_exp0 = 10'd834; a_exp1 = 10'd280; a_exp2 = 10'd132; a_exp3 = 10'd56;
b_exp0 = 10'd429; b_exp1 = 10'd537; b_exp2 = 10'd930; b_exp3 = 10'd163;
a_sign0 = 4'd10; a_sign1 = 4'd3; a_sign2 = 4'd15; a_sign3 = 4'd13;
b_sign0 = 4'd9; b_sign1 = 4'd13; b_sign2 = 4'd8; b_sign3 = 4'd15;
@(posedge clk_i);
shared_exps0 = 8'd115;
shared_exps1 = 8'd119;
a_mant0 = 8'd54; a_mant1 = 8'd117; a_mant2 = 8'd5; a_mant3 = 8'd206;
b_mant0 = 8'd179; b_mant1 = 8'd149; b_mant2 = 8'd216; b_mant3 = 8'd114;
a_exp0 = 10'd7; a_exp1 = 10'd213; a_exp2 = 10'd976; a_exp3 = 10'd402;
b_exp0 = 10'd232; b_exp1 = 10'd858; b_exp2 = 10'd828; b_exp3 = 10'd603;
a_sign0 = 4'd4; a_sign1 = 4'd16; a_sign2 = 4'd11; a_sign3 = 4'd15;
b_sign0 = 4'd16; b_sign1 = 4'd1; b_sign2 = 4'd6; b_sign3 = 4'd9;
@(posedge clk_i);
a_mant0 = 8'd196; a_mant1 = 8'd26; a_mant2 = 8'd61; a_mant3 = 8'd187;
b_mant0 = 8'd185; b_mant1 = 8'd39; b_mant2 = 8'd47; b_mant3 = 8'd169;
a_exp0 = 10'd131; a_exp1 = 10'd769; a_exp2 = 10'd59; a_exp3 = 10'd260;
b_exp0 = 10'd176; b_exp1 = 10'd685; b_exp2 = 10'd685; b_exp3 = 10'd872;
a_sign0 = 4'd4; a_sign1 = 4'd8; a_sign2 = 4'd13; a_sign3 = 4'd12;
b_sign0 = 4'd14; b_sign1 = 4'd6; b_sign2 = 4'd11; b_sign3 = 4'd12;
@(posedge clk_i);
a_mant0 = 8'd254; a_mant1 = 8'd107; a_mant2 = 8'd23; a_mant3 = 8'd229;
b_mant0 = 8'd58; b_mant1 = 8'd230; b_mant2 = 8'd137; b_mant3 = 8'd248;
a_exp0 = 10'd386; a_exp1 = 10'd213; a_exp2 = 10'd129; a_exp3 = 10'd135;
b_exp0 = 10'd424; b_exp1 = 10'd906; b_exp2 = 10'd646; b_exp3 = 10'd657;
a_sign0 = 4'd0; a_sign1 = 4'd3; a_sign2 = 4'd11; a_sign3 = 4'd5;
b_sign0 = 4'd6; b_sign1 = 4'd16; b_sign2 = 4'd8; b_sign3 = 4'd11;
@(posedge clk_i);
a_mant0 = 8'd65; a_mant1 = 8'd9; a_mant2 = 8'd215; a_mant3 = 8'd137;
b_mant0 = 8'd149; b_mant1 = 8'd117; b_mant2 = 8'd177; b_mant3 = 8'd37;
a_exp0 = 10'd883; a_exp1 = 10'd230; a_exp2 = 10'd523; a_exp3 = 10'd931;
b_exp0 = 10'd184; b_exp1 = 10'd263; b_exp2 = 10'd630; b_exp3 = 10'd425;
a_sign0 = 4'd6; a_sign1 = 4'd5; a_sign2 = 4'd4; a_sign3 = 4'd11;
b_sign0 = 4'd12; b_sign1 = 4'd8; b_sign2 = 4'd14; b_sign3 = 4'd0;
@(posedge clk_i);
a_mant0 = 8'd72; a_mant1 = 8'd209; a_mant2 = 8'd15; a_mant3 = 8'd138;
b_mant0 = 8'd19; b_mant1 = 8'd248; b_mant2 = 8'd251; b_mant3 = 8'd52;
a_exp0 = 10'd319; a_exp1 = 10'd686; a_exp2 = 10'd849; a_exp3 = 10'd727;
b_exp0 = 10'd249; b_exp1 = 10'd356; b_exp2 = 10'd978; b_exp3 = 10'd969;
a_sign0 = 4'd5; a_sign1 = 4'd11; a_sign2 = 4'd7; a_sign3 = 4'd15;
b_sign0 = 4'd6; b_sign1 = 4'd15; b_sign2 = 4'd3; b_sign3 = 4'd12;
@(posedge clk_i);
a_mant0 = 8'd254; a_mant1 = 8'd64; a_mant2 = 8'd114; a_mant3 = 8'd239;
b_mant0 = 8'd77; b_mant1 = 8'd9; b_mant2 = 8'd233; b_mant3 = 8'd161;
a_exp0 = 10'd347; a_exp1 = 10'd223; a_exp2 = 10'd584; a_exp3 = 10'd412;
b_exp0 = 10'd65; b_exp1 = 10'd796; b_exp2 = 10'd760; b_exp3 = 10'd89;
a_sign0 = 4'd2; a_sign1 = 4'd7; a_sign2 = 4'd14; a_sign3 = 4'd2;
b_sign0 = 4'd6; b_sign1 = 4'd3; b_sign2 = 4'd13; b_sign3 = 4'd7;
@(posedge clk_i);
a_mant0 = 8'd245; a_mant1 = 8'd76; a_mant2 = 8'd79; a_mant3 = 8'd215;
b_mant0 = 8'd189; b_mant1 = 8'd160; b_mant2 = 8'd14; b_mant3 = 8'd35;
a_exp0 = 10'd630; a_exp1 = 10'd975; a_exp2 = 10'd563; a_exp3 = 10'd190;
b_exp0 = 10'd680; b_exp1 = 10'd779; b_exp2 = 10'd526; b_exp3 = 10'd403;
a_sign0 = 4'd6; a_sign1 = 4'd10; a_sign2 = 4'd14; a_sign3 = 4'd4;
b_sign0 = 4'd12; b_sign1 = 4'd12; b_sign2 = 4'd0; b_sign3 = 4'd1;
@(posedge clk_i);
a_mant0 = 8'd29; a_mant1 = 8'd248; a_mant2 = 8'd177; a_mant3 = 8'd222;
b_mant0 = 8'd105; b_mant1 = 8'd129; b_mant2 = 8'd49; b_mant3 = 8'd82;
a_exp0 = 10'd716; a_exp1 = 10'd750; a_exp2 = 10'd860; a_exp3 = 10'd256;
b_exp0 = 10'd173; b_exp1 = 10'd964; b_exp2 = 10'd31; b_exp3 = 10'd382;
a_sign0 = 4'd2; a_sign1 = 4'd8; a_sign2 = 4'd2; a_sign3 = 4'd16;
b_sign0 = 4'd2; b_sign1 = 4'd8; b_sign2 = 4'd5; b_sign3 = 4'd3;
@(posedge clk_i);
shared_exps0 = 8'd125;
shared_exps1 = 8'd108;
a_mant0 = 8'd57; a_mant1 = 8'd230; a_mant2 = 8'd206; a_mant3 = 8'd203;
b_mant0 = 8'd114; b_mant1 = 8'd141; b_mant2 = 8'd31; b_mant3 = 8'd33;
a_exp0 = 10'd858; a_exp1 = 10'd937; a_exp2 = 10'd570; a_exp3 = 10'd71;
b_exp0 = 10'd119; b_exp1 = 10'd889; b_exp2 = 10'd544; b_exp3 = 10'd118;
a_sign0 = 4'd7; a_sign1 = 4'd6; a_sign2 = 4'd2; a_sign3 = 4'd5;
b_sign0 = 4'd2; b_sign1 = 4'd13; b_sign2 = 4'd14; b_sign3 = 4'd1;
@(posedge clk_i);
a_mant0 = 8'd172; a_mant1 = 8'd61; a_mant2 = 8'd22; a_mant3 = 8'd96;
b_mant0 = 8'd40; b_mant1 = 8'd173; b_mant2 = 8'd240; b_mant3 = 8'd224;
a_exp0 = 10'd796; a_exp1 = 10'd530; a_exp2 = 10'd58; a_exp3 = 10'd626;
b_exp0 = 10'd172; b_exp1 = 10'd112; b_exp2 = 10'd309; b_exp3 = 10'd300;
a_sign0 = 4'd12; a_sign1 = 4'd10; a_sign2 = 4'd7; a_sign3 = 4'd8;
b_sign0 = 4'd6; b_sign1 = 4'd11; b_sign2 = 4'd6; b_sign3 = 4'd12;
@(posedge clk_i);
a_mant0 = 8'd28; a_mant1 = 8'd227; a_mant2 = 8'd236; a_mant3 = 8'd111;
b_mant0 = 8'd0; b_mant1 = 8'd125; b_mant2 = 8'd111; b_mant3 = 8'd242;
a_exp0 = 10'd184; a_exp1 = 10'd779; a_exp2 = 10'd449; a_exp3 = 10'd860;
b_exp0 = 10'd933; b_exp1 = 10'd318; b_exp2 = 10'd292; b_exp3 = 10'd284;
a_sign0 = 4'd6; a_sign1 = 4'd8; a_sign2 = 4'd1; a_sign3 = 4'd1;
b_sign0 = 4'd10; b_sign1 = 4'd9; b_sign2 = 4'd7; b_sign3 = 4'd14;
@(posedge clk_i);
a_mant0 = 8'd15; a_mant1 = 8'd197; a_mant2 = 8'd84; a_mant3 = 8'd117;
b_mant0 = 8'd51; b_mant1 = 8'd67; b_mant2 = 8'd26; b_mant3 = 8'd173;
a_exp0 = 10'd378; a_exp1 = 10'd527; a_exp2 = 10'd195; a_exp3 = 10'd230;
b_exp0 = 10'd343; b_exp1 = 10'd845; b_exp2 = 10'd204; b_exp3 = 10'd972;
a_sign0 = 4'd4; a_sign1 = 4'd15; a_sign2 = 4'd12; a_sign3 = 4'd0;
b_sign0 = 4'd16; b_sign1 = 4'd7; b_sign2 = 4'd3; b_sign3 = 4'd1;
@(posedge clk_i);
a_mant0 = 8'd109; a_mant1 = 8'd57; a_mant2 = 8'd154; a_mant3 = 8'd96;
b_mant0 = 8'd217; b_mant1 = 8'd132; b_mant2 = 8'd85; b_mant3 = 8'd141;
a_exp0 = 10'd257; a_exp1 = 10'd427; a_exp2 = 10'd460; a_exp3 = 10'd450;
b_exp0 = 10'd98; b_exp1 = 10'd408; b_exp2 = 10'd901; b_exp3 = 10'd515;
a_sign0 = 4'd6; a_sign1 = 4'd1; a_sign2 = 4'd5; a_sign3 = 4'd11;
b_sign0 = 4'd1; b_sign1 = 4'd4; b_sign2 = 4'd0; b_sign3 = 4'd5;
@(posedge clk_i);
a_mant0 = 8'd100; a_mant1 = 8'd195; a_mant2 = 8'd53; a_mant3 = 8'd9;
b_mant0 = 8'd135; b_mant1 = 8'd6; b_mant2 = 8'd165; b_mant3 = 8'd114;
a_exp0 = 10'd112; a_exp1 = 10'd653; a_exp2 = 10'd123; a_exp3 = 10'd270;
b_exp0 = 10'd324; b_exp1 = 10'd944; b_exp2 = 10'd688; b_exp3 = 10'd518;
a_sign0 = 4'd5; a_sign1 = 4'd4; a_sign2 = 4'd9; a_sign3 = 4'd12;
b_sign0 = 4'd1; b_sign1 = 4'd1; b_sign2 = 4'd14; b_sign3 = 4'd10;
@(posedge clk_i);
a_mant0 = 8'd51; a_mant1 = 8'd165; a_mant2 = 8'd209; a_mant3 = 8'd65;
b_mant0 = 8'd131; b_mant1 = 8'd208; b_mant2 = 8'd47; b_mant3 = 8'd151;
a_exp0 = 10'd822; a_exp1 = 10'd807; a_exp2 = 10'd158; a_exp3 = 10'd291;
b_exp0 = 10'd653; b_exp1 = 10'd118; b_exp2 = 10'd982; b_exp3 = 10'd887;
a_sign0 = 4'd13; a_sign1 = 4'd6; a_sign2 = 4'd0; a_sign3 = 4'd10;
b_sign0 = 4'd13; b_sign1 = 4'd7; b_sign2 = 4'd12; b_sign3 = 4'd16;
@(posedge clk_i);
a_mant0 = 8'd166; a_mant1 = 8'd194; a_mant2 = 8'd104; a_mant3 = 8'd190;
b_mant0 = 8'd190; b_mant1 = 8'd73; b_mant2 = 8'd159; b_mant3 = 8'd37;
a_exp0 = 10'd386; a_exp1 = 10'd320; a_exp2 = 10'd174; a_exp3 = 10'd420;
b_exp0 = 10'd806; b_exp1 = 10'd278; b_exp2 = 10'd467; b_exp3 = 10'd788;
a_sign0 = 4'd10; a_sign1 = 4'd6; a_sign2 = 4'd4; a_sign3 = 4'd15;
b_sign0 = 4'd11; b_sign1 = 4'd13; b_sign2 = 4'd5; b_sign3 = 4'd13;
@(posedge clk_i);
shared_exps0 = 8'd120;
shared_exps1 = 8'd137;
a_mant0 = 8'd155; a_mant1 = 8'd239; a_mant2 = 8'd193; a_mant3 = 8'd213;
b_mant0 = 8'd141; b_mant1 = 8'd53; b_mant2 = 8'd93; b_mant3 = 8'd12;
a_exp0 = 10'd760; a_exp1 = 10'd714; a_exp2 = 10'd123; a_exp3 = 10'd682;
b_exp0 = 10'd89; b_exp1 = 10'd660; b_exp2 = 10'd349; b_exp3 = 10'd564;
a_sign0 = 4'd16; a_sign1 = 4'd0; a_sign2 = 4'd2; a_sign3 = 4'd11;
b_sign0 = 4'd4; b_sign1 = 4'd11; b_sign2 = 4'd4; b_sign3 = 4'd8;
@(posedge clk_i);
a_mant0 = 8'd239; a_mant1 = 8'd39; a_mant2 = 8'd88; a_mant3 = 8'd196;
b_mant0 = 8'd6; b_mant1 = 8'd15; b_mant2 = 8'd161; b_mant3 = 8'd220;
a_exp0 = 10'd613; a_exp1 = 10'd479; a_exp2 = 10'd67; a_exp3 = 10'd856;
b_exp0 = 10'd358; b_exp1 = 10'd635; b_exp2 = 10'd302; b_exp3 = 10'd544;
a_sign0 = 4'd10; a_sign1 = 4'd11; a_sign2 = 4'd14; a_sign3 = 4'd9;
b_sign0 = 4'd16; b_sign1 = 4'd9; b_sign2 = 4'd10; b_sign3 = 4'd14;
@(posedge clk_i);
a_mant0 = 8'd66; a_mant1 = 8'd52; a_mant2 = 8'd241; a_mant3 = 8'd52;
b_mant0 = 8'd118; b_mant1 = 8'd135; b_mant2 = 8'd119; b_mant3 = 8'd188;
a_exp0 = 10'd612; a_exp1 = 10'd985; a_exp2 = 10'd619; a_exp3 = 10'd233;
b_exp0 = 10'd767; b_exp1 = 10'd338; b_exp2 = 10'd312; b_exp3 = 10'd941;
a_sign0 = 4'd10; a_sign1 = 4'd14; a_sign2 = 4'd2; a_sign3 = 4'd1;
b_sign0 = 4'd4; b_sign1 = 4'd15; b_sign2 = 4'd10; b_sign3 = 4'd11;
@(posedge clk_i);
a_mant0 = 8'd197; a_mant1 = 8'd5; a_mant2 = 8'd159; a_mant3 = 8'd37;
b_mant0 = 8'd20; b_mant1 = 8'd106; b_mant2 = 8'd66; b_mant3 = 8'd22;
a_exp0 = 10'd311; a_exp1 = 10'd671; a_exp2 = 10'd956; a_exp3 = 10'd815;
b_exp0 = 10'd790; b_exp1 = 10'd9; b_exp2 = 10'd342; b_exp3 = 10'd442;
a_sign0 = 4'd3; a_sign1 = 4'd5; a_sign2 = 4'd0; a_sign3 = 4'd16;
b_sign0 = 4'd6; b_sign1 = 4'd1; b_sign2 = 4'd9; b_sign3 = 4'd4;
@(posedge clk_i);
a_mant0 = 8'd134; a_mant1 = 8'd132; a_mant2 = 8'd117; a_mant3 = 8'd234;
b_mant0 = 8'd44; b_mant1 = 8'd118; b_mant2 = 8'd129; b_mant3 = 8'd229;
a_exp0 = 10'd962; a_exp1 = 10'd102; a_exp2 = 10'd385; a_exp3 = 10'd342;
b_exp0 = 10'd236; b_exp1 = 10'd953; b_exp2 = 10'd772; b_exp3 = 10'd855;
a_sign0 = 4'd12; a_sign1 = 4'd7; a_sign2 = 4'd8; a_sign3 = 4'd10;
b_sign0 = 4'd13; b_sign1 = 4'd11; b_sign2 = 4'd12; b_sign3 = 4'd11;
@(posedge clk_i);
a_mant0 = 8'd3; a_mant1 = 8'd229; a_mant2 = 8'd157; a_mant3 = 8'd1;
b_mant0 = 8'd169; b_mant1 = 8'd54; b_mant2 = 8'd248; b_mant3 = 8'd34;
a_exp0 = 10'd108; a_exp1 = 10'd549; a_exp2 = 10'd601; a_exp3 = 10'd174;
b_exp0 = 10'd990; b_exp1 = 10'd672; b_exp2 = 10'd673; b_exp3 = 10'd683;
a_sign0 = 4'd16; a_sign1 = 4'd8; a_sign2 = 4'd11; a_sign3 = 4'd7;
b_sign0 = 4'd12; b_sign1 = 4'd11; b_sign2 = 4'd13; b_sign3 = 4'd5;
@(posedge clk_i);
a_mant0 = 8'd139; a_mant1 = 8'd85; a_mant2 = 8'd236; a_mant3 = 8'd196;
b_mant0 = 8'd5; b_mant1 = 8'd254; b_mant2 = 8'd47; b_mant3 = 8'd71;
a_exp0 = 10'd989; a_exp1 = 10'd971; a_exp2 = 10'd570; a_exp3 = 10'd753;
b_exp0 = 10'd872; b_exp1 = 10'd868; b_exp2 = 10'd671; b_exp3 = 10'd165;
a_sign0 = 4'd14; a_sign1 = 4'd7; a_sign2 = 4'd12; a_sign3 = 4'd2;
b_sign0 = 4'd0; b_sign1 = 4'd3; b_sign2 = 4'd16; b_sign3 = 4'd5;
@(posedge clk_i);
a_mant0 = 8'd3; a_mant1 = 8'd203; a_mant2 = 8'd139; a_mant3 = 8'd79;
b_mant0 = 8'd135; b_mant1 = 8'd136; b_mant2 = 8'd115; b_mant3 = 8'd9;
a_exp0 = 10'd120; a_exp1 = 10'd433; a_exp2 = 10'd546; a_exp3 = 10'd421;
b_exp0 = 10'd3; b_exp1 = 10'd434; b_exp2 = 10'd543; b_exp3 = 10'd274;
a_sign0 = 4'd11; a_sign1 = 4'd11; a_sign2 = 4'd10; a_sign3 = 4'd16;
b_sign0 = 4'd15; b_sign1 = 4'd11; b_sign2 = 4'd14; b_sign3 = 4'd11;
@(posedge clk_i);
shared_exps0 = 8'd131;
shared_exps1 = 8'd132;
rstn = 0;
@(posedge clk_i);
rstn = 1;
a_mant0 = 8'd254; a_mant1 = 8'd162; a_mant2 = 8'd90; a_mant3 = 8'd154;
b_mant0 = 8'd132; b_mant1 = 8'd249; b_mant2 = 8'd103; b_mant3 = 8'd57;
a_exp0 = 10'd243; a_exp1 = 10'd850; a_exp2 = 10'd839; a_exp3 = 10'd351;
b_exp0 = 10'd434; b_exp1 = 10'd339; b_exp2 = 10'd354; b_exp3 = 10'd52;
a_sign0 = 4'd3; a_sign1 = 4'd1; a_sign2 = 4'd6; a_sign3 = 4'd11;
b_sign0 = 4'd12; b_sign1 = 4'd6; b_sign2 = 4'd1; b_sign3 = 4'd14;
@(posedge clk_i);
a_mant0 = 8'd193; a_mant1 = 8'd156; a_mant2 = 8'd179; a_mant3 = 8'd199;
b_mant0 = 8'd238; b_mant1 = 8'd172; b_mant2 = 8'd49; b_mant3 = 8'd91;
a_exp0 = 10'd853; a_exp1 = 10'd47; a_exp2 = 10'd685; a_exp3 = 10'd358;
b_exp0 = 10'd455; b_exp1 = 10'd488; b_exp2 = 10'd765; b_exp3 = 10'd766;
a_sign0 = 4'd16; a_sign1 = 4'd8; a_sign2 = 4'd8; a_sign3 = 4'd6;
b_sign0 = 4'd9; b_sign1 = 4'd13; b_sign2 = 4'd3; b_sign3 = 4'd12;
@(posedge clk_i);
a_mant0 = 8'd33; a_mant1 = 8'd100; a_mant2 = 8'd61; a_mant3 = 8'd116;
b_mant0 = 8'd181; b_mant1 = 8'd202; b_mant2 = 8'd148; b_mant3 = 8'd90;
a_exp0 = 10'd379; a_exp1 = 10'd900; a_exp2 = 10'd90; a_exp3 = 10'd793;
b_exp0 = 10'd3; b_exp1 = 10'd951; b_exp2 = 10'd92; b_exp3 = 10'd349;
a_sign0 = 4'd13; a_sign1 = 4'd2; a_sign2 = 4'd3; a_sign3 = 4'd10;
b_sign0 = 4'd10; b_sign1 = 4'd8; b_sign2 = 4'd13; b_sign3 = 4'd7;
@(posedge clk_i);
a_mant0 = 8'd176; a_mant1 = 8'd50; a_mant2 = 8'd189; a_mant3 = 8'd14;
b_mant0 = 8'd78; b_mant1 = 8'd255; b_mant2 = 8'd208; b_mant3 = 8'd96;
a_exp0 = 10'd525; a_exp1 = 10'd159; a_exp2 = 10'd314; a_exp3 = 10'd634;
b_exp0 = 10'd333; b_exp1 = 10'd433; b_exp2 = 10'd588; b_exp3 = 10'd735;
a_sign0 = 4'd2; a_sign1 = 4'd0; a_sign2 = 4'd11; a_sign3 = 4'd10;
b_sign0 = 4'd5; b_sign1 = 4'd3; b_sign2 = 4'd1; b_sign3 = 4'd10;
@(posedge clk_i);
a_mant0 = 8'd72; a_mant1 = 8'd220; a_mant2 = 8'd9; a_mant3 = 8'd63;
b_mant0 = 8'd111; b_mant1 = 8'd28; b_mant2 = 8'd192; b_mant3 = 8'd142;
a_exp0 = 10'd135; a_exp1 = 10'd901; a_exp2 = 10'd255; a_exp3 = 10'd870;
b_exp0 = 10'd748; b_exp1 = 10'd398; b_exp2 = 10'd52; b_exp3 = 10'd196;
a_sign0 = 4'd5; a_sign1 = 4'd16; a_sign2 = 4'd0; a_sign3 = 4'd11;
b_sign0 = 4'd14; b_sign1 = 4'd8; b_sign2 = 4'd9; b_sign3 = 4'd10;
@(posedge clk_i);
a_mant0 = 8'd226; a_mant1 = 8'd235; a_mant2 = 8'd56; a_mant3 = 8'd89;
b_mant0 = 8'd192; b_mant1 = 8'd197; b_mant2 = 8'd154; b_mant3 = 8'd141;
a_exp0 = 10'd625; a_exp1 = 10'd975; a_exp2 = 10'd936; a_exp3 = 10'd709;
b_exp0 = 10'd5; b_exp1 = 10'd573; b_exp2 = 10'd812; b_exp3 = 10'd770;
a_sign0 = 4'd14; a_sign1 = 4'd1; a_sign2 = 4'd11; a_sign3 = 4'd12;
b_sign0 = 4'd12; b_sign1 = 4'd5; b_sign2 = 4'd0; b_sign3 = 4'd0;
@(posedge clk_i);
a_mant0 = 8'd216; a_mant1 = 8'd94; a_mant2 = 8'd76; a_mant3 = 8'd125;
b_mant0 = 8'd249; b_mant1 = 8'd105; b_mant2 = 8'd120; b_mant3 = 8'd27;
a_exp0 = 10'd331; a_exp1 = 10'd271; a_exp2 = 10'd619; a_exp3 = 10'd102;
b_exp0 = 10'd151; b_exp1 = 10'd320; b_exp2 = 10'd523; b_exp3 = 10'd436;
a_sign0 = 4'd4; a_sign1 = 4'd0; a_sign2 = 4'd3; a_sign3 = 4'd11;
b_sign0 = 4'd7; b_sign1 = 4'd13; b_sign2 = 4'd5; b_sign3 = 4'd16;
@(posedge clk_i);
shared_exps0 = 8'd143;
shared_exps1 = 8'd121;
a_mant0 = 8'd95; a_mant1 = 8'd226; a_mant2 = 8'd116; a_mant3 = 8'd46;
b_mant0 = 8'd156; b_mant1 = 8'd50; b_mant2 = 8'd87; b_mant3 = 8'd136;
a_exp0 = 10'd407; a_exp1 = 10'd883; a_exp2 = 10'd905; a_exp3 = 10'd236;
b_exp0 = 10'd425; b_exp1 = 10'd844; b_exp2 = 10'd373; b_exp3 = 10'd515;
a_sign0 = 4'd0; a_sign1 = 4'd8; a_sign2 = 4'd4; a_sign3 = 4'd1;
b_sign0 = 4'd4; b_sign1 = 4'd3; b_sign2 = 4'd13; b_sign3 = 4'd2;
@(posedge clk_i);
a_mant0 = 8'd56; a_mant1 = 8'd15; a_mant2 = 8'd96; a_mant3 = 8'd53;
b_mant0 = 8'd250; b_mant1 = 8'd217; b_mant2 = 8'd64; b_mant3 = 8'd187;
a_exp0 = 10'd92; a_exp1 = 10'd556; a_exp2 = 10'd517; a_exp3 = 10'd724;
b_exp0 = 10'd294; b_exp1 = 10'd856; b_exp2 = 10'd559; b_exp3 = 10'd196;
a_sign0 = 4'd7; a_sign1 = 4'd4; a_sign2 = 4'd9; a_sign3 = 4'd11;
b_sign0 = 4'd7; b_sign1 = 4'd10; b_sign2 = 4'd16; b_sign3 = 4'd5;
@(posedge clk_i);
a_mant0 = 8'd84; a_mant1 = 8'd23; a_mant2 = 8'd137; a_mant3 = 8'd190;
b_mant0 = 8'd80; b_mant1 = 8'd67; b_mant2 = 8'd245; b_mant3 = 8'd156;
a_exp0 = 10'd706; a_exp1 = 10'd699; a_exp2 = 10'd28; a_exp3 = 10'd1005;
b_exp0 = 10'd63; b_exp1 = 10'd468; b_exp2 = 10'd505; b_exp3 = 10'd799;
a_sign0 = 4'd11; a_sign1 = 4'd1; a_sign2 = 4'd9; a_sign3 = 4'd3;
b_sign0 = 4'd6; b_sign1 = 4'd4; b_sign2 = 4'd8; b_sign3 = 4'd1;
@(posedge clk_i);
a_mant0 = 8'd239; a_mant1 = 8'd175; a_mant2 = 8'd216; a_mant3 = 8'd20;
b_mant0 = 8'd108; b_mant1 = 8'd237; b_mant2 = 8'd176; b_mant3 = 8'd114;
a_exp0 = 10'd887; a_exp1 = 10'd154; a_exp2 = 10'd444; a_exp3 = 10'd555;
b_exp0 = 10'd728; b_exp1 = 10'd265; b_exp2 = 10'd356; b_exp3 = 10'd538;
a_sign0 = 4'd11; a_sign1 = 4'd7; a_sign2 = 4'd7; a_sign3 = 4'd8;
b_sign0 = 4'd2; b_sign1 = 4'd6; b_sign2 = 4'd12; b_sign3 = 4'd10;
@(posedge clk_i);
a_mant0 = 8'd27; a_mant1 = 8'd234; a_mant2 = 8'd66; a_mant3 = 8'd40;
b_mant0 = 8'd34; b_mant1 = 8'd93; b_mant2 = 8'd167; b_mant3 = 8'd32;
a_exp0 = 10'd575; a_exp1 = 10'd213; a_exp2 = 10'd142; a_exp3 = 10'd791;
b_exp0 = 10'd616; b_exp1 = 10'd369; b_exp2 = 10'd400; b_exp3 = 10'd657;
a_sign0 = 4'd12; a_sign1 = 4'd6; a_sign2 = 4'd9; a_sign3 = 4'd5;
b_sign0 = 4'd13; b_sign1 = 4'd2; b_sign2 = 4'd10; b_sign3 = 4'd13;
@(posedge clk_i);
a_mant0 = 8'd223; a_mant1 = 8'd88; a_mant2 = 8'd87; a_mant3 = 8'd104;
b_mant0 = 8'd9; b_mant1 = 8'd76; b_mant2 = 8'd138; b_mant3 = 8'd180;
a_exp0 = 10'd280; a_exp1 = 10'd863; a_exp2 = 10'd527; a_exp3 = 10'd279;
b_exp0 = 10'd64; b_exp1 = 10'd668; b_exp2 = 10'd79; b_exp3 = 10'd411;
a_sign0 = 4'd11; a_sign1 = 4'd9; a_sign2 = 4'd12; a_sign3 = 4'd0;
b_sign0 = 4'd11; b_sign1 = 4'd13; b_sign2 = 4'd9; b_sign3 = 4'd4;
@(posedge clk_i);
a_mant0 = 8'd32; a_mant1 = 8'd208; a_mant2 = 8'd169; a_mant3 = 8'd125;
b_mant0 = 8'd233; b_mant1 = 8'd155; b_mant2 = 8'd176; b_mant3 = 8'd94;
a_exp0 = 10'd130; a_exp1 = 10'd978; a_exp2 = 10'd15; a_exp3 = 10'd789;
b_exp0 = 10'd469; b_exp1 = 10'd863; b_exp2 = 10'd205; b_exp3 = 10'd821;
a_sign0 = 4'd5; a_sign1 = 4'd1; a_sign2 = 4'd10; a_sign3 = 4'd13;
b_sign0 = 4'd16; b_sign1 = 4'd3; b_sign2 = 4'd7; b_sign3 = 4'd7;
@(posedge clk_i);
a_mant0 = 8'd139; a_mant1 = 8'd131; a_mant2 = 8'd90; a_mant3 = 8'd203;
b_mant0 = 8'd100; b_mant1 = 8'd101; b_mant2 = 8'd61; b_mant3 = 8'd57;
a_exp0 = 10'd369; a_exp1 = 10'd751; a_exp2 = 10'd531; a_exp3 = 10'd781;
b_exp0 = 10'd200; b_exp1 = 10'd203; b_exp2 = 10'd1011; b_exp3 = 10'd182;
a_sign0 = 4'd5; a_sign1 = 4'd14; a_sign2 = 4'd10; a_sign3 = 4'd14;
b_sign0 = 4'd8; b_sign1 = 4'd9; b_sign2 = 4'd7; b_sign3 = 4'd5;
@(posedge clk_i);
shared_exps0 = 8'd118;
shared_exps1 = 8'd120;
a_mant0 = 8'd61; a_mant1 = 8'd38; a_mant2 = 8'd192; a_mant3 = 8'd12;
b_mant0 = 8'd83; b_mant1 = 8'd77; b_mant2 = 8'd104; b_mant3 = 8'd61;
a_exp0 = 10'd939; a_exp1 = 10'd134; a_exp2 = 10'd774; a_exp3 = 10'd786;
b_exp0 = 10'd100; b_exp1 = 10'd529; b_exp2 = 10'd679; b_exp3 = 10'd351;
a_sign0 = 4'd7; a_sign1 = 4'd13; a_sign2 = 4'd13; a_sign3 = 4'd12;
b_sign0 = 4'd1; b_sign1 = 4'd15; b_sign2 = 4'd9; b_sign3 = 4'd15;
@(posedge clk_i);
a_mant0 = 8'd83; a_mant1 = 8'd181; a_mant2 = 8'd131; a_mant3 = 8'd183;
b_mant0 = 8'd31; b_mant1 = 8'd11; b_mant2 = 8'd83; b_mant3 = 8'd217;
a_exp0 = 10'd624; a_exp1 = 10'd491; a_exp2 = 10'd148; a_exp3 = 10'd297;
b_exp0 = 10'd969; b_exp1 = 10'd420; b_exp2 = 10'd129; b_exp3 = 10'd972;
a_sign0 = 4'd9; a_sign1 = 4'd13; a_sign2 = 4'd5; a_sign3 = 4'd5;
b_sign0 = 4'd15; b_sign1 = 4'd10; b_sign2 = 4'd15; b_sign3 = 4'd5;
@(posedge clk_i);
a_mant0 = 8'd123; a_mant1 = 8'd121; a_mant2 = 8'd199; a_mant3 = 8'd42;
b_mant0 = 8'd75; b_mant1 = 8'd39; b_mant2 = 8'd100; b_mant3 = 8'd53;
a_exp0 = 10'd793; a_exp1 = 10'd230; a_exp2 = 10'd481; a_exp3 = 10'd768;
b_exp0 = 10'd891; b_exp1 = 10'd697; b_exp2 = 10'd665; b_exp3 = 10'd951;
a_sign0 = 4'd2; a_sign1 = 4'd4; a_sign2 = 4'd6; a_sign3 = 4'd16;
b_sign0 = 4'd2; b_sign1 = 4'd2; b_sign2 = 4'd7; b_sign3 = 4'd11;
@(posedge clk_i);
a_mant0 = 8'd0; a_mant1 = 8'd86; a_mant2 = 8'd229; a_mant3 = 8'd68;
b_mant0 = 8'd89; b_mant1 = 8'd182; b_mant2 = 8'd104; b_mant3 = 8'd7;
a_exp0 = 10'd542; a_exp1 = 10'd179; a_exp2 = 10'd435; a_exp3 = 10'd499;
b_exp0 = 10'd162; b_exp1 = 10'd841; b_exp2 = 10'd180; b_exp3 = 10'd683;
a_sign0 = 4'd2; a_sign1 = 4'd9; a_sign2 = 4'd2; a_sign3 = 4'd6;
b_sign0 = 4'd0; b_sign1 = 4'd12; b_sign2 = 4'd1; b_sign3 = 4'd6;
@(posedge clk_i);
a_mant0 = 8'd60; a_mant1 = 8'd12; a_mant2 = 8'd238; a_mant3 = 8'd166;
b_mant0 = 8'd183; b_mant1 = 8'd135; b_mant2 = 8'd219; b_mant3 = 8'd219;
a_exp0 = 10'd853; a_exp1 = 10'd937; a_exp2 = 10'd582; a_exp3 = 10'd26;
b_exp0 = 10'd293; b_exp1 = 10'd953; b_exp2 = 10'd526; b_exp3 = 10'd587;
a_sign0 = 4'd9; a_sign1 = 4'd1; a_sign2 = 4'd1; a_sign3 = 4'd12;
b_sign0 = 4'd14; b_sign1 = 4'd2; b_sign2 = 4'd14; b_sign3 = 4'd12;
@(posedge clk_i);
a_mant0 = 8'd156; a_mant1 = 8'd220; a_mant2 = 8'd17; a_mant3 = 8'd136;
b_mant0 = 8'd228; b_mant1 = 8'd226; b_mant2 = 8'd63; b_mant3 = 8'd82;
a_exp0 = 10'd79; a_exp1 = 10'd57; a_exp2 = 10'd14; a_exp3 = 10'd41;
b_exp0 = 10'd367; b_exp1 = 10'd85; b_exp2 = 10'd799; b_exp3 = 10'd384;
a_sign0 = 4'd13; a_sign1 = 4'd8; a_sign2 = 4'd10; a_sign3 = 4'd12;
b_sign0 = 4'd14; b_sign1 = 4'd5; b_sign2 = 4'd16; b_sign3 = 4'd9;
@(posedge clk_i);
a_mant0 = 8'd4; a_mant1 = 8'd172; a_mant2 = 8'd197; a_mant3 = 8'd138;
b_mant0 = 8'd51; b_mant1 = 8'd137; b_mant2 = 8'd81; b_mant3 = 8'd231;
a_exp0 = 10'd462; a_exp1 = 10'd471; a_exp2 = 10'd846; a_exp3 = 10'd277;
b_exp0 = 10'd890; b_exp1 = 10'd750; b_exp2 = 10'd165; b_exp3 = 10'd86;
a_sign0 = 4'd15; a_sign1 = 4'd10; a_sign2 = 4'd2; a_sign3 = 4'd16;
b_sign0 = 4'd3; b_sign1 = 4'd5; b_sign2 = 4'd9; b_sign3 = 4'd12;
@(posedge clk_i);
a_mant0 = 8'd183; a_mant1 = 8'd51; a_mant2 = 8'd199; a_mant3 = 8'd14;
b_mant0 = 8'd79; b_mant1 = 8'd58; b_mant2 = 8'd3; b_mant3 = 8'd63;
a_exp0 = 10'd746; a_exp1 = 10'd37; a_exp2 = 10'd712; a_exp3 = 10'd1021;
b_exp0 = 10'd407; b_exp1 = 10'd775; b_exp2 = 10'd940; b_exp3 = 10'd497;
a_sign0 = 4'd10; a_sign1 = 4'd7; a_sign2 = 4'd3; a_sign3 = 4'd4;
b_sign0 = 4'd0; b_sign1 = 4'd5; b_sign2 = 4'd11; b_sign3 = 4'd5;
@(posedge clk_i);
shared_exps0 = 8'd114;
shared_exps1 = 8'd126;
a_mant0 = 8'd50; a_mant1 = 8'd87; a_mant2 = 8'd64; a_mant3 = 8'd33;
b_mant0 = 8'd66; b_mant1 = 8'd36; b_mant2 = 8'd144; b_mant3 = 8'd21;
a_exp0 = 10'd133; a_exp1 = 10'd35; a_exp2 = 10'd1023; a_exp3 = 10'd43;
b_exp0 = 10'd450; b_exp1 = 10'd425; b_exp2 = 10'd909; b_exp3 = 10'd817;
a_sign0 = 4'd5; a_sign1 = 4'd0; a_sign2 = 4'd3; a_sign3 = 4'd4;
b_sign0 = 4'd7; b_sign1 = 4'd14; b_sign2 = 4'd2; b_sign3 = 4'd2;
@(posedge clk_i);
a_mant0 = 8'd186; a_mant1 = 8'd140; a_mant2 = 8'd194; a_mant3 = 8'd66;
b_mant0 = 8'd200; b_mant1 = 8'd100; b_mant2 = 8'd38; b_mant3 = 8'd59;
a_exp0 = 10'd874; a_exp1 = 10'd913; a_exp2 = 10'd1; a_exp3 = 10'd340;
b_exp0 = 10'd639; b_exp1 = 10'd383; b_exp2 = 10'd234; b_exp3 = 10'd338;
a_sign0 = 4'd5; a_sign1 = 4'd14; a_sign2 = 4'd2; a_sign3 = 4'd3;
b_sign0 = 4'd15; b_sign1 = 4'd14; b_sign2 = 4'd13; b_sign3 = 4'd6;
@(posedge clk_i);
a_mant0 = 8'd93; a_mant1 = 8'd180; a_mant2 = 8'd240; a_mant3 = 8'd142;
b_mant0 = 8'd78; b_mant1 = 8'd183; b_mant2 = 8'd128; b_mant3 = 8'd244;
a_exp0 = 10'd949; a_exp1 = 10'd250; a_exp2 = 10'd629; a_exp3 = 10'd592;
b_exp0 = 10'd967; b_exp1 = 10'd838; b_exp2 = 10'd523; b_exp3 = 10'd712;
a_sign0 = 4'd13; a_sign1 = 4'd11; a_sign2 = 4'd8; a_sign3 = 4'd14;
b_sign0 = 4'd13; b_sign1 = 4'd16; b_sign2 = 4'd0; b_sign3 = 4'd1;
@(posedge clk_i);
a_mant0 = 8'd120; a_mant1 = 8'd210; a_mant2 = 8'd29; a_mant3 = 8'd155;
b_mant0 = 8'd209; b_mant1 = 8'd162; b_mant2 = 8'd11; b_mant3 = 8'd194;
a_exp0 = 10'd857; a_exp1 = 10'd624; a_exp2 = 10'd675; a_exp3 = 10'd445;
b_exp0 = 10'd190; b_exp1 = 10'd659; b_exp2 = 10'd126; b_exp3 = 10'd788;
a_sign0 = 4'd11; a_sign1 = 4'd12; a_sign2 = 4'd5; a_sign3 = 4'd3;
b_sign0 = 4'd15; b_sign1 = 4'd8; b_sign2 = 4'd12; b_sign3 = 4'd1;
@(posedge clk_i);
a_mant0 = 8'd229; a_mant1 = 8'd89; a_mant2 = 8'd53; a_mant3 = 8'd96;
b_mant0 = 8'd121; b_mant1 = 8'd96; b_mant2 = 8'd16; b_mant3 = 8'd3;
a_exp0 = 10'd139; a_exp1 = 10'd675; a_exp2 = 10'd7; a_exp3 = 10'd321;
b_exp0 = 10'd365; b_exp1 = 10'd118; b_exp2 = 10'd267; b_exp3 = 10'd470;
a_sign0 = 4'd13; a_sign1 = 4'd4; a_sign2 = 4'd2; a_sign3 = 4'd3;
b_sign0 = 4'd4; b_sign1 = 4'd2; b_sign2 = 4'd5; b_sign3 = 4'd6;
@(posedge clk_i);
a_mant0 = 8'd203; a_mant1 = 8'd228; a_mant2 = 8'd192; a_mant3 = 8'd124;
b_mant0 = 8'd244; b_mant1 = 8'd176; b_mant2 = 8'd148; b_mant3 = 8'd29;
a_exp0 = 10'd846; a_exp1 = 10'd212; a_exp2 = 10'd814; a_exp3 = 10'd844;
b_exp0 = 10'd276; b_exp1 = 10'd171; b_exp2 = 10'd836; b_exp3 = 10'd430;
a_sign0 = 4'd4; a_sign1 = 4'd12; a_sign2 = 4'd7; a_sign3 = 4'd4;
b_sign0 = 4'd12; b_sign1 = 4'd15; b_sign2 = 4'd6; b_sign3 = 4'd15;
@(posedge clk_i);
a_mant0 = 8'd208; a_mant1 = 8'd183; a_mant2 = 8'd176; a_mant3 = 8'd185;
b_mant0 = 8'd42; b_mant1 = 8'd8; b_mant2 = 8'd35; b_mant3 = 8'd217;
a_exp0 = 10'd128; a_exp1 = 10'd622; a_exp2 = 10'd55; a_exp3 = 10'd427;
b_exp0 = 10'd559; b_exp1 = 10'd374; b_exp2 = 10'd707; b_exp3 = 10'd626;
a_sign0 = 4'd8; a_sign1 = 4'd15; a_sign2 = 4'd16; a_sign3 = 4'd12;
b_sign0 = 4'd3; b_sign1 = 4'd1; b_sign2 = 4'd4; b_sign3 = 4'd0;
@(posedge clk_i);
a_mant0 = 8'd184; a_mant1 = 8'd43; a_mant2 = 8'd58; a_mant3 = 8'd137;
b_mant0 = 8'd94; b_mant1 = 8'd241; b_mant2 = 8'd96; b_mant3 = 8'd88;
a_exp0 = 10'd766; a_exp1 = 10'd252; a_exp2 = 10'd663; a_exp3 = 10'd440;
b_exp0 = 10'd442; b_exp1 = 10'd346; b_exp2 = 10'd48; b_exp3 = 10'd138;
a_sign0 = 4'd0; a_sign1 = 4'd2; a_sign2 = 4'd10; a_sign3 = 4'd12;
b_sign0 = 4'd7; b_sign1 = 4'd2; b_sign2 = 4'd4; b_sign3 = 4'd6;
@(posedge clk_i);
shared_exps0 = 8'd100;
shared_exps1 = 8'd113;
rstn = 0;
@(posedge clk_i);
rstn = 1;
a_mant0 = 8'd50; a_mant1 = 8'd119; a_mant2 = 8'd198; a_mant3 = 8'd212;
b_mant0 = 8'd21; b_mant1 = 8'd227; b_mant2 = 8'd249; b_mant3 = 8'd60;
a_exp0 = 10'd865; a_exp1 = 10'd892; a_exp2 = 10'd457; a_exp3 = 10'd651;
b_exp0 = 10'd419; b_exp1 = 10'd561; b_exp2 = 10'd632; b_exp3 = 10'd266;
a_sign0 = 4'd16; a_sign1 = 4'd3; a_sign2 = 4'd3; a_sign3 = 4'd3;
b_sign0 = 4'd4; b_sign1 = 4'd11; b_sign2 = 4'd13; b_sign3 = 4'd8;
@(posedge clk_i);
a_mant0 = 8'd65; a_mant1 = 8'd77; a_mant2 = 8'd16; a_mant3 = 8'd16;
b_mant0 = 8'd120; b_mant1 = 8'd19; b_mant2 = 8'd12; b_mant3 = 8'd53;
a_exp0 = 10'd478; a_exp1 = 10'd973; a_exp2 = 10'd308; a_exp3 = 10'd648;
b_exp0 = 10'd899; b_exp1 = 10'd672; b_exp2 = 10'd21; b_exp3 = 10'd525;
a_sign0 = 4'd10; a_sign1 = 4'd8; a_sign2 = 4'd8; a_sign3 = 4'd13;
b_sign0 = 4'd1; b_sign1 = 4'd11; b_sign2 = 4'd6; b_sign3 = 4'd2;
@(posedge clk_i);
a_mant0 = 8'd13; a_mant1 = 8'd105; a_mant2 = 8'd10; a_mant3 = 8'd83;
b_mant0 = 8'd2; b_mant1 = 8'd28; b_mant2 = 8'd85; b_mant3 = 8'd24;
a_exp0 = 10'd264; a_exp1 = 10'd656; a_exp2 = 10'd919; a_exp3 = 10'd847;
b_exp0 = 10'd795; b_exp1 = 10'd687; b_exp2 = 10'd954; b_exp3 = 10'd557;
a_sign0 = 4'd16; a_sign1 = 4'd11; a_sign2 = 4'd1; a_sign3 = 4'd5;
b_sign0 = 4'd15; b_sign1 = 4'd4; b_sign2 = 4'd11; b_sign3 = 4'd8;
@(posedge clk_i);
a_mant0 = 8'd118; a_mant1 = 8'd148; a_mant2 = 8'd228; a_mant3 = 8'd72;
b_mant0 = 8'd134; b_mant1 = 8'd158; b_mant2 = 8'd90; b_mant3 = 8'd177;
a_exp0 = 10'd818; a_exp1 = 10'd629; a_exp2 = 10'd191; a_exp3 = 10'd84;
b_exp0 = 10'd752; b_exp1 = 10'd704; b_exp2 = 10'd772; b_exp3 = 10'd721;
a_sign0 = 4'd1; a_sign1 = 4'd11; a_sign2 = 4'd16; a_sign3 = 4'd14;
b_sign0 = 4'd10; b_sign1 = 4'd6; b_sign2 = 4'd4; b_sign3 = 4'd0;
@(posedge clk_i);
a_mant0 = 8'd73; a_mant1 = 8'd207; a_mant2 = 8'd224; a_mant3 = 8'd17;
b_mant0 = 8'd201; b_mant1 = 8'd161; b_mant2 = 8'd165; b_mant3 = 8'd134;
a_exp0 = 10'd196; a_exp1 = 10'd459; a_exp2 = 10'd609; a_exp3 = 10'd838;
b_exp0 = 10'd737; b_exp1 = 10'd106; b_exp2 = 10'd999; b_exp3 = 10'd97;
a_sign0 = 4'd9; a_sign1 = 4'd12; a_sign2 = 4'd13; a_sign3 = 4'd12;
b_sign0 = 4'd9; b_sign1 = 4'd1; b_sign2 = 4'd1; b_sign3 = 4'd2;
@(posedge clk_i);
a_mant0 = 8'd233; a_mant1 = 8'd249; a_mant2 = 8'd233; a_mant3 = 8'd158;
b_mant0 = 8'd200; b_mant1 = 8'd225; b_mant2 = 8'd230; b_mant3 = 8'd155;
a_exp0 = 10'd809; a_exp1 = 10'd237; a_exp2 = 10'd561; a_exp3 = 10'd477;
b_exp0 = 10'd394; b_exp1 = 10'd501; b_exp2 = 10'd134; b_exp3 = 10'd404;
a_sign0 = 4'd16; a_sign1 = 4'd3; a_sign2 = 4'd6; a_sign3 = 4'd4;
b_sign0 = 4'd8; b_sign1 = 4'd10; b_sign2 = 4'd4; b_sign3 = 4'd4;
@(posedge clk_i);
a_mant0 = 8'd10; a_mant1 = 8'd101; a_mant2 = 8'd31; a_mant3 = 8'd13;
b_mant0 = 8'd0; b_mant1 = 8'd198; b_mant2 = 8'd237; b_mant3 = 8'd122;
a_exp0 = 10'd863; a_exp1 = 10'd25; a_exp2 = 10'd852; a_exp3 = 10'd634;
b_exp0 = 10'd792; b_exp1 = 10'd653; b_exp2 = 10'd811; b_exp3 = 10'd903;
a_sign0 = 4'd5; a_sign1 = 4'd15; a_sign2 = 4'd16; a_sign3 = 4'd1;
b_sign0 = 4'd15; b_sign1 = 4'd6; b_sign2 = 4'd10; b_sign3 = 4'd3;
@(posedge clk_i);
shared_exps0 = 8'd136;
shared_exps1 = 8'd139;
a_mant0 = 8'd250; a_mant1 = 8'd239; a_mant2 = 8'd175; a_mant3 = 8'd136;
b_mant0 = 8'd34; b_mant1 = 8'd33; b_mant2 = 8'd87; b_mant3 = 8'd131;
a_exp0 = 10'd931; a_exp1 = 10'd907; a_exp2 = 10'd106; a_exp3 = 10'd118;
b_exp0 = 10'd413; b_exp1 = 10'd56; b_exp2 = 10'd113; b_exp3 = 10'd451;
a_sign0 = 4'd10; a_sign1 = 4'd14; a_sign2 = 4'd12; a_sign3 = 4'd10;
b_sign0 = 4'd13; b_sign1 = 4'd1; b_sign2 = 4'd7; b_sign3 = 4'd16;
@(posedge clk_i);
a_mant0 = 8'd198; a_mant1 = 8'd231; a_mant2 = 8'd175; a_mant3 = 8'd58;
b_mant0 = 8'd153; b_mant1 = 8'd183; b_mant2 = 8'd3; b_mant3 = 8'd70;
a_exp0 = 10'd99; a_exp1 = 10'd510; a_exp2 = 10'd61; a_exp3 = 10'd144;
b_exp0 = 10'd220; b_exp1 = 10'd14; b_exp2 = 10'd428; b_exp3 = 10'd279;
a_sign0 = 4'd9; a_sign1 = 4'd6; a_sign2 = 4'd10; a_sign3 = 4'd7;
b_sign0 = 4'd12; b_sign1 = 4'd15; b_sign2 = 4'd8; b_sign3 = 4'd7;
@(posedge clk_i);
a_mant0 = 8'd115; a_mant1 = 8'd191; a_mant2 = 8'd190; a_mant3 = 8'd2;
b_mant0 = 8'd107; b_mant1 = 8'd102; b_mant2 = 8'd42; b_mant3 = 8'd63;
a_exp0 = 10'd476; a_exp1 = 10'd181; a_exp2 = 10'd347; a_exp3 = 10'd465;
b_exp0 = 10'd367; b_exp1 = 10'd514; b_exp2 = 10'd795; b_exp3 = 10'd572;
a_sign0 = 4'd4; a_sign1 = 4'd6; a_sign2 = 4'd4; a_sign3 = 4'd8;
b_sign0 = 4'd10; b_sign1 = 4'd6; b_sign2 = 4'd12; b_sign3 = 4'd15;
@(posedge clk_i);
a_mant0 = 8'd167; a_mant1 = 8'd37; a_mant2 = 8'd7; a_mant3 = 8'd25;
b_mant0 = 8'd139; b_mant1 = 8'd39; b_mant2 = 8'd190; b_mant3 = 8'd249;
a_exp0 = 10'd473; a_exp1 = 10'd227; a_exp2 = 10'd414; a_exp3 = 10'd129;
b_exp0 = 10'd410; b_exp1 = 10'd851; b_exp2 = 10'd449; b_exp3 = 10'd287;
a_sign0 = 4'd11; a_sign1 = 4'd13; a_sign2 = 4'd14; a_sign3 = 4'd16;
b_sign0 = 4'd3; b_sign1 = 4'd12; b_sign2 = 4'd10; b_sign3 = 4'd5;
@(posedge clk_i);
a_mant0 = 8'd40; a_mant1 = 8'd128; a_mant2 = 8'd147; a_mant3 = 8'd135;
b_mant0 = 8'd166; b_mant1 = 8'd21; b_mant2 = 8'd48; b_mant3 = 8'd223;
a_exp0 = 10'd384; a_exp1 = 10'd209; a_exp2 = 10'd264; a_exp3 = 10'd809;
b_exp0 = 10'd597; b_exp1 = 10'd255; b_exp2 = 10'd507; b_exp3 = 10'd739;
a_sign0 = 4'd10; a_sign1 = 4'd12; a_sign2 = 4'd14; a_sign3 = 4'd0;
b_sign0 = 4'd14; b_sign1 = 4'd4; b_sign2 = 4'd10; b_sign3 = 4'd13;
@(posedge clk_i);
a_mant0 = 8'd6; a_mant1 = 8'd102; a_mant2 = 8'd118; a_mant3 = 8'd168;
b_mant0 = 8'd18; b_mant1 = 8'd147; b_mant2 = 8'd84; b_mant3 = 8'd107;
a_exp0 = 10'd739; a_exp1 = 10'd336; a_exp2 = 10'd176; a_exp3 = 10'd390;
b_exp0 = 10'd1006; b_exp1 = 10'd1017; b_exp2 = 10'd837; b_exp3 = 10'd748;
a_sign0 = 4'd12; a_sign1 = 4'd12; a_sign2 = 4'd16; a_sign3 = 4'd16;
b_sign0 = 4'd15; b_sign1 = 4'd11; b_sign2 = 4'd14; b_sign3 = 4'd13;
@(posedge clk_i);
a_mant0 = 8'd181; a_mant1 = 8'd200; a_mant2 = 8'd142; a_mant3 = 8'd162;
b_mant0 = 8'd149; b_mant1 = 8'd93; b_mant2 = 8'd58; b_mant3 = 8'd94;
a_exp0 = 10'd907; a_exp1 = 10'd822; a_exp2 = 10'd418; a_exp3 = 10'd841;
b_exp0 = 10'd180; b_exp1 = 10'd74; b_exp2 = 10'd55; b_exp3 = 10'd936;
a_sign0 = 4'd9; a_sign1 = 4'd0; a_sign2 = 4'd7; a_sign3 = 4'd0;
b_sign0 = 4'd7; b_sign1 = 4'd14; b_sign2 = 4'd14; b_sign3 = 4'd6;
@(posedge clk_i);
a_mant0 = 8'd243; a_mant1 = 8'd253; a_mant2 = 8'd200; a_mant3 = 8'd54;
b_mant0 = 8'd178; b_mant1 = 8'd124; b_mant2 = 8'd19; b_mant3 = 8'd54;
a_exp0 = 10'd839; a_exp1 = 10'd179; a_exp2 = 10'd110; a_exp3 = 10'd52;
b_exp0 = 10'd121; b_exp1 = 10'd65; b_exp2 = 10'd326; b_exp3 = 10'd257;
a_sign0 = 4'd2; a_sign1 = 4'd13; a_sign2 = 4'd10; a_sign3 = 4'd3;
b_sign0 = 4'd15; b_sign1 = 4'd2; b_sign2 = 4'd12; b_sign3 = 4'd2;
@(posedge clk_i);
shared_exps0 = 8'd130;
shared_exps1 = 8'd118;
a_mant0 = 8'd198; a_mant1 = 8'd119; a_mant2 = 8'd3; a_mant3 = 8'd233;
b_mant0 = 8'd239; b_mant1 = 8'd242; b_mant2 = 8'd118; b_mant3 = 8'd214;
a_exp0 = 10'd83; a_exp1 = 10'd233; a_exp2 = 10'd785; a_exp3 = 10'd507;
b_exp0 = 10'd486; b_exp1 = 10'd759; b_exp2 = 10'd101; b_exp3 = 10'd818;
a_sign0 = 4'd7; a_sign1 = 4'd6; a_sign2 = 4'd7; a_sign3 = 4'd15;
b_sign0 = 4'd2; b_sign1 = 4'd8; b_sign2 = 4'd5; b_sign3 = 4'd2;
@(posedge clk_i);
a_mant0 = 8'd199; a_mant1 = 8'd11; a_mant2 = 8'd254; a_mant3 = 8'd4;
b_mant0 = 8'd144; b_mant1 = 8'd51; b_mant2 = 8'd213; b_mant3 = 8'd233;
a_exp0 = 10'd671; a_exp1 = 10'd146; a_exp2 = 10'd79; a_exp3 = 10'd761;
b_exp0 = 10'd935; b_exp1 = 10'd334; b_exp2 = 10'd34; b_exp3 = 10'd502;
a_sign0 = 4'd9; a_sign1 = 4'd7; a_sign2 = 4'd4; a_sign3 = 4'd9;
b_sign0 = 4'd14; b_sign1 = 4'd15; b_sign2 = 4'd11; b_sign3 = 4'd12;
@(posedge clk_i);
a_mant0 = 8'd64; a_mant1 = 8'd235; a_mant2 = 8'd217; a_mant3 = 8'd1;
b_mant0 = 8'd196; b_mant1 = 8'd31; b_mant2 = 8'd19; b_mant3 = 8'd216;
a_exp0 = 10'd155; a_exp1 = 10'd340; a_exp2 = 10'd821; a_exp3 = 10'd103;
b_exp0 = 10'd175; b_exp1 = 10'd417; b_exp2 = 10'd555; b_exp3 = 10'd216;
a_sign0 = 4'd16; a_sign1 = 4'd2; a_sign2 = 4'd15; a_sign3 = 4'd3;
b_sign0 = 4'd5; b_sign1 = 4'd8; b_sign2 = 4'd7; b_sign3 = 4'd10;
@(posedge clk_i);
a_mant0 = 8'd80; a_mant1 = 8'd22; a_mant2 = 8'd85; a_mant3 = 8'd12;
b_mant0 = 8'd85; b_mant1 = 8'd125; b_mant2 = 8'd207; b_mant3 = 8'd145;
a_exp0 = 10'd589; a_exp1 = 10'd1012; a_exp2 = 10'd988; a_exp3 = 10'd814;
b_exp0 = 10'd288; b_exp1 = 10'd115; b_exp2 = 10'd36; b_exp3 = 10'd297;
a_sign0 = 4'd13; a_sign1 = 4'd1; a_sign2 = 4'd4; a_sign3 = 4'd12;
b_sign0 = 4'd1; b_sign1 = 4'd3; b_sign2 = 4'd15; b_sign3 = 4'd8;
@(posedge clk_i);
a_mant0 = 8'd207; a_mant1 = 8'd183; a_mant2 = 8'd80; a_mant3 = 8'd180;
b_mant0 = 8'd83; b_mant1 = 8'd217; b_mant2 = 8'd48; b_mant3 = 8'd102;
a_exp0 = 10'd78; a_exp1 = 10'd870; a_exp2 = 10'd832; a_exp3 = 10'd128;
b_exp0 = 10'd505; b_exp1 = 10'd482; b_exp2 = 10'd718; b_exp3 = 10'd90;
a_sign0 = 4'd11; a_sign1 = 4'd14; a_sign2 = 4'd8; a_sign3 = 4'd9;
b_sign0 = 4'd14; b_sign1 = 4'd11; b_sign2 = 4'd16; b_sign3 = 4'd16;
@(posedge clk_i);
a_mant0 = 8'd215; a_mant1 = 8'd203; a_mant2 = 8'd143; a_mant3 = 8'd60;
b_mant0 = 8'd28; b_mant1 = 8'd96; b_mant2 = 8'd151; b_mant3 = 8'd237;
a_exp0 = 10'd926; a_exp1 = 10'd88; a_exp2 = 10'd797; a_exp3 = 10'd572;
b_exp0 = 10'd236; b_exp1 = 10'd294; b_exp2 = 10'd21; b_exp3 = 10'd921;
a_sign0 = 4'd6; a_sign1 = 4'd15; a_sign2 = 4'd3; a_sign3 = 4'd0;
b_sign0 = 4'd4; b_sign1 = 4'd15; b_sign2 = 4'd9; b_sign3 = 4'd2;
@(posedge clk_i);
a_mant0 = 8'd159; a_mant1 = 8'd181; a_mant2 = 8'd3; a_mant3 = 8'd209;
b_mant0 = 8'd128; b_mant1 = 8'd192; b_mant2 = 8'd0; b_mant3 = 8'd18;
a_exp0 = 10'd859; a_exp1 = 10'd987; a_exp2 = 10'd2; a_exp3 = 10'd697;
b_exp0 = 10'd313; b_exp1 = 10'd536; b_exp2 = 10'd955; b_exp3 = 10'd262;
a_sign0 = 4'd11; a_sign1 = 4'd1; a_sign2 = 4'd2; a_sign3 = 4'd8;
b_sign0 = 4'd0; b_sign1 = 4'd10; b_sign2 = 4'd10; b_sign3 = 4'd9;
@(posedge clk_i);
a_mant0 = 8'd112; a_mant1 = 8'd170; a_mant2 = 8'd214; a_mant3 = 8'd16;
b_mant0 = 8'd110; b_mant1 = 8'd161; b_mant2 = 8'd68; b_mant3 = 8'd60;
a_exp0 = 10'd573; a_exp1 = 10'd45; a_exp2 = 10'd442; a_exp3 = 10'd10;
b_exp0 = 10'd931; b_exp1 = 10'd718; b_exp2 = 10'd310; b_exp3 = 10'd206;
a_sign0 = 4'd6; a_sign1 = 4'd1; a_sign2 = 4'd6; a_sign3 = 4'd2;
b_sign0 = 4'd9; b_sign1 = 4'd7; b_sign2 = 4'd6; b_sign3 = 4'd16;
@(posedge clk_i);
shared_exps0 = 8'd123;
shared_exps1 = 8'd152;
a_mant0 = 8'd3; a_mant1 = 8'd237; a_mant2 = 8'd36; a_mant3 = 8'd78;
b_mant0 = 8'd188; b_mant1 = 8'd43; b_mant2 = 8'd86; b_mant3 = 8'd230;
a_exp0 = 10'd990; a_exp1 = 10'd657; a_exp2 = 10'd706; a_exp3 = 10'd286;
b_exp0 = 10'd45; b_exp1 = 10'd962; b_exp2 = 10'd594; b_exp3 = 10'd546;
a_sign0 = 4'd1; a_sign1 = 4'd11; a_sign2 = 4'd15; a_sign3 = 4'd1;
b_sign0 = 4'd6; b_sign1 = 4'd15; b_sign2 = 4'd11; b_sign3 = 4'd2;
@(posedge clk_i);
a_mant0 = 8'd19; a_mant1 = 8'd146; a_mant2 = 8'd111; a_mant3 = 8'd150;
b_mant0 = 8'd43; b_mant1 = 8'd14; b_mant2 = 8'd45; b_mant3 = 8'd242;
a_exp0 = 10'd92; a_exp1 = 10'd424; a_exp2 = 10'd314; a_exp3 = 10'd721;
b_exp0 = 10'd641; b_exp1 = 10'd975; b_exp2 = 10'd253; b_exp3 = 10'd113;
a_sign0 = 4'd4; a_sign1 = 4'd8; a_sign2 = 4'd12; a_sign3 = 4'd7;
b_sign0 = 4'd13; b_sign1 = 4'd6; b_sign2 = 4'd16; b_sign3 = 4'd10;
@(posedge clk_i);
a_mant0 = 8'd253; a_mant1 = 8'd184; a_mant2 = 8'd120; a_mant3 = 8'd66;
b_mant0 = 8'd138; b_mant1 = 8'd238; b_mant2 = 8'd51; b_mant3 = 8'd233;
a_exp0 = 10'd566; a_exp1 = 10'd11; a_exp2 = 10'd434; a_exp3 = 10'd628;
b_exp0 = 10'd661; b_exp1 = 10'd778; b_exp2 = 10'd715; b_exp3 = 10'd184;
a_sign0 = 4'd4; a_sign1 = 4'd7; a_sign2 = 4'd7; a_sign3 = 4'd12;
b_sign0 = 4'd2; b_sign1 = 4'd5; b_sign2 = 4'd3; b_sign3 = 4'd1;
@(posedge clk_i);
a_mant0 = 8'd31; a_mant1 = 8'd197; a_mant2 = 8'd104; a_mant3 = 8'd63;
b_mant0 = 8'd116; b_mant1 = 8'd173; b_mant2 = 8'd103; b_mant3 = 8'd158;
a_exp0 = 10'd836; a_exp1 = 10'd361; a_exp2 = 10'd636; a_exp3 = 10'd140;
b_exp0 = 10'd989; b_exp1 = 10'd433; b_exp2 = 10'd972; b_exp3 = 10'd25;
a_sign0 = 4'd14; a_sign1 = 4'd15; a_sign2 = 4'd8; a_sign3 = 4'd2;
b_sign0 = 4'd15; b_sign1 = 4'd14; b_sign2 = 4'd7; b_sign3 = 4'd13;
@(posedge clk_i);
a_mant0 = 8'd7; a_mant1 = 8'd92; a_mant2 = 8'd73; a_mant3 = 8'd58;
b_mant0 = 8'd2; b_mant1 = 8'd54; b_mant2 = 8'd231; b_mant3 = 8'd250;
a_exp0 = 10'd305; a_exp1 = 10'd255; a_exp2 = 10'd85; a_exp3 = 10'd294;
b_exp0 = 10'd746; b_exp1 = 10'd681; b_exp2 = 10'd588; b_exp3 = 10'd792;
a_sign0 = 4'd11; a_sign1 = 4'd15; a_sign2 = 4'd8; a_sign3 = 4'd14;
b_sign0 = 4'd4; b_sign1 = 4'd14; b_sign2 = 4'd3; b_sign3 = 4'd3;
@(posedge clk_i);
a_mant0 = 8'd72; a_mant1 = 8'd250; a_mant2 = 8'd39; a_mant3 = 8'd104;
b_mant0 = 8'd140; b_mant1 = 8'd52; b_mant2 = 8'd214; b_mant3 = 8'd147;
a_exp0 = 10'd254; a_exp1 = 10'd632; a_exp2 = 10'd880; a_exp3 = 10'd610;
b_exp0 = 10'd364; b_exp1 = 10'd726; b_exp2 = 10'd729; b_exp3 = 10'd599;
a_sign0 = 4'd13; a_sign1 = 4'd8; a_sign2 = 4'd1; a_sign3 = 4'd10;
b_sign0 = 4'd2; b_sign1 = 4'd8; b_sign2 = 4'd14; b_sign3 = 4'd9;
@(posedge clk_i);
a_mant0 = 8'd188; a_mant1 = 8'd11; a_mant2 = 8'd251; a_mant3 = 8'd85;
b_mant0 = 8'd188; b_mant1 = 8'd238; b_mant2 = 8'd95; b_mant3 = 8'd233;
a_exp0 = 10'd139; a_exp1 = 10'd2; a_exp2 = 10'd292; a_exp3 = 10'd485;
b_exp0 = 10'd680; b_exp1 = 10'd706; b_exp2 = 10'd142; b_exp3 = 10'd960;
a_sign0 = 4'd3; a_sign1 = 4'd11; a_sign2 = 4'd6; a_sign3 = 4'd1;
b_sign0 = 4'd6; b_sign1 = 4'd12; b_sign2 = 4'd8; b_sign3 = 4'd16;
@(posedge clk_i);
a_mant0 = 8'd169; a_mant1 = 8'd180; a_mant2 = 8'd120; a_mant3 = 8'd167;
b_mant0 = 8'd130; b_mant1 = 8'd154; b_mant2 = 8'd51; b_mant3 = 8'd171;
a_exp0 = 10'd538; a_exp1 = 10'd815; a_exp2 = 10'd388; a_exp3 = 10'd866;
b_exp0 = 10'd594; b_exp1 = 10'd887; b_exp2 = 10'd527; b_exp3 = 10'd124;
a_sign0 = 4'd11; a_sign1 = 4'd11; a_sign2 = 4'd16; a_sign3 = 4'd11;
b_sign0 = 4'd8; b_sign1 = 4'd15; b_sign2 = 4'd14; b_sign3 = 4'd6;
@(posedge clk_i);
shared_exps0 = 8'd116;
shared_exps1 = 8'd142;
rstn = 0;
@(posedge clk_i);
rstn = 1;
a_mant0 = 8'd81; a_mant1 = 8'd48; a_mant2 = 8'd224; a_mant3 = 8'd69;
b_mant0 = 8'd16; b_mant1 = 8'd93; b_mant2 = 8'd39; b_mant3 = 8'd73;
a_exp0 = 10'd21; a_exp1 = 10'd261; a_exp2 = 10'd144; a_exp3 = 10'd473;
b_exp0 = 10'd364; b_exp1 = 10'd835; b_exp2 = 10'd71; b_exp3 = 10'd869;
a_sign0 = 4'd1; a_sign1 = 4'd0; a_sign2 = 4'd11; a_sign3 = 4'd1;
b_sign0 = 4'd7; b_sign1 = 4'd10; b_sign2 = 4'd7; b_sign3 = 4'd6;
@(posedge clk_i);
a_mant0 = 8'd174; a_mant1 = 8'd198; a_mant2 = 8'd25; a_mant3 = 8'd157;
b_mant0 = 8'd43; b_mant1 = 8'd60; b_mant2 = 8'd96; b_mant3 = 8'd109;
a_exp0 = 10'd530; a_exp1 = 10'd319; a_exp2 = 10'd1004; a_exp3 = 10'd578;
b_exp0 = 10'd277; b_exp1 = 10'd980; b_exp2 = 10'd355; b_exp3 = 10'd615;
a_sign0 = 4'd15; a_sign1 = 4'd12; a_sign2 = 4'd7; a_sign3 = 4'd5;
b_sign0 = 4'd6; b_sign1 = 4'd8; b_sign2 = 4'd4; b_sign3 = 4'd6;
@(posedge clk_i);
a_mant0 = 8'd78; a_mant1 = 8'd129; a_mant2 = 8'd176; a_mant3 = 8'd235;
b_mant0 = 8'd75; b_mant1 = 8'd20; b_mant2 = 8'd39; b_mant3 = 8'd99;
a_exp0 = 10'd703; a_exp1 = 10'd630; a_exp2 = 10'd704; a_exp3 = 10'd378;
b_exp0 = 10'd75; b_exp1 = 10'd13; b_exp2 = 10'd377; b_exp3 = 10'd402;
a_sign0 = 4'd13; a_sign1 = 4'd9; a_sign2 = 4'd3; a_sign3 = 4'd12;
b_sign0 = 4'd6; b_sign1 = 4'd0; b_sign2 = 4'd13; b_sign3 = 4'd8;
@(posedge clk_i);
a_mant0 = 8'd52; a_mant1 = 8'd57; a_mant2 = 8'd44; a_mant3 = 8'd197;
b_mant0 = 8'd182; b_mant1 = 8'd145; b_mant2 = 8'd113; b_mant3 = 8'd173;
a_exp0 = 10'd278; a_exp1 = 10'd233; a_exp2 = 10'd942; a_exp3 = 10'd343;
b_exp0 = 10'd2; b_exp1 = 10'd269; b_exp2 = 10'd307; b_exp3 = 10'd110;
a_sign0 = 4'd10; a_sign1 = 4'd12; a_sign2 = 4'd13; a_sign3 = 4'd6;
b_sign0 = 4'd10; b_sign1 = 4'd9; b_sign2 = 4'd13; b_sign3 = 4'd7;
@(posedge clk_i);
a_mant0 = 8'd10; a_mant1 = 8'd73; a_mant2 = 8'd170; a_mant3 = 8'd5;
b_mant0 = 8'd176; b_mant1 = 8'd245; b_mant2 = 8'd165; b_mant3 = 8'd242;
a_exp0 = 10'd396; a_exp1 = 10'd306; a_exp2 = 10'd616; a_exp3 = 10'd603;
b_exp0 = 10'd784; b_exp1 = 10'd646; b_exp2 = 10'd503; b_exp3 = 10'd113;
a_sign0 = 4'd8; a_sign1 = 4'd12; a_sign2 = 4'd13; a_sign3 = 4'd12;
b_sign0 = 4'd6; b_sign1 = 4'd11; b_sign2 = 4'd14; b_sign3 = 4'd11;
@(posedge clk_i);
a_mant0 = 8'd70; a_mant1 = 8'd85; a_mant2 = 8'd186; a_mant3 = 8'd229;
b_mant0 = 8'd176; b_mant1 = 8'd182; b_mant2 = 8'd243; b_mant3 = 8'd83;
a_exp0 = 10'd405; a_exp1 = 10'd609; a_exp2 = 10'd423; a_exp3 = 10'd623;
b_exp0 = 10'd92; b_exp1 = 10'd561; b_exp2 = 10'd85; b_exp3 = 10'd794;
a_sign0 = 4'd16; a_sign1 = 4'd16; a_sign2 = 4'd11; a_sign3 = 4'd11;
b_sign0 = 4'd6; b_sign1 = 4'd3; b_sign2 = 4'd12; b_sign3 = 4'd13;
@(posedge clk_i);
a_mant0 = 8'd44; a_mant1 = 8'd90; a_mant2 = 8'd254; a_mant3 = 8'd240;
b_mant0 = 8'd13; b_mant1 = 8'd44; b_mant2 = 8'd149; b_mant3 = 8'd122;
a_exp0 = 10'd172; a_exp1 = 10'd130; a_exp2 = 10'd540; a_exp3 = 10'd162;
b_exp0 = 10'd662; b_exp1 = 10'd811; b_exp2 = 10'd1011; b_exp3 = 10'd107;
a_sign0 = 4'd13; a_sign1 = 4'd10; a_sign2 = 4'd13; a_sign3 = 4'd15;
b_sign0 = 4'd5; b_sign1 = 4'd12; b_sign2 = 4'd12; b_sign3 = 4'd4;
@(posedge clk_i);
shared_exps0 = 8'd114;
shared_exps1 = 8'd124;
a_mant0 = 8'd234; a_mant1 = 8'd59; a_mant2 = 8'd134; a_mant3 = 8'd200;
b_mant0 = 8'd81; b_mant1 = 8'd236; b_mant2 = 8'd45; b_mant3 = 8'd10;
a_exp0 = 10'd401; a_exp1 = 10'd32; a_exp2 = 10'd686; a_exp3 = 10'd1004;
b_exp0 = 10'd341; b_exp1 = 10'd259; b_exp2 = 10'd166; b_exp3 = 10'd848;
a_sign0 = 4'd16; a_sign1 = 4'd11; a_sign2 = 4'd12; a_sign3 = 4'd8;
b_sign0 = 4'd1; b_sign1 = 4'd11; b_sign2 = 4'd0; b_sign3 = 4'd11;
@(posedge clk_i);
a_mant0 = 8'd204; a_mant1 = 8'd106; a_mant2 = 8'd248; a_mant3 = 8'd239;
b_mant0 = 8'd160; b_mant1 = 8'd63; b_mant2 = 8'd103; b_mant3 = 8'd155;
a_exp0 = 10'd905; a_exp1 = 10'd720; a_exp2 = 10'd906; a_exp3 = 10'd921;
b_exp0 = 10'd714; b_exp1 = 10'd372; b_exp2 = 10'd673; b_exp3 = 10'd923;
a_sign0 = 4'd0; a_sign1 = 4'd1; a_sign2 = 4'd8; a_sign3 = 4'd13;
b_sign0 = 4'd3; b_sign1 = 4'd15; b_sign2 = 4'd10; b_sign3 = 4'd0;
@(posedge clk_i);
a_mant0 = 8'd26; a_mant1 = 8'd228; a_mant2 = 8'd121; a_mant3 = 8'd153;
b_mant0 = 8'd135; b_mant1 = 8'd37; b_mant2 = 8'd94; b_mant3 = 8'd230;
a_exp0 = 10'd437; a_exp1 = 10'd902; a_exp2 = 10'd8; a_exp3 = 10'd101;
b_exp0 = 10'd965; b_exp1 = 10'd64; b_exp2 = 10'd548; b_exp3 = 10'd891;
a_sign0 = 4'd8; a_sign1 = 4'd10; a_sign2 = 4'd7; a_sign3 = 4'd0;
b_sign0 = 4'd7; b_sign1 = 4'd7; b_sign2 = 4'd5; b_sign3 = 4'd4;
@(posedge clk_i);
a_mant0 = 8'd165; a_mant1 = 8'd101; a_mant2 = 8'd226; a_mant3 = 8'd219;
b_mant0 = 8'd156; b_mant1 = 8'd71; b_mant2 = 8'd249; b_mant3 = 8'd116;
a_exp0 = 10'd443; a_exp1 = 10'd461; a_exp2 = 10'd384; a_exp3 = 10'd790;
b_exp0 = 10'd95; b_exp1 = 10'd84; b_exp2 = 10'd709; b_exp3 = 10'd535;
a_sign0 = 4'd6; a_sign1 = 4'd7; a_sign2 = 4'd10; a_sign3 = 4'd7;
b_sign0 = 4'd10; b_sign1 = 4'd15; b_sign2 = 4'd4; b_sign3 = 4'd4;
@(posedge clk_i);
a_mant0 = 8'd107; a_mant1 = 8'd229; a_mant2 = 8'd126; a_mant3 = 8'd71;
b_mant0 = 8'd23; b_mant1 = 8'd18; b_mant2 = 8'd129; b_mant3 = 8'd37;
a_exp0 = 10'd131; a_exp1 = 10'd924; a_exp2 = 10'd750; a_exp3 = 10'd159;
b_exp0 = 10'd210; b_exp1 = 10'd74; b_exp2 = 10'd56; b_exp3 = 10'd127;
a_sign0 = 4'd10; a_sign1 = 4'd13; a_sign2 = 4'd1; a_sign3 = 4'd2;
b_sign0 = 4'd4; b_sign1 = 4'd2; b_sign2 = 4'd9; b_sign3 = 4'd5;
@(posedge clk_i);
a_mant0 = 8'd199; a_mant1 = 8'd244; a_mant2 = 8'd203; a_mant3 = 8'd217;
b_mant0 = 8'd41; b_mant1 = 8'd32; b_mant2 = 8'd34; b_mant3 = 8'd23;
a_exp0 = 10'd272; a_exp1 = 10'd138; a_exp2 = 10'd246; a_exp3 = 10'd611;
b_exp0 = 10'd366; b_exp1 = 10'd976; b_exp2 = 10'd699; b_exp3 = 10'd851;
a_sign0 = 4'd0; a_sign1 = 4'd16; a_sign2 = 4'd14; a_sign3 = 4'd15;
b_sign0 = 4'd5; b_sign1 = 4'd0; b_sign2 = 4'd4; b_sign3 = 4'd8;
@(posedge clk_i);
a_mant0 = 8'd126; a_mant1 = 8'd187; a_mant2 = 8'd35; a_mant3 = 8'd208;
b_mant0 = 8'd115; b_mant1 = 8'd165; b_mant2 = 8'd43; b_mant3 = 8'd17;
a_exp0 = 10'd307; a_exp1 = 10'd558; a_exp2 = 10'd84; a_exp3 = 10'd171;
b_exp0 = 10'd855; b_exp1 = 10'd505; b_exp2 = 10'd541; b_exp3 = 10'd739;
a_sign0 = 4'd8; a_sign1 = 4'd8; a_sign2 = 4'd16; a_sign3 = 4'd13;
b_sign0 = 4'd8; b_sign1 = 4'd7; b_sign2 = 4'd14; b_sign3 = 4'd16;
@(posedge clk_i);
a_mant0 = 8'd15; a_mant1 = 8'd56; a_mant2 = 8'd168; a_mant3 = 8'd83;
b_mant0 = 8'd101; b_mant1 = 8'd123; b_mant2 = 8'd146; b_mant3 = 8'd122;
a_exp0 = 10'd729; a_exp1 = 10'd568; a_exp2 = 10'd111; a_exp3 = 10'd300;
b_exp0 = 10'd226; b_exp1 = 10'd411; b_exp2 = 10'd716; b_exp3 = 10'd444;
a_sign0 = 4'd9; a_sign1 = 4'd5; a_sign2 = 4'd5; a_sign3 = 4'd7;
b_sign0 = 4'd8; b_sign1 = 4'd3; b_sign2 = 4'd3; b_sign3 = 4'd4;
@(posedge clk_i);
shared_exps0 = 8'd150;
shared_exps1 = 8'd144;
a_mant0 = 8'd42; a_mant1 = 8'd38; a_mant2 = 8'd155; a_mant3 = 8'd138;
b_mant0 = 8'd28; b_mant1 = 8'd208; b_mant2 = 8'd148; b_mant3 = 8'd50;
a_exp0 = 10'd965; a_exp1 = 10'd496; a_exp2 = 10'd294; a_exp3 = 10'd178;
b_exp0 = 10'd69; b_exp1 = 10'd659; b_exp2 = 10'd590; b_exp3 = 10'd723;
a_sign0 = 4'd3; a_sign1 = 4'd3; a_sign2 = 4'd0; a_sign3 = 4'd7;
b_sign0 = 4'd8; b_sign1 = 4'd15; b_sign2 = 4'd8; b_sign3 = 4'd16;
@(posedge clk_i);
a_mant0 = 8'd60; a_mant1 = 8'd3; a_mant2 = 8'd222; a_mant3 = 8'd235;
b_mant0 = 8'd142; b_mant1 = 8'd9; b_mant2 = 8'd175; b_mant3 = 8'd125;
a_exp0 = 10'd282; a_exp1 = 10'd500; a_exp2 = 10'd977; a_exp3 = 10'd1008;
b_exp0 = 10'd163; b_exp1 = 10'd495; b_exp2 = 10'd249; b_exp3 = 10'd261;
a_sign0 = 4'd4; a_sign1 = 4'd15; a_sign2 = 4'd1; a_sign3 = 4'd13;
b_sign0 = 4'd9; b_sign1 = 4'd3; b_sign2 = 4'd4; b_sign3 = 4'd8;
@(posedge clk_i);
a_mant0 = 8'd121; a_mant1 = 8'd137; a_mant2 = 8'd234; a_mant3 = 8'd140;
b_mant0 = 8'd149; b_mant1 = 8'd53; b_mant2 = 8'd132; b_mant3 = 8'd215;
a_exp0 = 10'd514; a_exp1 = 10'd653; a_exp2 = 10'd269; a_exp3 = 10'd56;
b_exp0 = 10'd715; b_exp1 = 10'd141; b_exp2 = 10'd423; b_exp3 = 10'd368;
a_sign0 = 4'd12; a_sign1 = 4'd0; a_sign2 = 4'd1; a_sign3 = 4'd2;
b_sign0 = 4'd15; b_sign1 = 4'd0; b_sign2 = 4'd14; b_sign3 = 4'd1;
@(posedge clk_i);
a_mant0 = 8'd64; a_mant1 = 8'd127; a_mant2 = 8'd21; a_mant3 = 8'd36;
b_mant0 = 8'd180; b_mant1 = 8'd28; b_mant2 = 8'd233; b_mant3 = 8'd122;
a_exp0 = 10'd612; a_exp1 = 10'd427; a_exp2 = 10'd499; a_exp3 = 10'd650;
b_exp0 = 10'd1019; b_exp1 = 10'd539; b_exp2 = 10'd210; b_exp3 = 10'd657;
a_sign0 = 4'd4; a_sign1 = 4'd9; a_sign2 = 4'd12; a_sign3 = 4'd7;
b_sign0 = 4'd10; b_sign1 = 4'd8; b_sign2 = 4'd10; b_sign3 = 4'd6;
@(posedge clk_i);
a_mant0 = 8'd143; a_mant1 = 8'd79; a_mant2 = 8'd82; a_mant3 = 8'd139;
b_mant0 = 8'd166; b_mant1 = 8'd44; b_mant2 = 8'd38; b_mant3 = 8'd240;
a_exp0 = 10'd44; a_exp1 = 10'd607; a_exp2 = 10'd171; a_exp3 = 10'd594;
b_exp0 = 10'd420; b_exp1 = 10'd967; b_exp2 = 10'd126; b_exp3 = 10'd392;
a_sign0 = 4'd2; a_sign1 = 4'd12; a_sign2 = 4'd16; a_sign3 = 4'd11;
b_sign0 = 4'd7; b_sign1 = 4'd13; b_sign2 = 4'd15; b_sign3 = 4'd16;
@(posedge clk_i);
a_mant0 = 8'd223; a_mant1 = 8'd87; a_mant2 = 8'd193; a_mant3 = 8'd131;
b_mant0 = 8'd181; b_mant1 = 8'd49; b_mant2 = 8'd16; b_mant3 = 8'd89;
a_exp0 = 10'd286; a_exp1 = 10'd552; a_exp2 = 10'd779; a_exp3 = 10'd212;
b_exp0 = 10'd77; b_exp1 = 10'd182; b_exp2 = 10'd548; b_exp3 = 10'd486;
a_sign0 = 4'd4; a_sign1 = 4'd8; a_sign2 = 4'd3; a_sign3 = 4'd1;
b_sign0 = 4'd2; b_sign1 = 4'd3; b_sign2 = 4'd13; b_sign3 = 4'd2;
@(posedge clk_i);
a_mant0 = 8'd142; a_mant1 = 8'd6; a_mant2 = 8'd215; a_mant3 = 8'd245;
b_mant0 = 8'd208; b_mant1 = 8'd133; b_mant2 = 8'd83; b_mant3 = 8'd35;
a_exp0 = 10'd44; a_exp1 = 10'd319; a_exp2 = 10'd629; a_exp3 = 10'd844;
b_exp0 = 10'd883; b_exp1 = 10'd148; b_exp2 = 10'd32; b_exp3 = 10'd571;
a_sign0 = 4'd5; a_sign1 = 4'd12; a_sign2 = 4'd16; a_sign3 = 4'd11;
b_sign0 = 4'd2; b_sign1 = 4'd0; b_sign2 = 4'd6; b_sign3 = 4'd11;
@(posedge clk_i);
a_mant0 = 8'd115; a_mant1 = 8'd12; a_mant2 = 8'd170; a_mant3 = 8'd210;
b_mant0 = 8'd134; b_mant1 = 8'd37; b_mant2 = 8'd231; b_mant3 = 8'd145;
a_exp0 = 10'd451; a_exp1 = 10'd59; a_exp2 = 10'd214; a_exp3 = 10'd335;
b_exp0 = 10'd401; b_exp1 = 10'd77; b_exp2 = 10'd109; b_exp3 = 10'd609;
a_sign0 = 4'd14; a_sign1 = 4'd0; a_sign2 = 4'd16; a_sign3 = 4'd15;
b_sign0 = 4'd14; b_sign1 = 4'd5; b_sign2 = 4'd9; b_sign3 = 4'd8;
@(posedge clk_i);
shared_exps0 = 8'd117;
shared_exps1 = 8'd149;
a_mant0 = 8'd58; a_mant1 = 8'd103; a_mant2 = 8'd118; a_mant3 = 8'd38;
b_mant0 = 8'd71; b_mant1 = 8'd245; b_mant2 = 8'd138; b_mant3 = 8'd149;
a_exp0 = 10'd933; a_exp1 = 10'd1014; a_exp2 = 10'd651; a_exp3 = 10'd215;
b_exp0 = 10'd925; b_exp1 = 10'd340; b_exp2 = 10'd541; b_exp3 = 10'd134;
a_sign0 = 4'd16; a_sign1 = 4'd16; a_sign2 = 4'd1; a_sign3 = 4'd4;
b_sign0 = 4'd7; b_sign1 = 4'd1; b_sign2 = 4'd14; b_sign3 = 4'd8;
@(posedge clk_i);
a_mant0 = 8'd117; a_mant1 = 8'd131; a_mant2 = 8'd99; a_mant3 = 8'd207;
b_mant0 = 8'd205; b_mant1 = 8'd127; b_mant2 = 8'd27; b_mant3 = 8'd198;
a_exp0 = 10'd630; a_exp1 = 10'd508; a_exp2 = 10'd805; a_exp3 = 10'd36;
b_exp0 = 10'd164; b_exp1 = 10'd341; b_exp2 = 10'd401; b_exp3 = 10'd531;
a_sign0 = 4'd0; a_sign1 = 4'd3; a_sign2 = 4'd16; a_sign3 = 4'd13;
b_sign0 = 4'd16; b_sign1 = 4'd5; b_sign2 = 4'd3; b_sign3 = 4'd2;
@(posedge clk_i);
a_mant0 = 8'd223; a_mant1 = 8'd20; a_mant2 = 8'd107; a_mant3 = 8'd199;
b_mant0 = 8'd30; b_mant1 = 8'd229; b_mant2 = 8'd74; b_mant3 = 8'd107;
a_exp0 = 10'd857; a_exp1 = 10'd274; a_exp2 = 10'd375; a_exp3 = 10'd274;
b_exp0 = 10'd1012; b_exp1 = 10'd107; b_exp2 = 10'd712; b_exp3 = 10'd741;
a_sign0 = 4'd7; a_sign1 = 4'd12; a_sign2 = 4'd7; a_sign3 = 4'd15;
b_sign0 = 4'd10; b_sign1 = 4'd4; b_sign2 = 4'd9; b_sign3 = 4'd11;
@(posedge clk_i);
a_mant0 = 8'd199; a_mant1 = 8'd205; a_mant2 = 8'd103; a_mant3 = 8'd65;
b_mant0 = 8'd202; b_mant1 = 8'd195; b_mant2 = 8'd90; b_mant3 = 8'd190;
a_exp0 = 10'd139; a_exp1 = 10'd733; a_exp2 = 10'd790; a_exp3 = 10'd820;
b_exp0 = 10'd201; b_exp1 = 10'd481; b_exp2 = 10'd847; b_exp3 = 10'd596;
a_sign0 = 4'd7; a_sign1 = 4'd0; a_sign2 = 4'd0; a_sign3 = 4'd9;
b_sign0 = 4'd2; b_sign1 = 4'd1; b_sign2 = 4'd10; b_sign3 = 4'd3;
@(posedge clk_i);
a_mant0 = 8'd103; a_mant1 = 8'd131; a_mant2 = 8'd46; a_mant3 = 8'd152;
b_mant0 = 8'd135; b_mant1 = 8'd217; b_mant2 = 8'd11; b_mant3 = 8'd96;
a_exp0 = 10'd67; a_exp1 = 10'd810; a_exp2 = 10'd1020; a_exp3 = 10'd891;
b_exp0 = 10'd447; b_exp1 = 10'd984; b_exp2 = 10'd558; b_exp3 = 10'd501;
a_sign0 = 4'd1; a_sign1 = 4'd8; a_sign2 = 4'd0; a_sign3 = 4'd16;
b_sign0 = 4'd12; b_sign1 = 4'd9; b_sign2 = 4'd12; b_sign3 = 4'd10;
@(posedge clk_i);
a_mant0 = 8'd57; a_mant1 = 8'd78; a_mant2 = 8'd151; a_mant3 = 8'd206;
b_mant0 = 8'd118; b_mant1 = 8'd84; b_mant2 = 8'd162; b_mant3 = 8'd217;
a_exp0 = 10'd670; a_exp1 = 10'd356; a_exp2 = 10'd549; a_exp3 = 10'd543;
b_exp0 = 10'd766; b_exp1 = 10'd465; b_exp2 = 10'd616; b_exp3 = 10'd584;
a_sign0 = 4'd12; a_sign1 = 4'd8; a_sign2 = 4'd10; a_sign3 = 4'd12;
b_sign0 = 4'd8; b_sign1 = 4'd13; b_sign2 = 4'd1; b_sign3 = 4'd0;
@(posedge clk_i);
a_mant0 = 8'd212; a_mant1 = 8'd188; a_mant2 = 8'd19; a_mant3 = 8'd231;
b_mant0 = 8'd145; b_mant1 = 8'd233; b_mant2 = 8'd193; b_mant3 = 8'd1;
a_exp0 = 10'd686; a_exp1 = 10'd543; a_exp2 = 10'd13; a_exp3 = 10'd83;
b_exp0 = 10'd844; b_exp1 = 10'd39; b_exp2 = 10'd921; b_exp3 = 10'd93;
a_sign0 = 4'd1; a_sign1 = 4'd14; a_sign2 = 4'd5; a_sign3 = 4'd9;
b_sign0 = 4'd7; b_sign1 = 4'd14; b_sign2 = 4'd7; b_sign3 = 4'd1;
@(posedge clk_i);
a_mant0 = 8'd239; a_mant1 = 8'd62; a_mant2 = 8'd47; a_mant3 = 8'd160;
b_mant0 = 8'd43; b_mant1 = 8'd80; b_mant2 = 8'd172; b_mant3 = 8'd77;
a_exp0 = 10'd86; a_exp1 = 10'd652; a_exp2 = 10'd58; a_exp3 = 10'd764;
b_exp0 = 10'd933; b_exp1 = 10'd659; b_exp2 = 10'd802; b_exp3 = 10'd902;
a_sign0 = 4'd3; a_sign1 = 4'd3; a_sign2 = 4'd11; a_sign3 = 4'd2;
b_sign0 = 4'd9; b_sign1 = 4'd14; b_sign2 = 4'd13; b_sign3 = 4'd12;
@(posedge clk_i);
shared_exps0 = 8'd121;
shared_exps1 = 8'd136;
rstn = 0;
@(posedge clk_i);
rstn = 1;
a_mant0 = 8'd183; a_mant1 = 8'd242; a_mant2 = 8'd4; a_mant3 = 8'd175;
b_mant0 = 8'd220; b_mant1 = 8'd58; b_mant2 = 8'd150; b_mant3 = 8'd110;
a_exp0 = 10'd371; a_exp1 = 10'd654; a_exp2 = 10'd973; a_exp3 = 10'd1000;
b_exp0 = 10'd46; b_exp1 = 10'd797; b_exp2 = 10'd473; b_exp3 = 10'd896;
a_sign0 = 4'd3; a_sign1 = 4'd11; a_sign2 = 4'd9; a_sign3 = 4'd2;
b_sign0 = 4'd3; b_sign1 = 4'd8; b_sign2 = 4'd3; b_sign3 = 4'd11;
@(posedge clk_i);
a_mant0 = 8'd213; a_mant1 = 8'd59; a_mant2 = 8'd172; a_mant3 = 8'd228;
b_mant0 = 8'd75; b_mant1 = 8'd57; b_mant2 = 8'd13; b_mant3 = 8'd227;
a_exp0 = 10'd708; a_exp1 = 10'd856; a_exp2 = 10'd19; a_exp3 = 10'd323;
b_exp0 = 10'd962; b_exp1 = 10'd779; b_exp2 = 10'd204; b_exp3 = 10'd584;
a_sign0 = 4'd2; a_sign1 = 4'd14; a_sign2 = 4'd8; a_sign3 = 4'd2;
b_sign0 = 4'd15; b_sign1 = 4'd14; b_sign2 = 4'd9; b_sign3 = 4'd11;
@(posedge clk_i);
a_mant0 = 8'd214; a_mant1 = 8'd153; a_mant2 = 8'd174; a_mant3 = 8'd118;
b_mant0 = 8'd162; b_mant1 = 8'd253; b_mant2 = 8'd91; b_mant3 = 8'd231;
a_exp0 = 10'd443; a_exp1 = 10'd439; a_exp2 = 10'd701; a_exp3 = 10'd655;
b_exp0 = 10'd922; b_exp1 = 10'd180; b_exp2 = 10'd3; b_exp3 = 10'd214;
a_sign0 = 4'd13; a_sign1 = 4'd16; a_sign2 = 4'd15; a_sign3 = 4'd12;
b_sign0 = 4'd15; b_sign1 = 4'd14; b_sign2 = 4'd0; b_sign3 = 4'd6;
@(posedge clk_i);
a_mant0 = 8'd86; a_mant1 = 8'd190; a_mant2 = 8'd24; a_mant3 = 8'd89;
b_mant0 = 8'd180; b_mant1 = 8'd209; b_mant2 = 8'd102; b_mant3 = 8'd204;
a_exp0 = 10'd452; a_exp1 = 10'd278; a_exp2 = 10'd301; a_exp3 = 10'd403;
b_exp0 = 10'd461; b_exp1 = 10'd309; b_exp2 = 10'd469; b_exp3 = 10'd272;
a_sign0 = 4'd8; a_sign1 = 4'd9; a_sign2 = 4'd2; a_sign3 = 4'd5;
b_sign0 = 4'd1; b_sign1 = 4'd4; b_sign2 = 4'd6; b_sign3 = 4'd3;
@(posedge clk_i);
a_mant0 = 8'd108; a_mant1 = 8'd223; a_mant2 = 8'd199; a_mant3 = 8'd115;
b_mant0 = 8'd11; b_mant1 = 8'd168; b_mant2 = 8'd210; b_mant3 = 8'd234;
a_exp0 = 10'd65; a_exp1 = 10'd407; a_exp2 = 10'd329; a_exp3 = 10'd861;
b_exp0 = 10'd400; b_exp1 = 10'd172; b_exp2 = 10'd802; b_exp3 = 10'd306;
a_sign0 = 4'd0; a_sign1 = 4'd10; a_sign2 = 4'd12; a_sign3 = 4'd13;
b_sign0 = 4'd16; b_sign1 = 4'd14; b_sign2 = 4'd15; b_sign3 = 4'd3;
@(posedge clk_i);
a_mant0 = 8'd213; a_mant1 = 8'd173; a_mant2 = 8'd172; a_mant3 = 8'd22;
b_mant0 = 8'd209; b_mant1 = 8'd102; b_mant2 = 8'd206; b_mant3 = 8'd171;
a_exp0 = 10'd874; a_exp1 = 10'd473; a_exp2 = 10'd38; a_exp3 = 10'd711;
b_exp0 = 10'd943; b_exp1 = 10'd409; b_exp2 = 10'd142; b_exp3 = 10'd371;
a_sign0 = 4'd14; a_sign1 = 4'd3; a_sign2 = 4'd7; a_sign3 = 4'd1;
b_sign0 = 4'd10; b_sign1 = 4'd5; b_sign2 = 4'd6; b_sign3 = 4'd0;
@(posedge clk_i);
a_mant0 = 8'd163; a_mant1 = 8'd129; a_mant2 = 8'd181; a_mant3 = 8'd136;
b_mant0 = 8'd131; b_mant1 = 8'd118; b_mant2 = 8'd110; b_mant3 = 8'd230;
a_exp0 = 10'd962; a_exp1 = 10'd225; a_exp2 = 10'd354; a_exp3 = 10'd659;
b_exp0 = 10'd988; b_exp1 = 10'd497; b_exp2 = 10'd488; b_exp3 = 10'd157;
a_sign0 = 4'd4; a_sign1 = 4'd15; a_sign2 = 4'd10; a_sign3 = 4'd6;
b_sign0 = 4'd2; b_sign1 = 4'd15; b_sign2 = 4'd9; b_sign3 = 4'd14;
@(posedge clk_i);
shared_exps0 = 8'd129;
shared_exps1 = 8'd148;
a_mant0 = 8'd186; a_mant1 = 8'd228; a_mant2 = 8'd19; a_mant3 = 8'd120;
b_mant0 = 8'd56; b_mant1 = 8'd231; b_mant2 = 8'd228; b_mant3 = 8'd153;
a_exp0 = 10'd497; a_exp1 = 10'd156; a_exp2 = 10'd665; a_exp3 = 10'd608;
b_exp0 = 10'd442; b_exp1 = 10'd417; b_exp2 = 10'd235; b_exp3 = 10'd366;
a_sign0 = 4'd6; a_sign1 = 4'd0; a_sign2 = 4'd15; a_sign3 = 4'd3;
b_sign0 = 4'd9; b_sign1 = 4'd3; b_sign2 = 4'd3; b_sign3 = 4'd2;
@(posedge clk_i);
a_mant0 = 8'd53; a_mant1 = 8'd1; a_mant2 = 8'd105; a_mant3 = 8'd14;
b_mant0 = 8'd138; b_mant1 = 8'd180; b_mant2 = 8'd145; b_mant3 = 8'd125;
a_exp0 = 10'd519; a_exp1 = 10'd514; a_exp2 = 10'd537; a_exp3 = 10'd647;
b_exp0 = 10'd208; b_exp1 = 10'd165; b_exp2 = 10'd433; b_exp3 = 10'd846;
a_sign0 = 4'd7; a_sign1 = 4'd12; a_sign2 = 4'd6; a_sign3 = 4'd16;
b_sign0 = 4'd7; b_sign1 = 4'd13; b_sign2 = 4'd1; b_sign3 = 4'd9;
@(posedge clk_i);
a_mant0 = 8'd140; a_mant1 = 8'd228; a_mant2 = 8'd146; a_mant3 = 8'd31;
b_mant0 = 8'd236; b_mant1 = 8'd122; b_mant2 = 8'd128; b_mant3 = 8'd166;
a_exp0 = 10'd714; a_exp1 = 10'd405; a_exp2 = 10'd529; a_exp3 = 10'd746;
b_exp0 = 10'd807; b_exp1 = 10'd523; b_exp2 = 10'd508; b_exp3 = 10'd397;
a_sign0 = 4'd3; a_sign1 = 4'd9; a_sign2 = 4'd3; a_sign3 = 4'd10;
b_sign0 = 4'd14; b_sign1 = 4'd9; b_sign2 = 4'd9; b_sign3 = 4'd5;
@(posedge clk_i);
a_mant0 = 8'd75; a_mant1 = 8'd196; a_mant2 = 8'd77; a_mant3 = 8'd127;
b_mant0 = 8'd27; b_mant1 = 8'd51; b_mant2 = 8'd107; b_mant3 = 8'd118;
a_exp0 = 10'd998; a_exp1 = 10'd772; a_exp2 = 10'd241; a_exp3 = 10'd309;
b_exp0 = 10'd348; b_exp1 = 10'd676; b_exp2 = 10'd686; b_exp3 = 10'd391;
a_sign0 = 4'd0; a_sign1 = 4'd2; a_sign2 = 4'd10; a_sign3 = 4'd4;
b_sign0 = 4'd2; b_sign1 = 4'd5; b_sign2 = 4'd12; b_sign3 = 4'd2;
@(posedge clk_i);
a_mant0 = 8'd188; a_mant1 = 8'd252; a_mant2 = 8'd219; a_mant3 = 8'd119;
b_mant0 = 8'd214; b_mant1 = 8'd166; b_mant2 = 8'd40; b_mant3 = 8'd196;
a_exp0 = 10'd524; a_exp1 = 10'd303; a_exp2 = 10'd908; a_exp3 = 10'd15;
b_exp0 = 10'd711; b_exp1 = 10'd335; b_exp2 = 10'd692; b_exp3 = 10'd155;
a_sign0 = 4'd5; a_sign1 = 4'd13; a_sign2 = 4'd8; a_sign3 = 4'd13;
b_sign0 = 4'd6; b_sign1 = 4'd13; b_sign2 = 4'd9; b_sign3 = 4'd13;
@(posedge clk_i);
a_mant0 = 8'd196; a_mant1 = 8'd92; a_mant2 = 8'd2; a_mant3 = 8'd188;
b_mant0 = 8'd21; b_mant1 = 8'd245; b_mant2 = 8'd203; b_mant3 = 8'd35;
a_exp0 = 10'd638; a_exp1 = 10'd543; a_exp2 = 10'd754; a_exp3 = 10'd510;
b_exp0 = 10'd11; b_exp1 = 10'd171; b_exp2 = 10'd780; b_exp3 = 10'd62;
a_sign0 = 4'd12; a_sign1 = 4'd3; a_sign2 = 4'd14; a_sign3 = 4'd10;
b_sign0 = 4'd9; b_sign1 = 4'd6; b_sign2 = 4'd5; b_sign3 = 4'd7;
@(posedge clk_i);
a_mant0 = 8'd232; a_mant1 = 8'd178; a_mant2 = 8'd43; a_mant3 = 8'd228;
b_mant0 = 8'd223; b_mant1 = 8'd128; b_mant2 = 8'd143; b_mant3 = 8'd170;
a_exp0 = 10'd61; a_exp1 = 10'd728; a_exp2 = 10'd882; a_exp3 = 10'd992;
b_exp0 = 10'd299; b_exp1 = 10'd410; b_exp2 = 10'd562; b_exp3 = 10'd518;
a_sign0 = 4'd7; a_sign1 = 4'd15; a_sign2 = 4'd10; a_sign3 = 4'd1;
b_sign0 = 4'd10; b_sign1 = 4'd11; b_sign2 = 4'd2; b_sign3 = 4'd13;
@(posedge clk_i);
a_mant0 = 8'd26; a_mant1 = 8'd174; a_mant2 = 8'd171; a_mant3 = 8'd176;
b_mant0 = 8'd113; b_mant1 = 8'd34; b_mant2 = 8'd170; b_mant3 = 8'd120;
a_exp0 = 10'd313; a_exp1 = 10'd225; a_exp2 = 10'd84; a_exp3 = 10'd927;
b_exp0 = 10'd146; b_exp1 = 10'd311; b_exp2 = 10'd295; b_exp3 = 10'd947;
a_sign0 = 4'd1; a_sign1 = 4'd5; a_sign2 = 4'd4; a_sign3 = 4'd8;
b_sign0 = 4'd7; b_sign1 = 4'd9; b_sign2 = 4'd9; b_sign3 = 4'd15;
@(posedge clk_i);
shared_exps0 = 8'd117;
shared_exps1 = 8'd130;
a_mant0 = 8'd103; a_mant1 = 8'd206; a_mant2 = 8'd206; a_mant3 = 8'd178;
b_mant0 = 8'd58; b_mant1 = 8'd106; b_mant2 = 8'd71; b_mant3 = 8'd191;
a_exp0 = 10'd874; a_exp1 = 10'd273; a_exp2 = 10'd988; a_exp3 = 10'd218;
b_exp0 = 10'd295; b_exp1 = 10'd653; b_exp2 = 10'd442; b_exp3 = 10'd797;
a_sign0 = 4'd5; a_sign1 = 4'd8; a_sign2 = 4'd1; a_sign3 = 4'd10;
b_sign0 = 4'd5; b_sign1 = 4'd6; b_sign2 = 4'd11; b_sign3 = 4'd14;
@(posedge clk_i);
a_mant0 = 8'd14; a_mant1 = 8'd22; a_mant2 = 8'd150; a_mant3 = 8'd253;
b_mant0 = 8'd41; b_mant1 = 8'd145; b_mant2 = 8'd237; b_mant3 = 8'd111;
a_exp0 = 10'd235; a_exp1 = 10'd429; a_exp2 = 10'd896; a_exp3 = 10'd292;
b_exp0 = 10'd594; b_exp1 = 10'd851; b_exp2 = 10'd464; b_exp3 = 10'd621;
a_sign0 = 4'd9; a_sign1 = 4'd7; a_sign2 = 4'd15; a_sign3 = 4'd2;
b_sign0 = 4'd9; b_sign1 = 4'd8; b_sign2 = 4'd11; b_sign3 = 4'd9;
@(posedge clk_i);
a_mant0 = 8'd187; a_mant1 = 8'd140; a_mant2 = 8'd29; a_mant3 = 8'd218;
b_mant0 = 8'd0; b_mant1 = 8'd151; b_mant2 = 8'd151; b_mant3 = 8'd166;
a_exp0 = 10'd151; a_exp1 = 10'd353; a_exp2 = 10'd874; a_exp3 = 10'd71;
b_exp0 = 10'd658; b_exp1 = 10'd655; b_exp2 = 10'd802; b_exp3 = 10'd860;
a_sign0 = 4'd15; a_sign1 = 4'd16; a_sign2 = 4'd7; a_sign3 = 4'd11;
b_sign0 = 4'd2; b_sign1 = 4'd1; b_sign2 = 4'd15; b_sign3 = 4'd6;
@(posedge clk_i);
a_mant0 = 8'd138; a_mant1 = 8'd237; a_mant2 = 8'd171; a_mant3 = 8'd217;
b_mant0 = 8'd91; b_mant1 = 8'd80; b_mant2 = 8'd129; b_mant3 = 8'd154;
a_exp0 = 10'd129; a_exp1 = 10'd459; a_exp2 = 10'd633; a_exp3 = 10'd976;
b_exp0 = 10'd57; b_exp1 = 10'd55; b_exp2 = 10'd478; b_exp3 = 10'd408;
a_sign0 = 4'd6; a_sign1 = 4'd4; a_sign2 = 4'd12; a_sign3 = 4'd13;
b_sign0 = 4'd7; b_sign1 = 4'd15; b_sign2 = 4'd12; b_sign3 = 4'd15;
@(posedge clk_i);
a_mant0 = 8'd73; a_mant1 = 8'd23; a_mant2 = 8'd179; a_mant3 = 8'd31;
b_mant0 = 8'd148; b_mant1 = 8'd201; b_mant2 = 8'd156; b_mant3 = 8'd218;
a_exp0 = 10'd950; a_exp1 = 10'd59; a_exp2 = 10'd272; a_exp3 = 10'd553;
b_exp0 = 10'd886; b_exp1 = 10'd127; b_exp2 = 10'd136; b_exp3 = 10'd270;
a_sign0 = 4'd0; a_sign1 = 4'd8; a_sign2 = 4'd4; a_sign3 = 4'd5;
b_sign0 = 4'd2; b_sign1 = 4'd8; b_sign2 = 4'd9; b_sign3 = 4'd7;
@(posedge clk_i);
a_mant0 = 8'd206; a_mant1 = 8'd147; a_mant2 = 8'd105; a_mant3 = 8'd181;
b_mant0 = 8'd130; b_mant1 = 8'd39; b_mant2 = 8'd22; b_mant3 = 8'd99;
a_exp0 = 10'd102; a_exp1 = 10'd563; a_exp2 = 10'd115; a_exp3 = 10'd897;
b_exp0 = 10'd717; b_exp1 = 10'd62; b_exp2 = 10'd213; b_exp3 = 10'd614;
a_sign0 = 4'd0; a_sign1 = 4'd6; a_sign2 = 4'd5; a_sign3 = 4'd0;
b_sign0 = 4'd11; b_sign1 = 4'd9; b_sign2 = 4'd10; b_sign3 = 4'd0;
@(posedge clk_i);
a_mant0 = 8'd133; a_mant1 = 8'd174; a_mant2 = 8'd2; a_mant3 = 8'd129;
b_mant0 = 8'd18; b_mant1 = 8'd78; b_mant2 = 8'd166; b_mant3 = 8'd222;
a_exp0 = 10'd188; a_exp1 = 10'd473; a_exp2 = 10'd429; a_exp3 = 10'd930;
b_exp0 = 10'd890; b_exp1 = 10'd724; b_exp2 = 10'd468; b_exp3 = 10'd459;
a_sign0 = 4'd2; a_sign1 = 4'd9; a_sign2 = 4'd10; a_sign3 = 4'd7;
b_sign0 = 4'd0; b_sign1 = 4'd12; b_sign2 = 4'd4; b_sign3 = 4'd16;
@(posedge clk_i);
a_mant0 = 8'd154; a_mant1 = 8'd186; a_mant2 = 8'd175; a_mant3 = 8'd68;
b_mant0 = 8'd53; b_mant1 = 8'd99; b_mant2 = 8'd21; b_mant3 = 8'd150;
a_exp0 = 10'd308; a_exp1 = 10'd362; a_exp2 = 10'd975; a_exp3 = 10'd740;
b_exp0 = 10'd183; b_exp1 = 10'd333; b_exp2 = 10'd941; b_exp3 = 10'd691;
a_sign0 = 4'd9; a_sign1 = 4'd0; a_sign2 = 4'd3; a_sign3 = 4'd0;
b_sign0 = 4'd3; b_sign1 = 4'd5; b_sign2 = 4'd12; b_sign3 = 4'd3;
@(posedge clk_i);
shared_exps0 = 8'd140;
shared_exps1 = 8'd115;
a_mant0 = 8'd209; a_mant1 = 8'd23; a_mant2 = 8'd83; a_mant3 = 8'd116;
b_mant0 = 8'd224; b_mant1 = 8'd11; b_mant2 = 8'd245; b_mant3 = 8'd99;
a_exp0 = 10'd769; a_exp1 = 10'd359; a_exp2 = 10'd200; a_exp3 = 10'd486;
b_exp0 = 10'd387; b_exp1 = 10'd587; b_exp2 = 10'd723; b_exp3 = 10'd923;
a_sign0 = 4'd4; a_sign1 = 4'd9; a_sign2 = 4'd0; a_sign3 = 4'd12;
b_sign0 = 4'd15; b_sign1 = 4'd1; b_sign2 = 4'd2; b_sign3 = 4'd11;
@(posedge clk_i);
a_mant0 = 8'd13; a_mant1 = 8'd166; a_mant2 = 8'd32; a_mant3 = 8'd12;
b_mant0 = 8'd4; b_mant1 = 8'd74; b_mant2 = 8'd78; b_mant3 = 8'd214;
a_exp0 = 10'd266; a_exp1 = 10'd932; a_exp2 = 10'd975; a_exp3 = 10'd348;
b_exp0 = 10'd100; b_exp1 = 10'd661; b_exp2 = 10'd949; b_exp3 = 10'd656;
a_sign0 = 4'd16; a_sign1 = 4'd7; a_sign2 = 4'd10; a_sign3 = 4'd9;
b_sign0 = 4'd8; b_sign1 = 4'd0; b_sign2 = 4'd9; b_sign3 = 4'd5;
@(posedge clk_i);
a_mant0 = 8'd225; a_mant1 = 8'd190; a_mant2 = 8'd221; a_mant3 = 8'd204;
b_mant0 = 8'd188; b_mant1 = 8'd50; b_mant2 = 8'd150; b_mant3 = 8'd108;
a_exp0 = 10'd228; a_exp1 = 10'd985; a_exp2 = 10'd724; a_exp3 = 10'd957;
b_exp0 = 10'd763; b_exp1 = 10'd618; b_exp2 = 10'd158; b_exp3 = 10'd824;
a_sign0 = 4'd12; a_sign1 = 4'd10; a_sign2 = 4'd1; a_sign3 = 4'd3;
b_sign0 = 4'd13; b_sign1 = 4'd11; b_sign2 = 4'd3; b_sign3 = 4'd5;
@(posedge clk_i);
a_mant0 = 8'd216; a_mant1 = 8'd167; a_mant2 = 8'd137; a_mant3 = 8'd22;
b_mant0 = 8'd42; b_mant1 = 8'd147; b_mant2 = 8'd204; b_mant3 = 8'd40;
a_exp0 = 10'd1021; a_exp1 = 10'd441; a_exp2 = 10'd114; a_exp3 = 10'd861;
b_exp0 = 10'd902; b_exp1 = 10'd650; b_exp2 = 10'd165; b_exp3 = 10'd880;
a_sign0 = 4'd4; a_sign1 = 4'd10; a_sign2 = 4'd15; a_sign3 = 4'd16;
b_sign0 = 4'd11; b_sign1 = 4'd6; b_sign2 = 4'd11; b_sign3 = 4'd8;
@(posedge clk_i);
a_mant0 = 8'd134; a_mant1 = 8'd108; a_mant2 = 8'd150; a_mant3 = 8'd48;
b_mant0 = 8'd133; b_mant1 = 8'd240; b_mant2 = 8'd131; b_mant3 = 8'd84;
a_exp0 = 10'd798; a_exp1 = 10'd487; a_exp2 = 10'd748; a_exp3 = 10'd417;
b_exp0 = 10'd134; b_exp1 = 10'd84; b_exp2 = 10'd980; b_exp3 = 10'd646;
a_sign0 = 4'd2; a_sign1 = 4'd13; a_sign2 = 4'd4; a_sign3 = 4'd5;
b_sign0 = 4'd8; b_sign1 = 4'd2; b_sign2 = 4'd9; b_sign3 = 4'd5;
@(posedge clk_i);
a_mant0 = 8'd0; a_mant1 = 8'd48; a_mant2 = 8'd5; a_mant3 = 8'd138;
b_mant0 = 8'd122; b_mant1 = 8'd123; b_mant2 = 8'd33; b_mant3 = 8'd184;
a_exp0 = 10'd401; a_exp1 = 10'd606; a_exp2 = 10'd563; a_exp3 = 10'd68;
b_exp0 = 10'd890; b_exp1 = 10'd412; b_exp2 = 10'd715; b_exp3 = 10'd701;
a_sign0 = 4'd12; a_sign1 = 4'd16; a_sign2 = 4'd2; a_sign3 = 4'd5;
b_sign0 = 4'd10; b_sign1 = 4'd3; b_sign2 = 4'd12; b_sign3 = 4'd16;
@(posedge clk_i);
a_mant0 = 8'd91; a_mant1 = 8'd189; a_mant2 = 8'd213; a_mant3 = 8'd40;
b_mant0 = 8'd49; b_mant1 = 8'd19; b_mant2 = 8'd102; b_mant3 = 8'd182;
a_exp0 = 10'd904; a_exp1 = 10'd777; a_exp2 = 10'd445; a_exp3 = 10'd807;
b_exp0 = 10'd603; b_exp1 = 10'd906; b_exp2 = 10'd835; b_exp3 = 10'd906;
a_sign0 = 4'd10; a_sign1 = 4'd1; a_sign2 = 4'd16; a_sign3 = 4'd5;
b_sign0 = 4'd4; b_sign1 = 4'd10; b_sign2 = 4'd3; b_sign3 = 4'd15;
@(posedge clk_i);
a_mant0 = 8'd135; a_mant1 = 8'd23; a_mant2 = 8'd33; a_mant3 = 8'd74;
b_mant0 = 8'd175; b_mant1 = 8'd158; b_mant2 = 8'd132; b_mant3 = 8'd182;
a_exp0 = 10'd841; a_exp1 = 10'd5; a_exp2 = 10'd628; a_exp3 = 10'd820;
b_exp0 = 10'd822; b_exp1 = 10'd731; b_exp2 = 10'd621; b_exp3 = 10'd936;
a_sign0 = 4'd5; a_sign1 = 4'd16; a_sign2 = 4'd9; a_sign3 = 4'd13;
b_sign0 = 4'd6; b_sign1 = 4'd2; b_sign2 = 4'd1; b_sign3 = 4'd10;
@(posedge clk_i);
shared_exps0 = 8'd115;
shared_exps1 = 8'd122;
rstn = 0;
@(posedge clk_i);
rstn = 1;
a_mant0 = 8'd184; a_mant1 = 8'd36; a_mant2 = 8'd99; a_mant3 = 8'd81;
b_mant0 = 8'd33; b_mant1 = 8'd152; b_mant2 = 8'd210; b_mant3 = 8'd120;
a_exp0 = 10'd287; a_exp1 = 10'd273; a_exp2 = 10'd976; a_exp3 = 10'd768;
b_exp0 = 10'd142; b_exp1 = 10'd389; b_exp2 = 10'd1023; b_exp3 = 10'd876;
a_sign0 = 4'd15; a_sign1 = 4'd3; a_sign2 = 4'd12; a_sign3 = 4'd14;
b_sign0 = 4'd13; b_sign1 = 4'd13; b_sign2 = 4'd12; b_sign3 = 4'd6;
@(posedge clk_i);
a_mant0 = 8'd164; a_mant1 = 8'd241; a_mant2 = 8'd158; a_mant3 = 8'd5;
b_mant0 = 8'd82; b_mant1 = 8'd222; b_mant2 = 8'd152; b_mant3 = 8'd78;
a_exp0 = 10'd823; a_exp1 = 10'd411; a_exp2 = 10'd453; a_exp3 = 10'd848;
b_exp0 = 10'd38; b_exp1 = 10'd263; b_exp2 = 10'd302; b_exp3 = 10'd476;
a_sign0 = 4'd9; a_sign1 = 4'd4; a_sign2 = 4'd7; a_sign3 = 4'd4;
b_sign0 = 4'd9; b_sign1 = 4'd2; b_sign2 = 4'd8; b_sign3 = 4'd0;
@(posedge clk_i);
a_mant0 = 8'd180; a_mant1 = 8'd197; a_mant2 = 8'd117; a_mant3 = 8'd72;
b_mant0 = 8'd112; b_mant1 = 8'd109; b_mant2 = 8'd138; b_mant3 = 8'd52;
a_exp0 = 10'd366; a_exp1 = 10'd348; a_exp2 = 10'd331; a_exp3 = 10'd29;
b_exp0 = 10'd877; b_exp1 = 10'd355; b_exp2 = 10'd294; b_exp3 = 10'd339;
a_sign0 = 4'd6; a_sign1 = 4'd0; a_sign2 = 4'd2; a_sign3 = 4'd11;
b_sign0 = 4'd3; b_sign1 = 4'd9; b_sign2 = 4'd15; b_sign3 = 4'd7;
@(posedge clk_i);
a_mant0 = 8'd108; a_mant1 = 8'd215; a_mant2 = 8'd134; a_mant3 = 8'd70;
b_mant0 = 8'd210; b_mant1 = 8'd39; b_mant2 = 8'd178; b_mant3 = 8'd54;
a_exp0 = 10'd299; a_exp1 = 10'd498; a_exp2 = 10'd807; a_exp3 = 10'd61;
b_exp0 = 10'd291; b_exp1 = 10'd415; b_exp2 = 10'd464; b_exp3 = 10'd727;
a_sign0 = 4'd2; a_sign1 = 4'd6; a_sign2 = 4'd3; a_sign3 = 4'd0;
b_sign0 = 4'd6; b_sign1 = 4'd5; b_sign2 = 4'd15; b_sign3 = 4'd15;
@(posedge clk_i);
a_mant0 = 8'd90; a_mant1 = 8'd135; a_mant2 = 8'd149; a_mant3 = 8'd62;
b_mant0 = 8'd107; b_mant1 = 8'd199; b_mant2 = 8'd182; b_mant3 = 8'd238;
a_exp0 = 10'd810; a_exp1 = 10'd51; a_exp2 = 10'd724; a_exp3 = 10'd938;
b_exp0 = 10'd78; b_exp1 = 10'd18; b_exp2 = 10'd743; b_exp3 = 10'd840;
a_sign0 = 4'd3; a_sign1 = 4'd2; a_sign2 = 4'd10; a_sign3 = 4'd15;
b_sign0 = 4'd16; b_sign1 = 4'd6; b_sign2 = 4'd2; b_sign3 = 4'd4;
@(posedge clk_i);
a_mant0 = 8'd223; a_mant1 = 8'd47; a_mant2 = 8'd165; a_mant3 = 8'd200;
b_mant0 = 8'd53; b_mant1 = 8'd4; b_mant2 = 8'd62; b_mant3 = 8'd7;
a_exp0 = 10'd767; a_exp1 = 10'd597; a_exp2 = 10'd193; a_exp3 = 10'd429;
b_exp0 = 10'd207; b_exp1 = 10'd671; b_exp2 = 10'd382; b_exp3 = 10'd895;
a_sign0 = 4'd15; a_sign1 = 4'd0; a_sign2 = 4'd0; a_sign3 = 4'd5;
b_sign0 = 4'd6; b_sign1 = 4'd16; b_sign2 = 4'd2; b_sign3 = 4'd9;
@(posedge clk_i);
a_mant0 = 8'd211; a_mant1 = 8'd34; a_mant2 = 8'd1; a_mant3 = 8'd40;
b_mant0 = 8'd222; b_mant1 = 8'd240; b_mant2 = 8'd190; b_mant3 = 8'd156;
a_exp0 = 10'd602; a_exp1 = 10'd39; a_exp2 = 10'd694; a_exp3 = 10'd944;
b_exp0 = 10'd66; b_exp1 = 10'd964; b_exp2 = 10'd181; b_exp3 = 10'd349;
a_sign0 = 4'd2; a_sign1 = 4'd4; a_sign2 = 4'd10; a_sign3 = 4'd0;
b_sign0 = 4'd7; b_sign1 = 4'd15; b_sign2 = 4'd6; b_sign3 = 4'd0;
@(posedge clk_i);
shared_exps0 = 8'd113;
shared_exps1 = 8'd136;
a_mant0 = 8'd29; a_mant1 = 8'd198; a_mant2 = 8'd212; a_mant3 = 8'd185;
b_mant0 = 8'd97; b_mant1 = 8'd198; b_mant2 = 8'd126; b_mant3 = 8'd59;
a_exp0 = 10'd710; a_exp1 = 10'd1003; a_exp2 = 10'd832; a_exp3 = 10'd696;
b_exp0 = 10'd94; b_exp1 = 10'd345; b_exp2 = 10'd888; b_exp3 = 10'd335;
a_sign0 = 4'd1; a_sign1 = 4'd6; a_sign2 = 4'd10; a_sign3 = 4'd15;
b_sign0 = 4'd3; b_sign1 = 4'd13; b_sign2 = 4'd11; b_sign3 = 4'd3;
@(posedge clk_i);
a_mant0 = 8'd134; a_mant1 = 8'd60; a_mant2 = 8'd141; a_mant3 = 8'd22;
b_mant0 = 8'd201; b_mant1 = 8'd200; b_mant2 = 8'd206; b_mant3 = 8'd112;
a_exp0 = 10'd998; a_exp1 = 10'd195; a_exp2 = 10'd560; a_exp3 = 10'd678;
b_exp0 = 10'd101; b_exp1 = 10'd461; b_exp2 = 10'd560; b_exp3 = 10'd1000;
a_sign0 = 4'd5; a_sign1 = 4'd7; a_sign2 = 4'd7; a_sign3 = 4'd0;
b_sign0 = 4'd10; b_sign1 = 4'd16; b_sign2 = 4'd14; b_sign3 = 4'd2;
@(posedge clk_i);
a_mant0 = 8'd228; a_mant1 = 8'd200; a_mant2 = 8'd81; a_mant3 = 8'd70;
b_mant0 = 8'd115; b_mant1 = 8'd235; b_mant2 = 8'd222; b_mant3 = 8'd53;
a_exp0 = 10'd197; a_exp1 = 10'd786; a_exp2 = 10'd863; a_exp3 = 10'd795;
b_exp0 = 10'd769; b_exp1 = 10'd911; b_exp2 = 10'd983; b_exp3 = 10'd46;
a_sign0 = 4'd6; a_sign1 = 4'd10; a_sign2 = 4'd16; a_sign3 = 4'd10;
b_sign0 = 4'd4; b_sign1 = 4'd12; b_sign2 = 4'd3; b_sign3 = 4'd7;
@(posedge clk_i);
a_mant0 = 8'd125; a_mant1 = 8'd1; a_mant2 = 8'd207; a_mant3 = 8'd249;
b_mant0 = 8'd248; b_mant1 = 8'd218; b_mant2 = 8'd82; b_mant3 = 8'd95;
a_exp0 = 10'd593; a_exp1 = 10'd265; a_exp2 = 10'd38; a_exp3 = 10'd669;
b_exp0 = 10'd775; b_exp1 = 10'd219; b_exp2 = 10'd350; b_exp3 = 10'd456;
a_sign0 = 4'd16; a_sign1 = 4'd11; a_sign2 = 4'd14; a_sign3 = 4'd7;
b_sign0 = 4'd12; b_sign1 = 4'd10; b_sign2 = 4'd5; b_sign3 = 4'd16;
@(posedge clk_i);
a_mant0 = 8'd159; a_mant1 = 8'd6; a_mant2 = 8'd244; a_mant3 = 8'd220;
b_mant0 = 8'd3; b_mant1 = 8'd129; b_mant2 = 8'd1; b_mant3 = 8'd21;
a_exp0 = 10'd864; a_exp1 = 10'd999; a_exp2 = 10'd376; a_exp3 = 10'd491;
b_exp0 = 10'd697; b_exp1 = 10'd766; b_exp2 = 10'd872; b_exp3 = 10'd810;
a_sign0 = 4'd2; a_sign1 = 4'd9; a_sign2 = 4'd11; a_sign3 = 4'd16;
b_sign0 = 4'd1; b_sign1 = 4'd16; b_sign2 = 4'd11; b_sign3 = 4'd9;
@(posedge clk_i);
a_mant0 = 8'd73; a_mant1 = 8'd187; a_mant2 = 8'd224; a_mant3 = 8'd119;
b_mant0 = 8'd139; b_mant1 = 8'd188; b_mant2 = 8'd120; b_mant3 = 8'd127;
a_exp0 = 10'd516; a_exp1 = 10'd420; a_exp2 = 10'd968; a_exp3 = 10'd905;
b_exp0 = 10'd764; b_exp1 = 10'd787; b_exp2 = 10'd499; b_exp3 = 10'd780;
a_sign0 = 4'd16; a_sign1 = 4'd5; a_sign2 = 4'd6; a_sign3 = 4'd9;
b_sign0 = 4'd15; b_sign1 = 4'd6; b_sign2 = 4'd14; b_sign3 = 4'd14;
@(posedge clk_i);
a_mant0 = 8'd92; a_mant1 = 8'd14; a_mant2 = 8'd67; a_mant3 = 8'd248;
b_mant0 = 8'd204; b_mant1 = 8'd161; b_mant2 = 8'd63; b_mant3 = 8'd35;
a_exp0 = 10'd526; a_exp1 = 10'd603; a_exp2 = 10'd9; a_exp3 = 10'd367;
b_exp0 = 10'd735; b_exp1 = 10'd932; b_exp2 = 10'd351; b_exp3 = 10'd360;
a_sign0 = 4'd0; a_sign1 = 4'd0; a_sign2 = 4'd12; a_sign3 = 4'd11;
b_sign0 = 4'd0; b_sign1 = 4'd8; b_sign2 = 4'd8; b_sign3 = 4'd1;
@(posedge clk_i);
a_mant0 = 8'd33; a_mant1 = 8'd155; a_mant2 = 8'd55; a_mant3 = 8'd239;
b_mant0 = 8'd239; b_mant1 = 8'd156; b_mant2 = 8'd98; b_mant3 = 8'd105;
a_exp0 = 10'd156; a_exp1 = 10'd966; a_exp2 = 10'd354; a_exp3 = 10'd571;
b_exp0 = 10'd183; b_exp1 = 10'd913; b_exp2 = 10'd925; b_exp3 = 10'd412;
a_sign0 = 4'd9; a_sign1 = 4'd1; a_sign2 = 4'd10; a_sign3 = 4'd7;
b_sign0 = 4'd12; b_sign1 = 4'd10; b_sign2 = 4'd4; b_sign3 = 4'd9;
@(posedge clk_i);
shared_exps0 = 8'd124;
shared_exps1 = 8'd128;
a_mant0 = 8'd123; a_mant1 = 8'd109; a_mant2 = 8'd130; a_mant3 = 8'd228;
b_mant0 = 8'd46; b_mant1 = 8'd232; b_mant2 = 8'd178; b_mant3 = 8'd161;
a_exp0 = 10'd516; a_exp1 = 10'd547; a_exp2 = 10'd34; a_exp3 = 10'd816;
b_exp0 = 10'd536; b_exp1 = 10'd162; b_exp2 = 10'd373; b_exp3 = 10'd821;
a_sign0 = 4'd14; a_sign1 = 4'd15; a_sign2 = 4'd4; a_sign3 = 4'd13;
b_sign0 = 4'd6; b_sign1 = 4'd13; b_sign2 = 4'd13; b_sign3 = 4'd8;
@(posedge clk_i);
a_mant0 = 8'd87; a_mant1 = 8'd15; a_mant2 = 8'd52; a_mant3 = 8'd218;
b_mant0 = 8'd90; b_mant1 = 8'd157; b_mant2 = 8'd44; b_mant3 = 8'd157;
a_exp0 = 10'd320; a_exp1 = 10'd136; a_exp2 = 10'd968; a_exp3 = 10'd835;
b_exp0 = 10'd33; b_exp1 = 10'd168; b_exp2 = 10'd135; b_exp3 = 10'd295;
a_sign0 = 4'd0; a_sign1 = 4'd2; a_sign2 = 4'd6; a_sign3 = 4'd4;
b_sign0 = 4'd2; b_sign1 = 4'd12; b_sign2 = 4'd3; b_sign3 = 4'd15;
@(posedge clk_i);
a_mant0 = 8'd163; a_mant1 = 8'd4; a_mant2 = 8'd168; a_mant3 = 8'd172;
b_mant0 = 8'd244; b_mant1 = 8'd145; b_mant2 = 8'd88; b_mant3 = 8'd41;
a_exp0 = 10'd1000; a_exp1 = 10'd462; a_exp2 = 10'd727; a_exp3 = 10'd1008;
b_exp0 = 10'd497; b_exp1 = 10'd922; b_exp2 = 10'd222; b_exp3 = 10'd19;
a_sign0 = 4'd10; a_sign1 = 4'd2; a_sign2 = 4'd10; a_sign3 = 4'd4;
b_sign0 = 4'd0; b_sign1 = 4'd11; b_sign2 = 4'd14; b_sign3 = 4'd7;
@(posedge clk_i);
a_mant0 = 8'd141; a_mant1 = 8'd96; a_mant2 = 8'd57; a_mant3 = 8'd226;
b_mant0 = 8'd175; b_mant1 = 8'd37; b_mant2 = 8'd247; b_mant3 = 8'd73;
a_exp0 = 10'd55; a_exp1 = 10'd61; a_exp2 = 10'd860; a_exp3 = 10'd574;
b_exp0 = 10'd866; b_exp1 = 10'd192; b_exp2 = 10'd841; b_exp3 = 10'd872;
a_sign0 = 4'd15; a_sign1 = 4'd3; a_sign2 = 4'd11; a_sign3 = 4'd2;
b_sign0 = 4'd0; b_sign1 = 4'd11; b_sign2 = 4'd14; b_sign3 = 4'd1;
@(posedge clk_i);
a_mant0 = 8'd243; a_mant1 = 8'd133; a_mant2 = 8'd149; a_mant3 = 8'd251;
b_mant0 = 8'd61; b_mant1 = 8'd90; b_mant2 = 8'd67; b_mant3 = 8'd139;
a_exp0 = 10'd308; a_exp1 = 10'd804; a_exp2 = 10'd39; a_exp3 = 10'd306;
b_exp0 = 10'd982; b_exp1 = 10'd500; b_exp2 = 10'd816; b_exp3 = 10'd793;
a_sign0 = 4'd14; a_sign1 = 4'd12; a_sign2 = 4'd5; a_sign3 = 4'd8;
b_sign0 = 4'd16; b_sign1 = 4'd2; b_sign2 = 4'd15; b_sign3 = 4'd12;
@(posedge clk_i);
a_mant0 = 8'd70; a_mant1 = 8'd66; a_mant2 = 8'd119; a_mant3 = 8'd79;
b_mant0 = 8'd190; b_mant1 = 8'd128; b_mant2 = 8'd225; b_mant3 = 8'd167;
a_exp0 = 10'd660; a_exp1 = 10'd239; a_exp2 = 10'd515; a_exp3 = 10'd239;
b_exp0 = 10'd313; b_exp1 = 10'd716; b_exp2 = 10'd711; b_exp3 = 10'd683;
a_sign0 = 4'd7; a_sign1 = 4'd10; a_sign2 = 4'd10; a_sign3 = 4'd2;
b_sign0 = 4'd5; b_sign1 = 4'd14; b_sign2 = 4'd10; b_sign3 = 4'd1;
@(posedge clk_i);
a_mant0 = 8'd202; a_mant1 = 8'd204; a_mant2 = 8'd165; a_mant3 = 8'd25;
b_mant0 = 8'd223; b_mant1 = 8'd45; b_mant2 = 8'd130; b_mant3 = 8'd47;
a_exp0 = 10'd1023; a_exp1 = 10'd90; a_exp2 = 10'd63; a_exp3 = 10'd80;
b_exp0 = 10'd922; b_exp1 = 10'd132; b_exp2 = 10'd214; b_exp3 = 10'd1;
a_sign0 = 4'd13; a_sign1 = 4'd4; a_sign2 = 4'd7; a_sign3 = 4'd4;
b_sign0 = 4'd5; b_sign1 = 4'd13; b_sign2 = 4'd10; b_sign3 = 4'd4;
@(posedge clk_i);
a_mant0 = 8'd8; a_mant1 = 8'd216; a_mant2 = 8'd18; a_mant3 = 8'd233;
b_mant0 = 8'd180; b_mant1 = 8'd24; b_mant2 = 8'd171; b_mant3 = 8'd200;
a_exp0 = 10'd175; a_exp1 = 10'd433; a_exp2 = 10'd538; a_exp3 = 10'd645;
b_exp0 = 10'd160; b_exp1 = 10'd539; b_exp2 = 10'd778; b_exp3 = 10'd556;
a_sign0 = 4'd7; a_sign1 = 4'd10; a_sign2 = 4'd7; a_sign3 = 4'd4;
b_sign0 = 4'd16; b_sign1 = 4'd13; b_sign2 = 4'd2; b_sign3 = 4'd4;
@(posedge clk_i);
shared_exps0 = 8'd116;
shared_exps1 = 8'd140;
a_mant0 = 8'd116; a_mant1 = 8'd214; a_mant2 = 8'd59; a_mant3 = 8'd18;
b_mant0 = 8'd177; b_mant1 = 8'd103; b_mant2 = 8'd72; b_mant3 = 8'd223;
a_exp0 = 10'd152; a_exp1 = 10'd234; a_exp2 = 10'd0; a_exp3 = 10'd866;
b_exp0 = 10'd146; b_exp1 = 10'd104; b_exp2 = 10'd129; b_exp3 = 10'd940;
a_sign0 = 4'd13; a_sign1 = 4'd9; a_sign2 = 4'd0; a_sign3 = 4'd14;
b_sign0 = 4'd3; b_sign1 = 4'd7; b_sign2 = 4'd6; b_sign3 = 4'd3;
@(posedge clk_i);
a_mant0 = 8'd138; a_mant1 = 8'd87; a_mant2 = 8'd205; a_mant3 = 8'd35;
b_mant0 = 8'd96; b_mant1 = 8'd18; b_mant2 = 8'd60; b_mant3 = 8'd9;
a_exp0 = 10'd665; a_exp1 = 10'd360; a_exp2 = 10'd999; a_exp3 = 10'd519;
b_exp0 = 10'd955; b_exp1 = 10'd850; b_exp2 = 10'd26; b_exp3 = 10'd1015;
a_sign0 = 4'd9; a_sign1 = 4'd3; a_sign2 = 4'd3; a_sign3 = 4'd6;
b_sign0 = 4'd13; b_sign1 = 4'd8; b_sign2 = 4'd6; b_sign3 = 4'd16;
@(posedge clk_i);
a_mant0 = 8'd61; a_mant1 = 8'd244; a_mant2 = 8'd58; a_mant3 = 8'd74;
b_mant0 = 8'd31; b_mant1 = 8'd98; b_mant2 = 8'd191; b_mant3 = 8'd142;
a_exp0 = 10'd987; a_exp1 = 10'd659; a_exp2 = 10'd1019; a_exp3 = 10'd363;
b_exp0 = 10'd816; b_exp1 = 10'd958; b_exp2 = 10'd845; b_exp3 = 10'd584;
a_sign0 = 4'd0; a_sign1 = 4'd4; a_sign2 = 4'd16; a_sign3 = 4'd0;
b_sign0 = 4'd15; b_sign1 = 4'd11; b_sign2 = 4'd3; b_sign3 = 4'd15;
@(posedge clk_i);
a_mant0 = 8'd121; a_mant1 = 8'd181; a_mant2 = 8'd184; a_mant3 = 8'd227;
b_mant0 = 8'd160; b_mant1 = 8'd94; b_mant2 = 8'd220; b_mant3 = 8'd103;
a_exp0 = 10'd980; a_exp1 = 10'd16; a_exp2 = 10'd845; a_exp3 = 10'd770;
b_exp0 = 10'd185; b_exp1 = 10'd527; b_exp2 = 10'd494; b_exp3 = 10'd194;
a_sign0 = 4'd5; a_sign1 = 4'd0; a_sign2 = 4'd13; a_sign3 = 4'd1;
b_sign0 = 4'd16; b_sign1 = 4'd10; b_sign2 = 4'd7; b_sign3 = 4'd4;
@(posedge clk_i);
a_mant0 = 8'd198; a_mant1 = 8'd218; a_mant2 = 8'd41; a_mant3 = 8'd135;
b_mant0 = 8'd14; b_mant1 = 8'd81; b_mant2 = 8'd113; b_mant3 = 8'd208;
a_exp0 = 10'd1; a_exp1 = 10'd547; a_exp2 = 10'd211; a_exp3 = 10'd898;
b_exp0 = 10'd883; b_exp1 = 10'd429; b_exp2 = 10'd939; b_exp3 = 10'd153;
a_sign0 = 4'd7; a_sign1 = 4'd9; a_sign2 = 4'd7; a_sign3 = 4'd7;
b_sign0 = 4'd16; b_sign1 = 4'd15; b_sign2 = 4'd3; b_sign3 = 4'd8;
@(posedge clk_i);
a_mant0 = 8'd207; a_mant1 = 8'd20; a_mant2 = 8'd249; a_mant3 = 8'd214;
b_mant0 = 8'd123; b_mant1 = 8'd133; b_mant2 = 8'd250; b_mant3 = 8'd243;
a_exp0 = 10'd186; a_exp1 = 10'd185; a_exp2 = 10'd457; a_exp3 = 10'd660;
b_exp0 = 10'd943; b_exp1 = 10'd470; b_exp2 = 10'd254; b_exp3 = 10'd531;
a_sign0 = 4'd7; a_sign1 = 4'd6; a_sign2 = 4'd9; a_sign3 = 4'd5;
b_sign0 = 4'd3; b_sign1 = 4'd13; b_sign2 = 4'd1; b_sign3 = 4'd5;
@(posedge clk_i);
a_mant0 = 8'd222; a_mant1 = 8'd57; a_mant2 = 8'd45; a_mant3 = 8'd139;
b_mant0 = 8'd14; b_mant1 = 8'd105; b_mant2 = 8'd255; b_mant3 = 8'd166;
a_exp0 = 10'd9; a_exp1 = 10'd555; a_exp2 = 10'd347; a_exp3 = 10'd867;
b_exp0 = 10'd494; b_exp1 = 10'd283; b_exp2 = 10'd768; b_exp3 = 10'd800;
a_sign0 = 4'd4; a_sign1 = 4'd0; a_sign2 = 4'd8; a_sign3 = 4'd14;
b_sign0 = 4'd1; b_sign1 = 4'd14; b_sign2 = 4'd12; b_sign3 = 4'd11;
@(posedge clk_i);
a_mant0 = 8'd85; a_mant1 = 8'd213; a_mant2 = 8'd131; a_mant3 = 8'd233;
b_mant0 = 8'd24; b_mant1 = 8'd1; b_mant2 = 8'd66; b_mant3 = 8'd75;
a_exp0 = 10'd775; a_exp1 = 10'd175; a_exp2 = 10'd697; a_exp3 = 10'd605;
b_exp0 = 10'd454; b_exp1 = 10'd878; b_exp2 = 10'd721; b_exp3 = 10'd274;
a_sign0 = 4'd13; a_sign1 = 4'd9; a_sign2 = 4'd4; a_sign3 = 4'd1;
b_sign0 = 4'd13; b_sign1 = 4'd2; b_sign2 = 4'd2; b_sign3 = 4'd2;
@(posedge clk_i);
shared_exps0 = 8'd145;
shared_exps1 = 8'd123;
rstn = 0;
@(posedge clk_i);
rstn = 1;
a_mant0 = 8'd86; a_mant1 = 8'd233; a_mant2 = 8'd153; a_mant3 = 8'd253;
b_mant0 = 8'd80; b_mant1 = 8'd8; b_mant2 = 8'd44; b_mant3 = 8'd89;
a_exp0 = 10'd415; a_exp1 = 10'd162; a_exp2 = 10'd282; a_exp3 = 10'd671;
b_exp0 = 10'd852; b_exp1 = 10'd886; b_exp2 = 10'd14; b_exp3 = 10'd780;
a_sign0 = 4'd11; a_sign1 = 4'd13; a_sign2 = 4'd3; a_sign3 = 4'd2;
b_sign0 = 4'd2; b_sign1 = 4'd11; b_sign2 = 4'd14; b_sign3 = 4'd3;
@(posedge clk_i);
a_mant0 = 8'd172; a_mant1 = 8'd140; a_mant2 = 8'd113; a_mant3 = 8'd43;
b_mant0 = 8'd37; b_mant1 = 8'd36; b_mant2 = 8'd219; b_mant3 = 8'd144;
a_exp0 = 10'd644; a_exp1 = 10'd117; a_exp2 = 10'd476; a_exp3 = 10'd713;
b_exp0 = 10'd115; b_exp1 = 10'd682; b_exp2 = 10'd441; b_exp3 = 10'd568;
a_sign0 = 4'd12; a_sign1 = 4'd6; a_sign2 = 4'd11; a_sign3 = 4'd1;
b_sign0 = 4'd14; b_sign1 = 4'd6; b_sign2 = 4'd8; b_sign3 = 4'd13;
@(posedge clk_i);
a_mant0 = 8'd28; a_mant1 = 8'd33; a_mant2 = 8'd88; a_mant3 = 8'd79;
b_mant0 = 8'd230; b_mant1 = 8'd222; b_mant2 = 8'd62; b_mant3 = 8'd7;
a_exp0 = 10'd582; a_exp1 = 10'd337; a_exp2 = 10'd667; a_exp3 = 10'd159;
b_exp0 = 10'd638; b_exp1 = 10'd94; b_exp2 = 10'd727; b_exp3 = 10'd546;
a_sign0 = 4'd4; a_sign1 = 4'd11; a_sign2 = 4'd1; a_sign3 = 4'd4;
b_sign0 = 4'd11; b_sign1 = 4'd13; b_sign2 = 4'd15; b_sign3 = 4'd8;
@(posedge clk_i);
a_mant0 = 8'd64; a_mant1 = 8'd202; a_mant2 = 8'd111; a_mant3 = 8'd79;
b_mant0 = 8'd232; b_mant1 = 8'd62; b_mant2 = 8'd175; b_mant3 = 8'd38;
a_exp0 = 10'd558; a_exp1 = 10'd417; a_exp2 = 10'd105; a_exp3 = 10'd633;
b_exp0 = 10'd884; b_exp1 = 10'd643; b_exp2 = 10'd263; b_exp3 = 10'd548;
a_sign0 = 4'd13; a_sign1 = 4'd3; a_sign2 = 4'd0; a_sign3 = 4'd5;
b_sign0 = 4'd3; b_sign1 = 4'd12; b_sign2 = 4'd3; b_sign3 = 4'd15;
@(posedge clk_i);
a_mant0 = 8'd130; a_mant1 = 8'd148; a_mant2 = 8'd126; a_mant3 = 8'd103;
b_mant0 = 8'd28; b_mant1 = 8'd42; b_mant2 = 8'd72; b_mant3 = 8'd132;
a_exp0 = 10'd710; a_exp1 = 10'd665; a_exp2 = 10'd38; a_exp3 = 10'd52;
b_exp0 = 10'd183; b_exp1 = 10'd980; b_exp2 = 10'd34; b_exp3 = 10'd958;
a_sign0 = 4'd16; a_sign1 = 4'd0; a_sign2 = 4'd6; a_sign3 = 4'd2;
b_sign0 = 4'd1; b_sign1 = 4'd13; b_sign2 = 4'd0; b_sign3 = 4'd15;
@(posedge clk_i);
a_mant0 = 8'd57; a_mant1 = 8'd21; a_mant2 = 8'd184; a_mant3 = 8'd100;
b_mant0 = 8'd140; b_mant1 = 8'd53; b_mant2 = 8'd20; b_mant3 = 8'd163;
a_exp0 = 10'd935; a_exp1 = 10'd64; a_exp2 = 10'd330; a_exp3 = 10'd486;
b_exp0 = 10'd507; b_exp1 = 10'd978; b_exp2 = 10'd163; b_exp3 = 10'd447;
a_sign0 = 4'd12; a_sign1 = 4'd9; a_sign2 = 4'd5; a_sign3 = 4'd2;
b_sign0 = 4'd10; b_sign1 = 4'd15; b_sign2 = 4'd15; b_sign3 = 4'd13;
@(posedge clk_i);
a_mant0 = 8'd58; a_mant1 = 8'd24; a_mant2 = 8'd156; a_mant3 = 8'd20;
b_mant0 = 8'd247; b_mant1 = 8'd179; b_mant2 = 8'd240; b_mant3 = 8'd247;
a_exp0 = 10'd860; a_exp1 = 10'd48; a_exp2 = 10'd156; a_exp3 = 10'd141;
b_exp0 = 10'd671; b_exp1 = 10'd61; b_exp2 = 10'd793; b_exp3 = 10'd843;
a_sign0 = 4'd16; a_sign1 = 4'd10; a_sign2 = 4'd16; a_sign3 = 4'd3;
b_sign0 = 4'd3; b_sign1 = 4'd15; b_sign2 = 4'd4; b_sign3 = 4'd15;
@(posedge clk_i);
shared_exps0 = 8'd155;
shared_exps1 = 8'd128;
a_mant0 = 8'd131; a_mant1 = 8'd174; a_mant2 = 8'd21; a_mant3 = 8'd3;
b_mant0 = 8'd250; b_mant1 = 8'd116; b_mant2 = 8'd179; b_mant3 = 8'd38;
a_exp0 = 10'd875; a_exp1 = 10'd820; a_exp2 = 10'd190; a_exp3 = 10'd97;
b_exp0 = 10'd451; b_exp1 = 10'd389; b_exp2 = 10'd693; b_exp3 = 10'd988;
a_sign0 = 4'd10; a_sign1 = 4'd0; a_sign2 = 4'd5; a_sign3 = 4'd0;
b_sign0 = 4'd10; b_sign1 = 4'd2; b_sign2 = 4'd7; b_sign3 = 4'd3;
@(posedge clk_i);
a_mant0 = 8'd113; a_mant1 = 8'd218; a_mant2 = 8'd42; a_mant3 = 8'd1;
b_mant0 = 8'd185; b_mant1 = 8'd135; b_mant2 = 8'd131; b_mant3 = 8'd158;
a_exp0 = 10'd546; a_exp1 = 10'd564; a_exp2 = 10'd565; a_exp3 = 10'd329;
b_exp0 = 10'd948; b_exp1 = 10'd227; b_exp2 = 10'd574; b_exp3 = 10'd302;
a_sign0 = 4'd14; a_sign1 = 4'd4; a_sign2 = 4'd5; a_sign3 = 4'd5;
b_sign0 = 4'd7; b_sign1 = 4'd6; b_sign2 = 4'd5; b_sign3 = 4'd7;
@(posedge clk_i);
a_mant0 = 8'd51; a_mant1 = 8'd104; a_mant2 = 8'd19; a_mant3 = 8'd42;
b_mant0 = 8'd15; b_mant1 = 8'd68; b_mant2 = 8'd176; b_mant3 = 8'd181;
a_exp0 = 10'd909; a_exp1 = 10'd564; a_exp2 = 10'd385; a_exp3 = 10'd690;
b_exp0 = 10'd483; b_exp1 = 10'd182; b_exp2 = 10'd651; b_exp3 = 10'd572;
a_sign0 = 4'd1; a_sign1 = 4'd10; a_sign2 = 4'd16; a_sign3 = 4'd3;
b_sign0 = 4'd0; b_sign1 = 4'd8; b_sign2 = 4'd5; b_sign3 = 4'd3;
@(posedge clk_i);
a_mant0 = 8'd217; a_mant1 = 8'd215; a_mant2 = 8'd122; a_mant3 = 8'd96;
b_mant0 = 8'd210; b_mant1 = 8'd5; b_mant2 = 8'd62; b_mant3 = 8'd219;
a_exp0 = 10'd730; a_exp1 = 10'd767; a_exp2 = 10'd1003; a_exp3 = 10'd79;
b_exp0 = 10'd872; b_exp1 = 10'd169; b_exp2 = 10'd155; b_exp3 = 10'd4;
a_sign0 = 4'd6; a_sign1 = 4'd2; a_sign2 = 4'd11; a_sign3 = 4'd5;
b_sign0 = 4'd0; b_sign1 = 4'd12; b_sign2 = 4'd2; b_sign3 = 4'd14;
@(posedge clk_i);
a_mant0 = 8'd40; a_mant1 = 8'd34; a_mant2 = 8'd182; a_mant3 = 8'd143;
b_mant0 = 8'd75; b_mant1 = 8'd100; b_mant2 = 8'd103; b_mant3 = 8'd57;
a_exp0 = 10'd816; a_exp1 = 10'd626; a_exp2 = 10'd799; a_exp3 = 10'd110;
b_exp0 = 10'd909; b_exp1 = 10'd686; b_exp2 = 10'd739; b_exp3 = 10'd165;
a_sign0 = 4'd5; a_sign1 = 4'd9; a_sign2 = 4'd8; a_sign3 = 4'd1;
b_sign0 = 4'd13; b_sign1 = 4'd10; b_sign2 = 4'd2; b_sign3 = 4'd16;
@(posedge clk_i);
a_mant0 = 8'd52; a_mant1 = 8'd176; a_mant2 = 8'd31; a_mant3 = 8'd33;
b_mant0 = 8'd40; b_mant1 = 8'd14; b_mant2 = 8'd185; b_mant3 = 8'd130;
a_exp0 = 10'd823; a_exp1 = 10'd270; a_exp2 = 10'd643; a_exp3 = 10'd590;
b_exp0 = 10'd634; b_exp1 = 10'd41; b_exp2 = 10'd582; b_exp3 = 10'd704;
a_sign0 = 4'd7; a_sign1 = 4'd7; a_sign2 = 4'd11; a_sign3 = 4'd12;
b_sign0 = 4'd4; b_sign1 = 4'd6; b_sign2 = 4'd2; b_sign3 = 4'd15;
@(posedge clk_i);
a_mant0 = 8'd41; a_mant1 = 8'd50; a_mant2 = 8'd236; a_mant3 = 8'd45;
b_mant0 = 8'd103; b_mant1 = 8'd3; b_mant2 = 8'd24; b_mant3 = 8'd51;
a_exp0 = 10'd315; a_exp1 = 10'd594; a_exp2 = 10'd55; a_exp3 = 10'd177;
b_exp0 = 10'd602; b_exp1 = 10'd1007; b_exp2 = 10'd212; b_exp3 = 10'd670;
a_sign0 = 4'd3; a_sign1 = 4'd0; a_sign2 = 4'd5; a_sign3 = 4'd11;
b_sign0 = 4'd14; b_sign1 = 4'd8; b_sign2 = 4'd6; b_sign3 = 4'd7;
@(posedge clk_i);
a_mant0 = 8'd236; a_mant1 = 8'd242; a_mant2 = 8'd232; a_mant3 = 8'd2;
b_mant0 = 8'd210; b_mant1 = 8'd233; b_mant2 = 8'd221; b_mant3 = 8'd76;
a_exp0 = 10'd9; a_exp1 = 10'd789; a_exp2 = 10'd249; a_exp3 = 10'd833;
b_exp0 = 10'd715; b_exp1 = 10'd44; b_exp2 = 10'd719; b_exp3 = 10'd495;
a_sign0 = 4'd13; a_sign1 = 4'd6; a_sign2 = 4'd2; a_sign3 = 4'd10;
b_sign0 = 4'd8; b_sign1 = 4'd3; b_sign2 = 4'd9; b_sign3 = 4'd1;
@(posedge clk_i);
shared_exps0 = 8'd117;
shared_exps1 = 8'd106;
a_mant0 = 8'd57; a_mant1 = 8'd82; a_mant2 = 8'd30; a_mant3 = 8'd76;
b_mant0 = 8'd57; b_mant1 = 8'd103; b_mant2 = 8'd7; b_mant3 = 8'd106;
a_exp0 = 10'd451; a_exp1 = 10'd252; a_exp2 = 10'd588; a_exp3 = 10'd931;
b_exp0 = 10'd1001; b_exp1 = 10'd28; b_exp2 = 10'd983; b_exp3 = 10'd675;
a_sign0 = 4'd15; a_sign1 = 4'd5; a_sign2 = 4'd7; a_sign3 = 4'd0;
b_sign0 = 4'd3; b_sign1 = 4'd4; b_sign2 = 4'd0; b_sign3 = 4'd12;
@(posedge clk_i);
a_mant0 = 8'd73; a_mant1 = 8'd67; a_mant2 = 8'd21; a_mant3 = 8'd24;
b_mant0 = 8'd123; b_mant1 = 8'd56; b_mant2 = 8'd151; b_mant3 = 8'd243;
a_exp0 = 10'd702; a_exp1 = 10'd67; a_exp2 = 10'd863; a_exp3 = 10'd564;
b_exp0 = 10'd435; b_exp1 = 10'd127; b_exp2 = 10'd507; b_exp3 = 10'd425;
a_sign0 = 4'd2; a_sign1 = 4'd6; a_sign2 = 4'd11; a_sign3 = 4'd15;
b_sign0 = 4'd14; b_sign1 = 4'd0; b_sign2 = 4'd8; b_sign3 = 4'd10;
@(posedge clk_i);
a_mant0 = 8'd249; a_mant1 = 8'd71; a_mant2 = 8'd202; a_mant3 = 8'd86;
b_mant0 = 8'd98; b_mant1 = 8'd224; b_mant2 = 8'd101; b_mant3 = 8'd58;
a_exp0 = 10'd849; a_exp1 = 10'd509; a_exp2 = 10'd958; a_exp3 = 10'd394;
b_exp0 = 10'd571; b_exp1 = 10'd823; b_exp2 = 10'd516; b_exp3 = 10'd553;
a_sign0 = 4'd16; a_sign1 = 4'd14; a_sign2 = 4'd12; a_sign3 = 4'd11;
b_sign0 = 4'd2; b_sign1 = 4'd15; b_sign2 = 4'd0; b_sign3 = 4'd11;
@(posedge clk_i);
a_mant0 = 8'd118; a_mant1 = 8'd29; a_mant2 = 8'd67; a_mant3 = 8'd70;
b_mant0 = 8'd100; b_mant1 = 8'd171; b_mant2 = 8'd131; b_mant3 = 8'd28;
a_exp0 = 10'd58; a_exp1 = 10'd426; a_exp2 = 10'd378; a_exp3 = 10'd564;
b_exp0 = 10'd626; b_exp1 = 10'd248; b_exp2 = 10'd984; b_exp3 = 10'd948;
a_sign0 = 4'd4; a_sign1 = 4'd12; a_sign2 = 4'd16; a_sign3 = 4'd10;
b_sign0 = 4'd11; b_sign1 = 4'd5; b_sign2 = 4'd16; b_sign3 = 4'd2;
@(posedge clk_i);
a_mant0 = 8'd201; a_mant1 = 8'd48; a_mant2 = 8'd7; a_mant3 = 8'd14;
b_mant0 = 8'd49; b_mant1 = 8'd162; b_mant2 = 8'd40; b_mant3 = 8'd86;
a_exp0 = 10'd913; a_exp1 = 10'd720; a_exp2 = 10'd835; a_exp3 = 10'd907;
b_exp0 = 10'd276; b_exp1 = 10'd540; b_exp2 = 10'd570; b_exp3 = 10'd1010;
a_sign0 = 4'd1; a_sign1 = 4'd9; a_sign2 = 4'd16; a_sign3 = 4'd2;
b_sign0 = 4'd9; b_sign1 = 4'd0; b_sign2 = 4'd7; b_sign3 = 4'd10;
@(posedge clk_i);
a_mant0 = 8'd33; a_mant1 = 8'd120; a_mant2 = 8'd37; a_mant3 = 8'd39;
b_mant0 = 8'd146; b_mant1 = 8'd102; b_mant2 = 8'd204; b_mant3 = 8'd189;
a_exp0 = 10'd335; a_exp1 = 10'd550; a_exp2 = 10'd677; a_exp3 = 10'd130;
b_exp0 = 10'd864; b_exp1 = 10'd499; b_exp2 = 10'd174; b_exp3 = 10'd846;
a_sign0 = 4'd1; a_sign1 = 4'd10; a_sign2 = 4'd11; a_sign3 = 4'd3;
b_sign0 = 4'd15; b_sign1 = 4'd4; b_sign2 = 4'd16; b_sign3 = 4'd14;
@(posedge clk_i);
a_mant0 = 8'd181; a_mant1 = 8'd152; a_mant2 = 8'd28; a_mant3 = 8'd71;
b_mant0 = 8'd204; b_mant1 = 8'd96; b_mant2 = 8'd215; b_mant3 = 8'd5;
a_exp0 = 10'd634; a_exp1 = 10'd1002; a_exp2 = 10'd725; a_exp3 = 10'd870;
b_exp0 = 10'd781; b_exp1 = 10'd932; b_exp2 = 10'd896; b_exp3 = 10'd465;
a_sign0 = 4'd16; a_sign1 = 4'd5; a_sign2 = 4'd10; a_sign3 = 4'd10;
b_sign0 = 4'd11; b_sign1 = 4'd13; b_sign2 = 4'd4; b_sign3 = 4'd5;
@(posedge clk_i);
a_mant0 = 8'd123; a_mant1 = 8'd201; a_mant2 = 8'd178; a_mant3 = 8'd120;
b_mant0 = 8'd170; b_mant1 = 8'd0; b_mant2 = 8'd94; b_mant3 = 8'd155;
a_exp0 = 10'd572; a_exp1 = 10'd1009; a_exp2 = 10'd952; a_exp3 = 10'd476;
b_exp0 = 10'd255; b_exp1 = 10'd814; b_exp2 = 10'd399; b_exp3 = 10'd892;
a_sign0 = 4'd11; a_sign1 = 4'd10; a_sign2 = 4'd5; a_sign3 = 4'd3;
b_sign0 = 4'd5; b_sign1 = 4'd2; b_sign2 = 4'd10; b_sign3 = 4'd4;
@(posedge clk_i);
shared_exps0 = 8'd131;
shared_exps1 = 8'd123;
a_mant0 = 8'd196; a_mant1 = 8'd122; a_mant2 = 8'd249; a_mant3 = 8'd244;
b_mant0 = 8'd121; b_mant1 = 8'd223; b_mant2 = 8'd130; b_mant3 = 8'd164;
a_exp0 = 10'd29; a_exp1 = 10'd759; a_exp2 = 10'd365; a_exp3 = 10'd606;
b_exp0 = 10'd831; b_exp1 = 10'd542; b_exp2 = 10'd24; b_exp3 = 10'd684;
a_sign0 = 4'd0; a_sign1 = 4'd1; a_sign2 = 4'd11; a_sign3 = 4'd11;
b_sign0 = 4'd15; b_sign1 = 4'd9; b_sign2 = 4'd16; b_sign3 = 4'd15;
@(posedge clk_i);
a_mant0 = 8'd125; a_mant1 = 8'd166; a_mant2 = 8'd237; a_mant3 = 8'd125;
b_mant0 = 8'd205; b_mant1 = 8'd250; b_mant2 = 8'd43; b_mant3 = 8'd68;
a_exp0 = 10'd151; a_exp1 = 10'd334; a_exp2 = 10'd377; a_exp3 = 10'd961;
b_exp0 = 10'd655; b_exp1 = 10'd607; b_exp2 = 10'd886; b_exp3 = 10'd679;
a_sign0 = 4'd8; a_sign1 = 4'd12; a_sign2 = 4'd11; a_sign3 = 4'd14;
b_sign0 = 4'd7; b_sign1 = 4'd15; b_sign2 = 4'd3; b_sign3 = 4'd15;
@(posedge clk_i);
a_mant0 = 8'd250; a_mant1 = 8'd17; a_mant2 = 8'd97; a_mant3 = 8'd30;
b_mant0 = 8'd21; b_mant1 = 8'd14; b_mant2 = 8'd107; b_mant3 = 8'd5;
a_exp0 = 10'd896; a_exp1 = 10'd251; a_exp2 = 10'd723; a_exp3 = 10'd218;
b_exp0 = 10'd260; b_exp1 = 10'd211; b_exp2 = 10'd824; b_exp3 = 10'd782;
a_sign0 = 4'd8; a_sign1 = 4'd6; a_sign2 = 4'd2; a_sign3 = 4'd3;
b_sign0 = 4'd14; b_sign1 = 4'd8; b_sign2 = 4'd12; b_sign3 = 4'd15;
@(posedge clk_i);
a_mant0 = 8'd254; a_mant1 = 8'd85; a_mant2 = 8'd91; a_mant3 = 8'd244;
b_mant0 = 8'd192; b_mant1 = 8'd219; b_mant2 = 8'd135; b_mant3 = 8'd1;
a_exp0 = 10'd256; a_exp1 = 10'd36; a_exp2 = 10'd968; a_exp3 = 10'd649;
b_exp0 = 10'd119; b_exp1 = 10'd1011; b_exp2 = 10'd101; b_exp3 = 10'd960;
a_sign0 = 4'd13; a_sign1 = 4'd12; a_sign2 = 4'd2; a_sign3 = 4'd5;
b_sign0 = 4'd4; b_sign1 = 4'd3; b_sign2 = 4'd4; b_sign3 = 4'd1;
@(posedge clk_i);
a_mant0 = 8'd139; a_mant1 = 8'd58; a_mant2 = 8'd195; a_mant3 = 8'd199;
b_mant0 = 8'd204; b_mant1 = 8'd132; b_mant2 = 8'd66; b_mant3 = 8'd246;
a_exp0 = 10'd447; a_exp1 = 10'd828; a_exp2 = 10'd628; a_exp3 = 10'd632;
b_exp0 = 10'd199; b_exp1 = 10'd320; b_exp2 = 10'd382; b_exp3 = 10'd953;
a_sign0 = 4'd6; a_sign1 = 4'd12; a_sign2 = 4'd7; a_sign3 = 4'd2;
b_sign0 = 4'd3; b_sign1 = 4'd12; b_sign2 = 4'd11; b_sign3 = 4'd6;
@(posedge clk_i);
a_mant0 = 8'd40; a_mant1 = 8'd203; a_mant2 = 8'd50; a_mant3 = 8'd72;
b_mant0 = 8'd68; b_mant1 = 8'd198; b_mant2 = 8'd22; b_mant3 = 8'd154;
a_exp0 = 10'd692; a_exp1 = 10'd509; a_exp2 = 10'd438; a_exp3 = 10'd213;
b_exp0 = 10'd252; b_exp1 = 10'd322; b_exp2 = 10'd667; b_exp3 = 10'd589;
a_sign0 = 4'd13; a_sign1 = 4'd16; a_sign2 = 4'd1; a_sign3 = 4'd14;
b_sign0 = 4'd14; b_sign1 = 4'd1; b_sign2 = 4'd0; b_sign3 = 4'd3;
@(posedge clk_i);
a_mant0 = 8'd127; a_mant1 = 8'd227; a_mant2 = 8'd28; a_mant3 = 8'd43;
b_mant0 = 8'd128; b_mant1 = 8'd9; b_mant2 = 8'd155; b_mant3 = 8'd245;
a_exp0 = 10'd217; a_exp1 = 10'd126; a_exp2 = 10'd943; a_exp3 = 10'd1008;
b_exp0 = 10'd347; b_exp1 = 10'd63; b_exp2 = 10'd629; b_exp3 = 10'd1019;
a_sign0 = 4'd0; a_sign1 = 4'd3; a_sign2 = 4'd8; a_sign3 = 4'd10;
b_sign0 = 4'd16; b_sign1 = 4'd3; b_sign2 = 4'd5; b_sign3 = 4'd3;
@(posedge clk_i);
a_mant0 = 8'd33; a_mant1 = 8'd57; a_mant2 = 8'd8; a_mant3 = 8'd107;
b_mant0 = 8'd131; b_mant1 = 8'd101; b_mant2 = 8'd67; b_mant3 = 8'd81;
a_exp0 = 10'd852; a_exp1 = 10'd583; a_exp2 = 10'd755; a_exp3 = 10'd661;
b_exp0 = 10'd920; b_exp1 = 10'd334; b_exp2 = 10'd719; b_exp3 = 10'd88;
a_sign0 = 4'd9; a_sign1 = 4'd3; a_sign2 = 4'd15; a_sign3 = 4'd8;
b_sign0 = 4'd14; b_sign1 = 4'd12; b_sign2 = 4'd9; b_sign3 = 4'd12;
@(posedge clk_i);
shared_exps0 = 8'd139;
shared_exps1 = 8'd148;
rstn = 0;
@(posedge clk_i);
rstn = 1;
a_mant0 = 8'd31; a_mant1 = 8'd64; a_mant2 = 8'd20; a_mant3 = 8'd232;
b_mant0 = 8'd148; b_mant1 = 8'd78; b_mant2 = 8'd184; b_mant3 = 8'd144;
a_exp0 = 10'd279; a_exp1 = 10'd49; a_exp2 = 10'd322; a_exp3 = 10'd279;
b_exp0 = 10'd402; b_exp1 = 10'd893; b_exp2 = 10'd277; b_exp3 = 10'd12;
a_sign0 = 4'd15; a_sign1 = 4'd6; a_sign2 = 4'd2; a_sign3 = 4'd16;
b_sign0 = 4'd16; b_sign1 = 4'd3; b_sign2 = 4'd12; b_sign3 = 4'd5;
@(posedge clk_i);
a_mant0 = 8'd207; a_mant1 = 8'd82; a_mant2 = 8'd95; a_mant3 = 8'd72;
b_mant0 = 8'd158; b_mant1 = 8'd116; b_mant2 = 8'd8; b_mant3 = 8'd15;
a_exp0 = 10'd455; a_exp1 = 10'd43; a_exp2 = 10'd598; a_exp3 = 10'd464;
b_exp0 = 10'd204; b_exp1 = 10'd609; b_exp2 = 10'd909; b_exp3 = 10'd743;
a_sign0 = 4'd14; a_sign1 = 4'd7; a_sign2 = 4'd12; a_sign3 = 4'd9;
b_sign0 = 4'd10; b_sign1 = 4'd16; b_sign2 = 4'd4; b_sign3 = 4'd8;
@(posedge clk_i);
a_mant0 = 8'd167; a_mant1 = 8'd111; a_mant2 = 8'd96; a_mant3 = 8'd39;
b_mant0 = 8'd150; b_mant1 = 8'd136; b_mant2 = 8'd71; b_mant3 = 8'd135;
a_exp0 = 10'd853; a_exp1 = 10'd503; a_exp2 = 10'd886; a_exp3 = 10'd640;
b_exp0 = 10'd12; b_exp1 = 10'd457; b_exp2 = 10'd399; b_exp3 = 10'd588;
a_sign0 = 4'd9; a_sign1 = 4'd8; a_sign2 = 4'd10; a_sign3 = 4'd2;
b_sign0 = 4'd9; b_sign1 = 4'd8; b_sign2 = 4'd4; b_sign3 = 4'd6;
@(posedge clk_i);
a_mant0 = 8'd78; a_mant1 = 8'd141; a_mant2 = 8'd242; a_mant3 = 8'd172;
b_mant0 = 8'd118; b_mant1 = 8'd249; b_mant2 = 8'd156; b_mant3 = 8'd117;
a_exp0 = 10'd716; a_exp1 = 10'd880; a_exp2 = 10'd905; a_exp3 = 10'd994;
b_exp0 = 10'd195; b_exp1 = 10'd340; b_exp2 = 10'd977; b_exp3 = 10'd864;
a_sign0 = 4'd8; a_sign1 = 4'd14; a_sign2 = 4'd14; a_sign3 = 4'd13;
b_sign0 = 4'd2; b_sign1 = 4'd1; b_sign2 = 4'd14; b_sign3 = 4'd13;
@(posedge clk_i);
a_mant0 = 8'd169; a_mant1 = 8'd184; a_mant2 = 8'd55; a_mant3 = 8'd13;
b_mant0 = 8'd32; b_mant1 = 8'd112; b_mant2 = 8'd79; b_mant3 = 8'd4;
a_exp0 = 10'd158; a_exp1 = 10'd810; a_exp2 = 10'd621; a_exp3 = 10'd277;
b_exp0 = 10'd357; b_exp1 = 10'd124; b_exp2 = 10'd582; b_exp3 = 10'd1014;
a_sign0 = 4'd4; a_sign1 = 4'd4; a_sign2 = 4'd14; a_sign3 = 4'd10;
b_sign0 = 4'd3; b_sign1 = 4'd0; b_sign2 = 4'd3; b_sign3 = 4'd13;
@(posedge clk_i);
a_mant0 = 8'd161; a_mant1 = 8'd212; a_mant2 = 8'd7; a_mant3 = 8'd214;
b_mant0 = 8'd166; b_mant1 = 8'd190; b_mant2 = 8'd62; b_mant3 = 8'd79;
a_exp0 = 10'd329; a_exp1 = 10'd841; a_exp2 = 10'd146; a_exp3 = 10'd188;
b_exp0 = 10'd757; b_exp1 = 10'd64; b_exp2 = 10'd184; b_exp3 = 10'd556;
a_sign0 = 4'd12; a_sign1 = 4'd13; a_sign2 = 4'd9; a_sign3 = 4'd7;
b_sign0 = 4'd7; b_sign1 = 4'd14; b_sign2 = 4'd1; b_sign3 = 4'd6;
@(posedge clk_i);
a_mant0 = 8'd105; a_mant1 = 8'd135; a_mant2 = 8'd144; a_mant3 = 8'd52;
b_mant0 = 8'd195; b_mant1 = 8'd233; b_mant2 = 8'd46; b_mant3 = 8'd134;
a_exp0 = 10'd796; a_exp1 = 10'd89; a_exp2 = 10'd1012; a_exp3 = 10'd656;
b_exp0 = 10'd87; b_exp1 = 10'd837; b_exp2 = 10'd730; b_exp3 = 10'd678;
a_sign0 = 4'd4; a_sign1 = 4'd1; a_sign2 = 4'd10; a_sign3 = 4'd16;
b_sign0 = 4'd11; b_sign1 = 4'd15; b_sign2 = 4'd11; b_sign3 = 4'd16;
@(posedge clk_i);
shared_exps0 = 8'd101;
shared_exps1 = 8'd114;
a_mant0 = 8'd158; a_mant1 = 8'd0; a_mant2 = 8'd74; a_mant3 = 8'd93;
b_mant0 = 8'd38; b_mant1 = 8'd141; b_mant2 = 8'd141; b_mant3 = 8'd74;
a_exp0 = 10'd147; a_exp1 = 10'd148; a_exp2 = 10'd481; a_exp3 = 10'd560;
b_exp0 = 10'd859; b_exp1 = 10'd194; b_exp2 = 10'd784; b_exp3 = 10'd96;
a_sign0 = 4'd3; a_sign1 = 4'd2; a_sign2 = 4'd14; a_sign3 = 4'd3;
b_sign0 = 4'd16; b_sign1 = 4'd13; b_sign2 = 4'd12; b_sign3 = 4'd7;
@(posedge clk_i);
a_mant0 = 8'd11; a_mant1 = 8'd229; a_mant2 = 8'd10; a_mant3 = 8'd55;
b_mant0 = 8'd29; b_mant1 = 8'd49; b_mant2 = 8'd30; b_mant3 = 8'd7;
a_exp0 = 10'd779; a_exp1 = 10'd633; a_exp2 = 10'd373; a_exp3 = 10'd637;
b_exp0 = 10'd435; b_exp1 = 10'd889; b_exp2 = 10'd566; b_exp3 = 10'd812;
a_sign0 = 4'd5; a_sign1 = 4'd3; a_sign2 = 4'd14; a_sign3 = 4'd4;
b_sign0 = 4'd16; b_sign1 = 4'd5; b_sign2 = 4'd0; b_sign3 = 4'd2;
@(posedge clk_i);
a_mant0 = 8'd238; a_mant1 = 8'd151; a_mant2 = 8'd25; a_mant3 = 8'd47;
b_mant0 = 8'd47; b_mant1 = 8'd27; b_mant2 = 8'd24; b_mant3 = 8'd119;
a_exp0 = 10'd345; a_exp1 = 10'd166; a_exp2 = 10'd109; a_exp3 = 10'd935;
b_exp0 = 10'd174; b_exp1 = 10'd322; b_exp2 = 10'd851; b_exp3 = 10'd576;
a_sign0 = 4'd8; a_sign1 = 4'd13; a_sign2 = 4'd11; a_sign3 = 4'd1;
b_sign0 = 4'd0; b_sign1 = 4'd7; b_sign2 = 4'd4; b_sign3 = 4'd0;
@(posedge clk_i);
a_mant0 = 8'd121; a_mant1 = 8'd67; a_mant2 = 8'd68; a_mant3 = 8'd210;
b_mant0 = 8'd254; b_mant1 = 8'd47; b_mant2 = 8'd64; b_mant3 = 8'd94;
a_exp0 = 10'd602; a_exp1 = 10'd68; a_exp2 = 10'd744; a_exp3 = 10'd124;
b_exp0 = 10'd97; b_exp1 = 10'd88; b_exp2 = 10'd26; b_exp3 = 10'd568;
a_sign0 = 4'd9; a_sign1 = 4'd8; a_sign2 = 4'd8; a_sign3 = 4'd0;
b_sign0 = 4'd15; b_sign1 = 4'd5; b_sign2 = 4'd10; b_sign3 = 4'd14;
@(posedge clk_i);
a_mant0 = 8'd35; a_mant1 = 8'd40; a_mant2 = 8'd64; a_mant3 = 8'd58;
b_mant0 = 8'd117; b_mant1 = 8'd98; b_mant2 = 8'd87; b_mant3 = 8'd106;
a_exp0 = 10'd568; a_exp1 = 10'd97; a_exp2 = 10'd621; a_exp3 = 10'd152;
b_exp0 = 10'd399; b_exp1 = 10'd981; b_exp2 = 10'd189; b_exp3 = 10'd493;
a_sign0 = 4'd16; a_sign1 = 4'd15; a_sign2 = 4'd5; a_sign3 = 4'd13;
b_sign0 = 4'd6; b_sign1 = 4'd11; b_sign2 = 4'd16; b_sign3 = 4'd8;
@(posedge clk_i);
a_mant0 = 8'd77; a_mant1 = 8'd146; a_mant2 = 8'd98; a_mant3 = 8'd23;
b_mant0 = 8'd252; b_mant1 = 8'd78; b_mant2 = 8'd149; b_mant3 = 8'd229;
a_exp0 = 10'd380; a_exp1 = 10'd453; a_exp2 = 10'd763; a_exp3 = 10'd980;
b_exp0 = 10'd587; b_exp1 = 10'd368; b_exp2 = 10'd770; b_exp3 = 10'd148;
a_sign0 = 4'd6; a_sign1 = 4'd15; a_sign2 = 4'd1; a_sign3 = 4'd12;
b_sign0 = 4'd5; b_sign1 = 4'd12; b_sign2 = 4'd4; b_sign3 = 4'd12;
@(posedge clk_i);
a_mant0 = 8'd10; a_mant1 = 8'd192; a_mant2 = 8'd35; a_mant3 = 8'd237;
b_mant0 = 8'd122; b_mant1 = 8'd171; b_mant2 = 8'd78; b_mant3 = 8'd114;
a_exp0 = 10'd556; a_exp1 = 10'd878; a_exp2 = 10'd384; a_exp3 = 10'd251;
b_exp0 = 10'd579; b_exp1 = 10'd750; b_exp2 = 10'd817; b_exp3 = 10'd33;
a_sign0 = 4'd11; a_sign1 = 4'd11; a_sign2 = 4'd15; a_sign3 = 4'd10;
b_sign0 = 4'd4; b_sign1 = 4'd7; b_sign2 = 4'd13; b_sign3 = 4'd0;
@(posedge clk_i);
a_mant0 = 8'd200; a_mant1 = 8'd2; a_mant2 = 8'd137; a_mant3 = 8'd126;
b_mant0 = 8'd78; b_mant1 = 8'd188; b_mant2 = 8'd197; b_mant3 = 8'd240;
a_exp0 = 10'd475; a_exp1 = 10'd911; a_exp2 = 10'd947; a_exp3 = 10'd453;
b_exp0 = 10'd920; b_exp1 = 10'd247; b_exp2 = 10'd875; b_exp3 = 10'd98;
a_sign0 = 4'd16; a_sign1 = 4'd10; a_sign2 = 4'd7; a_sign3 = 4'd16;
b_sign0 = 4'd8; b_sign1 = 4'd0; b_sign2 = 4'd10; b_sign3 = 4'd2;
@(posedge clk_i);
shared_exps0 = 8'd120;
shared_exps1 = 8'd121;
a_mant0 = 8'd127; a_mant1 = 8'd81; a_mant2 = 8'd127; a_mant3 = 8'd97;
b_mant0 = 8'd60; b_mant1 = 8'd222; b_mant2 = 8'd138; b_mant3 = 8'd29;
a_exp0 = 10'd986; a_exp1 = 10'd504; a_exp2 = 10'd364; a_exp3 = 10'd211;
b_exp0 = 10'd476; b_exp1 = 10'd321; b_exp2 = 10'd239; b_exp3 = 10'd138;
a_sign0 = 4'd4; a_sign1 = 4'd5; a_sign2 = 4'd4; a_sign3 = 4'd3;
b_sign0 = 4'd9; b_sign1 = 4'd1; b_sign2 = 4'd9; b_sign3 = 4'd5;
@(posedge clk_i);
a_mant0 = 8'd255; a_mant1 = 8'd209; a_mant2 = 8'd75; a_mant3 = 8'd5;
b_mant0 = 8'd194; b_mant1 = 8'd44; b_mant2 = 8'd164; b_mant3 = 8'd185;
a_exp0 = 10'd847; a_exp1 = 10'd697; a_exp2 = 10'd1012; a_exp3 = 10'd141;
b_exp0 = 10'd826; b_exp1 = 10'd641; b_exp2 = 10'd13; b_exp3 = 10'd827;
a_sign0 = 4'd12; a_sign1 = 4'd11; a_sign2 = 4'd7; a_sign3 = 4'd11;
b_sign0 = 4'd1; b_sign1 = 4'd10; b_sign2 = 4'd0; b_sign3 = 4'd2;
@(posedge clk_i);
a_mant0 = 8'd125; a_mant1 = 8'd218; a_mant2 = 8'd214; a_mant3 = 8'd129;
b_mant0 = 8'd107; b_mant1 = 8'd144; b_mant2 = 8'd28; b_mant3 = 8'd216;
a_exp0 = 10'd966; a_exp1 = 10'd1013; a_exp2 = 10'd282; a_exp3 = 10'd470;
b_exp0 = 10'd541; b_exp1 = 10'd915; b_exp2 = 10'd642; b_exp3 = 10'd353;
a_sign0 = 4'd0; a_sign1 = 4'd15; a_sign2 = 4'd5; a_sign3 = 4'd5;
b_sign0 = 4'd6; b_sign1 = 4'd14; b_sign2 = 4'd8; b_sign3 = 4'd5;
@(posedge clk_i);
a_mant0 = 8'd220; a_mant1 = 8'd36; a_mant2 = 8'd60; a_mant3 = 8'd201;
b_mant0 = 8'd143; b_mant1 = 8'd189; b_mant2 = 8'd66; b_mant3 = 8'd48;
a_exp0 = 10'd977; a_exp1 = 10'd843; a_exp2 = 10'd184; a_exp3 = 10'd683;
b_exp0 = 10'd73; b_exp1 = 10'd839; b_exp2 = 10'd255; b_exp3 = 10'd842;
a_sign0 = 4'd5; a_sign1 = 4'd13; a_sign2 = 4'd4; a_sign3 = 4'd6;
b_sign0 = 4'd13; b_sign1 = 4'd5; b_sign2 = 4'd16; b_sign3 = 4'd12;
@(posedge clk_i);
a_mant0 = 8'd82; a_mant1 = 8'd109; a_mant2 = 8'd37; a_mant3 = 8'd70;
b_mant0 = 8'd195; b_mant1 = 8'd168; b_mant2 = 8'd200; b_mant3 = 8'd144;
a_exp0 = 10'd199; a_exp1 = 10'd477; a_exp2 = 10'd274; a_exp3 = 10'd263;
b_exp0 = 10'd216; b_exp1 = 10'd236; b_exp2 = 10'd280; b_exp3 = 10'd65;
a_sign0 = 4'd11; a_sign1 = 4'd9; a_sign2 = 4'd2; a_sign3 = 4'd14;
b_sign0 = 4'd12; b_sign1 = 4'd7; b_sign2 = 4'd10; b_sign3 = 4'd13;
@(posedge clk_i);
a_mant0 = 8'd71; a_mant1 = 8'd61; a_mant2 = 8'd199; a_mant3 = 8'd107;
b_mant0 = 8'd63; b_mant1 = 8'd98; b_mant2 = 8'd156; b_mant3 = 8'd118;
a_exp0 = 10'd446; a_exp1 = 10'd282; a_exp2 = 10'd850; a_exp3 = 10'd8;
b_exp0 = 10'd723; b_exp1 = 10'd408; b_exp2 = 10'd431; b_exp3 = 10'd633;
a_sign0 = 4'd0; a_sign1 = 4'd4; a_sign2 = 4'd15; a_sign3 = 4'd3;
b_sign0 = 4'd0; b_sign1 = 4'd2; b_sign2 = 4'd15; b_sign3 = 4'd1;
@(posedge clk_i);
a_mant0 = 8'd228; a_mant1 = 8'd48; a_mant2 = 8'd59; a_mant3 = 8'd13;
b_mant0 = 8'd242; b_mant1 = 8'd130; b_mant2 = 8'd102; b_mant3 = 8'd34;
a_exp0 = 10'd246; a_exp1 = 10'd258; a_exp2 = 10'd1018; a_exp3 = 10'd330;
b_exp0 = 10'd751; b_exp1 = 10'd493; b_exp2 = 10'd611; b_exp3 = 10'd622;
a_sign0 = 4'd2; a_sign1 = 4'd8; a_sign2 = 4'd13; a_sign3 = 4'd4;
b_sign0 = 4'd12; b_sign1 = 4'd3; b_sign2 = 4'd7; b_sign3 = 4'd5;
@(posedge clk_i);
a_mant0 = 8'd91; a_mant1 = 8'd212; a_mant2 = 8'd83; a_mant3 = 8'd136;
b_mant0 = 8'd241; b_mant1 = 8'd144; b_mant2 = 8'd162; b_mant3 = 8'd211;
a_exp0 = 10'd830; a_exp1 = 10'd658; a_exp2 = 10'd576; a_exp3 = 10'd339;
b_exp0 = 10'd818; b_exp1 = 10'd665; b_exp2 = 10'd193; b_exp3 = 10'd285;
a_sign0 = 4'd12; a_sign1 = 4'd11; a_sign2 = 4'd1; a_sign3 = 4'd6;
b_sign0 = 4'd11; b_sign1 = 4'd3; b_sign2 = 4'd10; b_sign3 = 4'd4;
@(posedge clk_i);
shared_exps0 = 8'd142;
shared_exps1 = 8'd161;
a_mant0 = 8'd203; a_mant1 = 8'd230; a_mant2 = 8'd255; a_mant3 = 8'd13;
b_mant0 = 8'd106; b_mant1 = 8'd3; b_mant2 = 8'd93; b_mant3 = 8'd34;
a_exp0 = 10'd167; a_exp1 = 10'd303; a_exp2 = 10'd269; a_exp3 = 10'd630;
b_exp0 = 10'd897; b_exp1 = 10'd231; b_exp2 = 10'd847; b_exp3 = 10'd450;
a_sign0 = 4'd13; a_sign1 = 4'd2; a_sign2 = 4'd4; a_sign3 = 4'd14;
b_sign0 = 4'd9; b_sign1 = 4'd12; b_sign2 = 4'd5; b_sign3 = 4'd16;
@(posedge clk_i);
a_mant0 = 8'd165; a_mant1 = 8'd128; a_mant2 = 8'd185; a_mant3 = 8'd118;
b_mant0 = 8'd196; b_mant1 = 8'd51; b_mant2 = 8'd195; b_mant3 = 8'd126;
a_exp0 = 10'd912; a_exp1 = 10'd694; a_exp2 = 10'd363; a_exp3 = 10'd949;
b_exp0 = 10'd158; b_exp1 = 10'd631; b_exp2 = 10'd413; b_exp3 = 10'd909;
a_sign0 = 4'd13; a_sign1 = 4'd3; a_sign2 = 4'd15; a_sign3 = 4'd4;
b_sign0 = 4'd13; b_sign1 = 4'd9; b_sign2 = 4'd2; b_sign3 = 4'd3;
@(posedge clk_i);
a_mant0 = 8'd235; a_mant1 = 8'd127; a_mant2 = 8'd121; a_mant3 = 8'd218;
b_mant0 = 8'd196; b_mant1 = 8'd97; b_mant2 = 8'd226; b_mant3 = 8'd87;
a_exp0 = 10'd478; a_exp1 = 10'd474; a_exp2 = 10'd733; a_exp3 = 10'd163;
b_exp0 = 10'd474; b_exp1 = 10'd172; b_exp2 = 10'd314; b_exp3 = 10'd944;
a_sign0 = 4'd12; a_sign1 = 4'd16; a_sign2 = 4'd16; a_sign3 = 4'd8;
b_sign0 = 4'd11; b_sign1 = 4'd13; b_sign2 = 4'd13; b_sign3 = 4'd0;
@(posedge clk_i);
a_mant0 = 8'd231; a_mant1 = 8'd33; a_mant2 = 8'd215; a_mant3 = 8'd8;
b_mant0 = 8'd115; b_mant1 = 8'd162; b_mant2 = 8'd58; b_mant3 = 8'd130;
a_exp0 = 10'd755; a_exp1 = 10'd890; a_exp2 = 10'd347; a_exp3 = 10'd170;
b_exp0 = 10'd651; b_exp1 = 10'd14; b_exp2 = 10'd308; b_exp3 = 10'd618;
a_sign0 = 4'd7; a_sign1 = 4'd7; a_sign2 = 4'd3; a_sign3 = 4'd0;
b_sign0 = 4'd12; b_sign1 = 4'd3; b_sign2 = 4'd15; b_sign3 = 4'd15;
@(posedge clk_i);
a_mant0 = 8'd245; a_mant1 = 8'd91; a_mant2 = 8'd233; a_mant3 = 8'd93;
b_mant0 = 8'd106; b_mant1 = 8'd203; b_mant2 = 8'd83; b_mant3 = 8'd245;
a_exp0 = 10'd508; a_exp1 = 10'd119; a_exp2 = 10'd62; a_exp3 = 10'd453;
b_exp0 = 10'd344; b_exp1 = 10'd422; b_exp2 = 10'd824; b_exp3 = 10'd954;
a_sign0 = 4'd15; a_sign1 = 4'd16; a_sign2 = 4'd6; a_sign3 = 4'd14;
b_sign0 = 4'd3; b_sign1 = 4'd3; b_sign2 = 4'd8; b_sign3 = 4'd6;
@(posedge clk_i);
a_mant0 = 8'd46; a_mant1 = 8'd187; a_mant2 = 8'd224; a_mant3 = 8'd149;
b_mant0 = 8'd126; b_mant1 = 8'd117; b_mant2 = 8'd95; b_mant3 = 8'd154;
a_exp0 = 10'd977; a_exp1 = 10'd679; a_exp2 = 10'd597; a_exp3 = 10'd303;
b_exp0 = 10'd175; b_exp1 = 10'd873; b_exp2 = 10'd438; b_exp3 = 10'd69;
a_sign0 = 4'd5; a_sign1 = 4'd4; a_sign2 = 4'd9; a_sign3 = 4'd5;
b_sign0 = 4'd1; b_sign1 = 4'd13; b_sign2 = 4'd13; b_sign3 = 4'd15;
@(posedge clk_i);
a_mant0 = 8'd118; a_mant1 = 8'd44; a_mant2 = 8'd241; a_mant3 = 8'd105;
b_mant0 = 8'd222; b_mant1 = 8'd219; b_mant2 = 8'd15; b_mant3 = 8'd42;
a_exp0 = 10'd257; a_exp1 = 10'd380; a_exp2 = 10'd689; a_exp3 = 10'd26;
b_exp0 = 10'd420; b_exp1 = 10'd703; b_exp2 = 10'd930; b_exp3 = 10'd112;
a_sign0 = 4'd12; a_sign1 = 4'd14; a_sign2 = 4'd12; a_sign3 = 4'd2;
b_sign0 = 4'd8; b_sign1 = 4'd3; b_sign2 = 4'd16; b_sign3 = 4'd2;
@(posedge clk_i);
a_mant0 = 8'd155; a_mant1 = 8'd196; a_mant2 = 8'd152; a_mant3 = 8'd65;
b_mant0 = 8'd88; b_mant1 = 8'd145; b_mant2 = 8'd116; b_mant3 = 8'd221;
a_exp0 = 10'd601; a_exp1 = 10'd827; a_exp2 = 10'd947; a_exp3 = 10'd483;
b_exp0 = 10'd665; b_exp1 = 10'd144; b_exp2 = 10'd72; b_exp3 = 10'd630;
a_sign0 = 4'd14; a_sign1 = 4'd11; a_sign2 = 4'd16; a_sign3 = 4'd0;
b_sign0 = 4'd11; b_sign1 = 4'd8; b_sign2 = 4'd1; b_sign3 = 4'd15;
@(posedge clk_i);
shared_exps0 = 8'd134;
shared_exps1 = 8'd151;
rstn = 0;
@(posedge clk_i);
rstn = 1;
a_mant0 = 8'd235; a_mant1 = 8'd130; a_mant2 = 8'd47; a_mant3 = 8'd1;
b_mant0 = 8'd75; b_mant1 = 8'd124; b_mant2 = 8'd124; b_mant3 = 8'd178;
a_exp0 = 10'd852; a_exp1 = 10'd682; a_exp2 = 10'd980; a_exp3 = 10'd879;
b_exp0 = 10'd514; b_exp1 = 10'd257; b_exp2 = 10'd742; b_exp3 = 10'd712;
a_sign0 = 4'd6; a_sign1 = 4'd10; a_sign2 = 4'd14; a_sign3 = 4'd8;
b_sign0 = 4'd16; b_sign1 = 4'd11; b_sign2 = 4'd12; b_sign3 = 4'd15;
@(posedge clk_i);
a_mant0 = 8'd78; a_mant1 = 8'd109; a_mant2 = 8'd61; a_mant3 = 8'd217;
b_mant0 = 8'd101; b_mant1 = 8'd195; b_mant2 = 8'd250; b_mant3 = 8'd52;
a_exp0 = 10'd397; a_exp1 = 10'd369; a_exp2 = 10'd71; a_exp3 = 10'd858;
b_exp0 = 10'd684; b_exp1 = 10'd204; b_exp2 = 10'd858; b_exp3 = 10'd645;
a_sign0 = 4'd13; a_sign1 = 4'd5; a_sign2 = 4'd16; a_sign3 = 4'd7;
b_sign0 = 4'd2; b_sign1 = 4'd3; b_sign2 = 4'd8; b_sign3 = 4'd11;
@(posedge clk_i);
a_mant0 = 8'd219; a_mant1 = 8'd253; a_mant2 = 8'd253; a_mant3 = 8'd38;
b_mant0 = 8'd74; b_mant1 = 8'd102; b_mant2 = 8'd150; b_mant3 = 8'd21;
a_exp0 = 10'd350; a_exp1 = 10'd440; a_exp2 = 10'd512; a_exp3 = 10'd473;
b_exp0 = 10'd340; b_exp1 = 10'd39; b_exp2 = 10'd991; b_exp3 = 10'd777;
a_sign0 = 4'd5; a_sign1 = 4'd13; a_sign2 = 4'd15; a_sign3 = 4'd3;
b_sign0 = 4'd6; b_sign1 = 4'd6; b_sign2 = 4'd3; b_sign3 = 4'd12;
@(posedge clk_i);
a_mant0 = 8'd91; a_mant1 = 8'd40; a_mant2 = 8'd142; a_mant3 = 8'd242;
b_mant0 = 8'd100; b_mant1 = 8'd197; b_mant2 = 8'd96; b_mant3 = 8'd230;
a_exp0 = 10'd429; a_exp1 = 10'd417; a_exp2 = 10'd515; a_exp3 = 10'd142;
b_exp0 = 10'd540; b_exp1 = 10'd79; b_exp2 = 10'd488; b_exp3 = 10'd328;
a_sign0 = 4'd16; a_sign1 = 4'd16; a_sign2 = 4'd11; a_sign3 = 4'd3;
b_sign0 = 4'd11; b_sign1 = 4'd8; b_sign2 = 4'd3; b_sign3 = 4'd6;
@(posedge clk_i);
a_mant0 = 8'd160; a_mant1 = 8'd56; a_mant2 = 8'd152; a_mant3 = 8'd197;
b_mant0 = 8'd31; b_mant1 = 8'd5; b_mant2 = 8'd180; b_mant3 = 8'd216;
a_exp0 = 10'd504; a_exp1 = 10'd957; a_exp2 = 10'd732; a_exp3 = 10'd686;
b_exp0 = 10'd836; b_exp1 = 10'd800; b_exp2 = 10'd526; b_exp3 = 10'd177;
a_sign0 = 4'd11; a_sign1 = 4'd15; a_sign2 = 4'd0; a_sign3 = 4'd9;
b_sign0 = 4'd16; b_sign1 = 4'd3; b_sign2 = 4'd15; b_sign3 = 4'd5;
@(posedge clk_i);
a_mant0 = 8'd155; a_mant1 = 8'd98; a_mant2 = 8'd159; a_mant3 = 8'd169;
b_mant0 = 8'd27; b_mant1 = 8'd163; b_mant2 = 8'd15; b_mant3 = 8'd90;
a_exp0 = 10'd654; a_exp1 = 10'd144; a_exp2 = 10'd612; a_exp3 = 10'd408;
b_exp0 = 10'd64; b_exp1 = 10'd411; b_exp2 = 10'd520; b_exp3 = 10'd379;
a_sign0 = 4'd2; a_sign1 = 4'd12; a_sign2 = 4'd12; a_sign3 = 4'd5;
b_sign0 = 4'd5; b_sign1 = 4'd11; b_sign2 = 4'd6; b_sign3 = 4'd1;
@(posedge clk_i);
a_mant0 = 8'd48; a_mant1 = 8'd32; a_mant2 = 8'd242; a_mant3 = 8'd1;
b_mant0 = 8'd114; b_mant1 = 8'd162; b_mant2 = 8'd218; b_mant3 = 8'd51;
a_exp0 = 10'd748; a_exp1 = 10'd202; a_exp2 = 10'd13; a_exp3 = 10'd175;
b_exp0 = 10'd548; b_exp1 = 10'd726; b_exp2 = 10'd164; b_exp3 = 10'd940;
a_sign0 = 4'd1; a_sign1 = 4'd3; a_sign2 = 4'd14; a_sign3 = 4'd13;
b_sign0 = 4'd6; b_sign1 = 4'd10; b_sign2 = 4'd8; b_sign3 = 4'd10;
@(posedge clk_i);
shared_exps0 = 8'd104;
shared_exps1 = 8'd131;
a_mant0 = 8'd153; a_mant1 = 8'd122; a_mant2 = 8'd98; a_mant3 = 8'd53;
b_mant0 = 8'd62; b_mant1 = 8'd18; b_mant2 = 8'd248; b_mant3 = 8'd181;
a_exp0 = 10'd144; a_exp1 = 10'd930; a_exp2 = 10'd496; a_exp3 = 10'd105;
b_exp0 = 10'd749; b_exp1 = 10'd922; b_exp2 = 10'd662; b_exp3 = 10'd786;
a_sign0 = 4'd9; a_sign1 = 4'd10; a_sign2 = 4'd4; a_sign3 = 4'd16;
b_sign0 = 4'd2; b_sign1 = 4'd13; b_sign2 = 4'd8; b_sign3 = 4'd14;
@(posedge clk_i);
a_mant0 = 8'd105; a_mant1 = 8'd99; a_mant2 = 8'd9; a_mant3 = 8'd68;
b_mant0 = 8'd184; b_mant1 = 8'd121; b_mant2 = 8'd129; b_mant3 = 8'd137;
a_exp0 = 10'd298; a_exp1 = 10'd602; a_exp2 = 10'd33; a_exp3 = 10'd196;
b_exp0 = 10'd880; b_exp1 = 10'd164; b_exp2 = 10'd48; b_exp3 = 10'd646;
a_sign0 = 4'd11; a_sign1 = 4'd15; a_sign2 = 4'd16; a_sign3 = 4'd7;
b_sign0 = 4'd16; b_sign1 = 4'd12; b_sign2 = 4'd15; b_sign3 = 4'd3;
@(posedge clk_i);
a_mant0 = 8'd90; a_mant1 = 8'd160; a_mant2 = 8'd211; a_mant3 = 8'd55;
b_mant0 = 8'd31; b_mant1 = 8'd120; b_mant2 = 8'd4; b_mant3 = 8'd156;
a_exp0 = 10'd359; a_exp1 = 10'd176; a_exp2 = 10'd1019; a_exp3 = 10'd358;
b_exp0 = 10'd790; b_exp1 = 10'd876; b_exp2 = 10'd664; b_exp3 = 10'd633;
a_sign0 = 4'd12; a_sign1 = 4'd8; a_sign2 = 4'd5; a_sign3 = 4'd8;
b_sign0 = 4'd7; b_sign1 = 4'd9; b_sign2 = 4'd15; b_sign3 = 4'd13;
@(posedge clk_i);
a_mant0 = 8'd253; a_mant1 = 8'd139; a_mant2 = 8'd166; a_mant3 = 8'd35;
b_mant0 = 8'd59; b_mant1 = 8'd98; b_mant2 = 8'd178; b_mant3 = 8'd25;
a_exp0 = 10'd618; a_exp1 = 10'd571; a_exp2 = 10'd216; a_exp3 = 10'd647;
b_exp0 = 10'd283; b_exp1 = 10'd582; b_exp2 = 10'd496; b_exp3 = 10'd467;
a_sign0 = 4'd0; a_sign1 = 4'd12; a_sign2 = 4'd4; a_sign3 = 4'd12;
b_sign0 = 4'd13; b_sign1 = 4'd11; b_sign2 = 4'd15; b_sign3 = 4'd14;
@(posedge clk_i);
a_mant0 = 8'd244; a_mant1 = 8'd217; a_mant2 = 8'd155; a_mant3 = 8'd6;
b_mant0 = 8'd29; b_mant1 = 8'd84; b_mant2 = 8'd250; b_mant3 = 8'd164;
a_exp0 = 10'd187; a_exp1 = 10'd1002; a_exp2 = 10'd761; a_exp3 = 10'd283;
b_exp0 = 10'd670; b_exp1 = 10'd858; b_exp2 = 10'd290; b_exp3 = 10'd289;
a_sign0 = 4'd7; a_sign1 = 4'd0; a_sign2 = 4'd5; a_sign3 = 4'd11;
b_sign0 = 4'd10; b_sign1 = 4'd10; b_sign2 = 4'd14; b_sign3 = 4'd7;
@(posedge clk_i);
a_mant0 = 8'd234; a_mant1 = 8'd231; a_mant2 = 8'd18; a_mant3 = 8'd245;
b_mant0 = 8'd120; b_mant1 = 8'd103; b_mant2 = 8'd190; b_mant3 = 8'd211;
a_exp0 = 10'd314; a_exp1 = 10'd283; a_exp2 = 10'd624; a_exp3 = 10'd305;
b_exp0 = 10'd188; b_exp1 = 10'd855; b_exp2 = 10'd206; b_exp3 = 10'd785;
a_sign0 = 4'd8; a_sign1 = 4'd13; a_sign2 = 4'd3; a_sign3 = 4'd2;
b_sign0 = 4'd3; b_sign1 = 4'd15; b_sign2 = 4'd14; b_sign3 = 4'd7;
@(posedge clk_i);
a_mant0 = 8'd169; a_mant1 = 8'd248; a_mant2 = 8'd200; a_mant3 = 8'd180;
b_mant0 = 8'd89; b_mant1 = 8'd234; b_mant2 = 8'd226; b_mant3 = 8'd42;
a_exp0 = 10'd85; a_exp1 = 10'd33; a_exp2 = 10'd243; a_exp3 = 10'd250;
b_exp0 = 10'd589; b_exp1 = 10'd192; b_exp2 = 10'd477; b_exp3 = 10'd968;
a_sign0 = 4'd3; a_sign1 = 4'd3; a_sign2 = 4'd6; a_sign3 = 4'd9;
b_sign0 = 4'd13; b_sign1 = 4'd5; b_sign2 = 4'd4; b_sign3 = 4'd11;
@(posedge clk_i);
a_mant0 = 8'd29; a_mant1 = 8'd141; a_mant2 = 8'd137; a_mant3 = 8'd143;
b_mant0 = 8'd164; b_mant1 = 8'd221; b_mant2 = 8'd20; b_mant3 = 8'd177;
a_exp0 = 10'd838; a_exp1 = 10'd441; a_exp2 = 10'd771; a_exp3 = 10'd627;
b_exp0 = 10'd730; b_exp1 = 10'd432; b_exp2 = 10'd172; b_exp3 = 10'd93;
a_sign0 = 4'd4; a_sign1 = 4'd2; a_sign2 = 4'd15; a_sign3 = 4'd2;
b_sign0 = 4'd8; b_sign1 = 4'd0; b_sign2 = 4'd9; b_sign3 = 4'd3;
@(posedge clk_i);
shared_exps0 = 8'd127;
shared_exps1 = 8'd131;
a_mant0 = 8'd220; a_mant1 = 8'd43; a_mant2 = 8'd240; a_mant3 = 8'd124;
b_mant0 = 8'd87; b_mant1 = 8'd146; b_mant2 = 8'd73; b_mant3 = 8'd176;
a_exp0 = 10'd784; a_exp1 = 10'd353; a_exp2 = 10'd189; a_exp3 = 10'd787;
b_exp0 = 10'd292; b_exp1 = 10'd789; b_exp2 = 10'd700; b_exp3 = 10'd714;
a_sign0 = 4'd13; a_sign1 = 4'd15; a_sign2 = 4'd4; a_sign3 = 4'd15;
b_sign0 = 4'd10; b_sign1 = 4'd12; b_sign2 = 4'd0; b_sign3 = 4'd16;
@(posedge clk_i);
a_mant0 = 8'd19; a_mant1 = 8'd66; a_mant2 = 8'd71; a_mant3 = 8'd226;
b_mant0 = 8'd197; b_mant1 = 8'd102; b_mant2 = 8'd174; b_mant3 = 8'd190;
a_exp0 = 10'd645; a_exp1 = 10'd1005; a_exp2 = 10'd237; a_exp3 = 10'd928;
b_exp0 = 10'd914; b_exp1 = 10'd148; b_exp2 = 10'd986; b_exp3 = 10'd348;
a_sign0 = 4'd13; a_sign1 = 4'd9; a_sign2 = 4'd10; a_sign3 = 4'd4;
b_sign0 = 4'd7; b_sign1 = 4'd1; b_sign2 = 4'd9; b_sign3 = 4'd7;
@(posedge clk_i);
a_mant0 = 8'd113; a_mant1 = 8'd205; a_mant2 = 8'd167; a_mant3 = 8'd51;
b_mant0 = 8'd0; b_mant1 = 8'd240; b_mant2 = 8'd195; b_mant3 = 8'd254;
a_exp0 = 10'd699; a_exp1 = 10'd314; a_exp2 = 10'd57; a_exp3 = 10'd639;
b_exp0 = 10'd870; b_exp1 = 10'd268; b_exp2 = 10'd464; b_exp3 = 10'd44;
a_sign0 = 4'd10; a_sign1 = 4'd14; a_sign2 = 4'd16; a_sign3 = 4'd0;
b_sign0 = 4'd1; b_sign1 = 4'd9; b_sign2 = 4'd1; b_sign3 = 4'd4;
@(posedge clk_i);
a_mant0 = 8'd245; a_mant1 = 8'd128; a_mant2 = 8'd114; a_mant3 = 8'd11;
b_mant0 = 8'd106; b_mant1 = 8'd159; b_mant2 = 8'd171; b_mant3 = 8'd94;
a_exp0 = 10'd975; a_exp1 = 10'd185; a_exp2 = 10'd893; a_exp3 = 10'd544;
b_exp0 = 10'd382; b_exp1 = 10'd927; b_exp2 = 10'd635; b_exp3 = 10'd195;
a_sign0 = 4'd3; a_sign1 = 4'd7; a_sign2 = 4'd10; a_sign3 = 4'd2;
b_sign0 = 4'd9; b_sign1 = 4'd11; b_sign2 = 4'd8; b_sign3 = 4'd1;
@(posedge clk_i);
a_mant0 = 8'd213; a_mant1 = 8'd126; a_mant2 = 8'd107; a_mant3 = 8'd20;
b_mant0 = 8'd250; b_mant1 = 8'd235; b_mant2 = 8'd196; b_mant3 = 8'd103;
a_exp0 = 10'd740; a_exp1 = 10'd431; a_exp2 = 10'd591; a_exp3 = 10'd463;
b_exp0 = 10'd458; b_exp1 = 10'd689; b_exp2 = 10'd44; b_exp3 = 10'd898;
a_sign0 = 4'd8; a_sign1 = 4'd11; a_sign2 = 4'd1; a_sign3 = 4'd1;
b_sign0 = 4'd9; b_sign1 = 4'd15; b_sign2 = 4'd15; b_sign3 = 4'd1;
@(posedge clk_i);
a_mant0 = 8'd89; a_mant1 = 8'd24; a_mant2 = 8'd222; a_mant3 = 8'd175;
b_mant0 = 8'd1; b_mant1 = 8'd209; b_mant2 = 8'd177; b_mant3 = 8'd221;
a_exp0 = 10'd783; a_exp1 = 10'd309; a_exp2 = 10'd859; a_exp3 = 10'd676;
b_exp0 = 10'd589; b_exp1 = 10'd26; b_exp2 = 10'd196; b_exp3 = 10'd816;
a_sign0 = 4'd10; a_sign1 = 4'd6; a_sign2 = 4'd6; a_sign3 = 4'd2;
b_sign0 = 4'd1; b_sign1 = 4'd11; b_sign2 = 4'd3; b_sign3 = 4'd9;
@(posedge clk_i);
a_mant0 = 8'd30; a_mant1 = 8'd208; a_mant2 = 8'd214; a_mant3 = 8'd73;
b_mant0 = 8'd154; b_mant1 = 8'd20; b_mant2 = 8'd179; b_mant3 = 8'd130;
a_exp0 = 10'd896; a_exp1 = 10'd728; a_exp2 = 10'd681; a_exp3 = 10'd401;
b_exp0 = 10'd584; b_exp1 = 10'd219; b_exp2 = 10'd315; b_exp3 = 10'd616;
a_sign0 = 4'd7; a_sign1 = 4'd5; a_sign2 = 4'd4; a_sign3 = 4'd14;
b_sign0 = 4'd14; b_sign1 = 4'd11; b_sign2 = 4'd3; b_sign3 = 4'd9;
@(posedge clk_i);
a_mant0 = 8'd148; a_mant1 = 8'd181; a_mant2 = 8'd26; a_mant3 = 8'd111;
b_mant0 = 8'd146; b_mant1 = 8'd11; b_mant2 = 8'd248; b_mant3 = 8'd230;
a_exp0 = 10'd609; a_exp1 = 10'd74; a_exp2 = 10'd489; a_exp3 = 10'd200;
b_exp0 = 10'd456; b_exp1 = 10'd716; b_exp2 = 10'd489; b_exp3 = 10'd98;
a_sign0 = 4'd4; a_sign1 = 4'd6; a_sign2 = 4'd13; a_sign3 = 4'd13;
b_sign0 = 4'd13; b_sign1 = 4'd3; b_sign2 = 4'd4; b_sign3 = 4'd15;
@(posedge clk_i);
shared_exps0 = 8'd146;
shared_exps1 = 8'd121;
a_mant0 = 8'd31; a_mant1 = 8'd191; a_mant2 = 8'd153; a_mant3 = 8'd17;
b_mant0 = 8'd23; b_mant1 = 8'd20; b_mant2 = 8'd224; b_mant3 = 8'd190;
a_exp0 = 10'd700; a_exp1 = 10'd999; a_exp2 = 10'd30; a_exp3 = 10'd270;
b_exp0 = 10'd433; b_exp1 = 10'd639; b_exp2 = 10'd184; b_exp3 = 10'd548;
a_sign0 = 4'd0; a_sign1 = 4'd9; a_sign2 = 4'd7; a_sign3 = 4'd12;
b_sign0 = 4'd7; b_sign1 = 4'd11; b_sign2 = 4'd1; b_sign3 = 4'd11;
@(posedge clk_i);
a_mant0 = 8'd75; a_mant1 = 8'd192; a_mant2 = 8'd192; a_mant3 = 8'd186;
b_mant0 = 8'd151; b_mant1 = 8'd117; b_mant2 = 8'd31; b_mant3 = 8'd65;
a_exp0 = 10'd830; a_exp1 = 10'd724; a_exp2 = 10'd762; a_exp3 = 10'd766;
b_exp0 = 10'd973; b_exp1 = 10'd418; b_exp2 = 10'd10; b_exp3 = 10'd1018;
a_sign0 = 4'd16; a_sign1 = 4'd11; a_sign2 = 4'd0; a_sign3 = 4'd8;
b_sign0 = 4'd3; b_sign1 = 4'd8; b_sign2 = 4'd12; b_sign3 = 4'd14;
@(posedge clk_i);
a_mant0 = 8'd169; a_mant1 = 8'd132; a_mant2 = 8'd85; a_mant3 = 8'd176;
b_mant0 = 8'd162; b_mant1 = 8'd154; b_mant2 = 8'd138; b_mant3 = 8'd27;
a_exp0 = 10'd293; a_exp1 = 10'd918; a_exp2 = 10'd408; a_exp3 = 10'd300;
b_exp0 = 10'd922; b_exp1 = 10'd104; b_exp2 = 10'd13; b_exp3 = 10'd456;
a_sign0 = 4'd3; a_sign1 = 4'd12; a_sign2 = 4'd5; a_sign3 = 4'd9;
b_sign0 = 4'd13; b_sign1 = 4'd16; b_sign2 = 4'd11; b_sign3 = 4'd10;
@(posedge clk_i);
a_mant0 = 8'd22; a_mant1 = 8'd96; a_mant2 = 8'd250; a_mant3 = 8'd31;
b_mant0 = 8'd192; b_mant1 = 8'd249; b_mant2 = 8'd47; b_mant3 = 8'd208;
a_exp0 = 10'd577; a_exp1 = 10'd212; a_exp2 = 10'd68; a_exp3 = 10'd345;
b_exp0 = 10'd573; b_exp1 = 10'd510; b_exp2 = 10'd302; b_exp3 = 10'd585;
a_sign0 = 4'd6; a_sign1 = 4'd1; a_sign2 = 4'd2; a_sign3 = 4'd11;
b_sign0 = 4'd2; b_sign1 = 4'd4; b_sign2 = 4'd6; b_sign3 = 4'd10;
@(posedge clk_i);
a_mant0 = 8'd138; a_mant1 = 8'd157; a_mant2 = 8'd180; a_mant3 = 8'd92;
b_mant0 = 8'd8; b_mant1 = 8'd2; b_mant2 = 8'd230; b_mant3 = 8'd148;
a_exp0 = 10'd119; a_exp1 = 10'd657; a_exp2 = 10'd37; a_exp3 = 10'd841;
b_exp0 = 10'd545; b_exp1 = 10'd536; b_exp2 = 10'd1001; b_exp3 = 10'd759;
a_sign0 = 4'd11; a_sign1 = 4'd13; a_sign2 = 4'd7; a_sign3 = 4'd14;
b_sign0 = 4'd5; b_sign1 = 4'd9; b_sign2 = 4'd8; b_sign3 = 4'd1;
@(posedge clk_i);
a_mant0 = 8'd110; a_mant1 = 8'd239; a_mant2 = 8'd11; a_mant3 = 8'd54;
b_mant0 = 8'd121; b_mant1 = 8'd149; b_mant2 = 8'd101; b_mant3 = 8'd68;
a_exp0 = 10'd103; a_exp1 = 10'd72; a_exp2 = 10'd614; a_exp3 = 10'd76;
b_exp0 = 10'd404; b_exp1 = 10'd648; b_exp2 = 10'd691; b_exp3 = 10'd87;
a_sign0 = 4'd16; a_sign1 = 4'd10; a_sign2 = 4'd14; a_sign3 = 4'd16;
b_sign0 = 4'd15; b_sign1 = 4'd4; b_sign2 = 4'd9; b_sign3 = 4'd9;
@(posedge clk_i);
a_mant0 = 8'd0; a_mant1 = 8'd196; a_mant2 = 8'd105; a_mant3 = 8'd121;
b_mant0 = 8'd203; b_mant1 = 8'd160; b_mant2 = 8'd205; b_mant3 = 8'd128;
a_exp0 = 10'd491; a_exp1 = 10'd177; a_exp2 = 10'd552; a_exp3 = 10'd792;
b_exp0 = 10'd597; b_exp1 = 10'd736; b_exp2 = 10'd217; b_exp3 = 10'd328;
a_sign0 = 4'd9; a_sign1 = 4'd1; a_sign2 = 4'd2; a_sign3 = 4'd16;
b_sign0 = 4'd15; b_sign1 = 4'd4; b_sign2 = 4'd5; b_sign3 = 4'd10;
@(posedge clk_i);
a_mant0 = 8'd232; a_mant1 = 8'd142; a_mant2 = 8'd61; a_mant3 = 8'd104;
b_mant0 = 8'd160; b_mant1 = 8'd90; b_mant2 = 8'd70; b_mant3 = 8'd121;
a_exp0 = 10'd656; a_exp1 = 10'd898; a_exp2 = 10'd70; a_exp3 = 10'd664;
b_exp0 = 10'd174; b_exp1 = 10'd45; b_exp2 = 10'd392; b_exp3 = 10'd301;
a_sign0 = 4'd10; a_sign1 = 4'd14; a_sign2 = 4'd13; a_sign3 = 4'd1;
b_sign0 = 4'd14; b_sign1 = 4'd12; b_sign2 = 4'd6; b_sign3 = 4'd9;
@(posedge clk_i);
shared_exps0 = 8'd110;
shared_exps1 = 8'd79;
rstn = 0;
@(posedge clk_i);
rstn = 1;
a_mant0 = 8'd245; a_mant1 = 8'd80; a_mant2 = 8'd173; a_mant3 = 8'd103;
b_mant0 = 8'd38; b_mant1 = 8'd118; b_mant2 = 8'd138; b_mant3 = 8'd67;
a_exp0 = 10'd121; a_exp1 = 10'd651; a_exp2 = 10'd821; a_exp3 = 10'd535;
b_exp0 = 10'd687; b_exp1 = 10'd570; b_exp2 = 10'd495; b_exp3 = 10'd326;
a_sign0 = 4'd4; a_sign1 = 4'd2; a_sign2 = 4'd3; a_sign3 = 4'd3;
b_sign0 = 4'd5; b_sign1 = 4'd12; b_sign2 = 4'd8; b_sign3 = 4'd13;
@(posedge clk_i);
a_mant0 = 8'd73; a_mant1 = 8'd155; a_mant2 = 8'd148; a_mant3 = 8'd131;
b_mant0 = 8'd21; b_mant1 = 8'd139; b_mant2 = 8'd106; b_mant3 = 8'd119;
a_exp0 = 10'd758; a_exp1 = 10'd409; a_exp2 = 10'd506; a_exp3 = 10'd90;
b_exp0 = 10'd389; b_exp1 = 10'd687; b_exp2 = 10'd499; b_exp3 = 10'd530;
a_sign0 = 4'd15; a_sign1 = 4'd5; a_sign2 = 4'd5; a_sign3 = 4'd16;
b_sign0 = 4'd4; b_sign1 = 4'd4; b_sign2 = 4'd5; b_sign3 = 4'd2;
@(posedge clk_i);
a_mant0 = 8'd51; a_mant1 = 8'd227; a_mant2 = 8'd86; a_mant3 = 8'd236;
b_mant0 = 8'd199; b_mant1 = 8'd11; b_mant2 = 8'd207; b_mant3 = 8'd14;
a_exp0 = 10'd163; a_exp1 = 10'd583; a_exp2 = 10'd779; a_exp3 = 10'd876;
b_exp0 = 10'd224; b_exp1 = 10'd80; b_exp2 = 10'd469; b_exp3 = 10'd261;
a_sign0 = 4'd1; a_sign1 = 4'd5; a_sign2 = 4'd7; a_sign3 = 4'd13;
b_sign0 = 4'd12; b_sign1 = 4'd5; b_sign2 = 4'd3; b_sign3 = 4'd14;
@(posedge clk_i);
a_mant0 = 8'd251; a_mant1 = 8'd251; a_mant2 = 8'd137; a_mant3 = 8'd170;
b_mant0 = 8'd151; b_mant1 = 8'd106; b_mant2 = 8'd250; b_mant3 = 8'd18;
a_exp0 = 10'd434; a_exp1 = 10'd379; a_exp2 = 10'd953; a_exp3 = 10'd301;
b_exp0 = 10'd349; b_exp1 = 10'd285; b_exp2 = 10'd753; b_exp3 = 10'd929;
a_sign0 = 4'd0; a_sign1 = 4'd2; a_sign2 = 4'd13; a_sign3 = 4'd14;
b_sign0 = 4'd9; b_sign1 = 4'd13; b_sign2 = 4'd8; b_sign3 = 4'd10;
@(posedge clk_i);
a_mant0 = 8'd36; a_mant1 = 8'd191; a_mant2 = 8'd64; a_mant3 = 8'd18;
b_mant0 = 8'd112; b_mant1 = 8'd247; b_mant2 = 8'd251; b_mant3 = 8'd167;
a_exp0 = 10'd426; a_exp1 = 10'd521; a_exp2 = 10'd102; a_exp3 = 10'd312;
b_exp0 = 10'd744; b_exp1 = 10'd652; b_exp2 = 10'd179; b_exp3 = 10'd539;
a_sign0 = 4'd1; a_sign1 = 4'd13; a_sign2 = 4'd11; a_sign3 = 4'd12;
b_sign0 = 4'd9; b_sign1 = 4'd14; b_sign2 = 4'd12; b_sign3 = 4'd4;
@(posedge clk_i);
a_mant0 = 8'd122; a_mant1 = 8'd48; a_mant2 = 8'd117; a_mant3 = 8'd126;
b_mant0 = 8'd111; b_mant1 = 8'd33; b_mant2 = 8'd178; b_mant3 = 8'd204;
a_exp0 = 10'd800; a_exp1 = 10'd197; a_exp2 = 10'd388; a_exp3 = 10'd487;
b_exp0 = 10'd104; b_exp1 = 10'd975; b_exp2 = 10'd887; b_exp3 = 10'd620;
a_sign0 = 4'd15; a_sign1 = 4'd7; a_sign2 = 4'd7; a_sign3 = 4'd2;
b_sign0 = 4'd5; b_sign1 = 4'd1; b_sign2 = 4'd16; b_sign3 = 4'd1;
@(posedge clk_i);
a_mant0 = 8'd58; a_mant1 = 8'd192; a_mant2 = 8'd191; a_mant3 = 8'd228;
b_mant0 = 8'd113; b_mant1 = 8'd190; b_mant2 = 8'd239; b_mant3 = 8'd128;
a_exp0 = 10'd20; a_exp1 = 10'd143; a_exp2 = 10'd438; a_exp3 = 10'd530;
b_exp0 = 10'd132; b_exp1 = 10'd674; b_exp2 = 10'd907; b_exp3 = 10'd301;
a_sign0 = 4'd8; a_sign1 = 4'd13; a_sign2 = 4'd9; a_sign3 = 4'd16;
b_sign0 = 4'd6; b_sign1 = 4'd13; b_sign2 = 4'd0; b_sign3 = 4'd7;
@(posedge clk_i);
shared_exps0 = 8'd128;
shared_exps1 = 8'd126;
a_mant0 = 8'd157; a_mant1 = 8'd75; a_mant2 = 8'd121; a_mant3 = 8'd86;
b_mant0 = 8'd4; b_mant1 = 8'd183; b_mant2 = 8'd77; b_mant3 = 8'd173;
a_exp0 = 10'd760; a_exp1 = 10'd242; a_exp2 = 10'd37; a_exp3 = 10'd1012;
b_exp0 = 10'd168; b_exp1 = 10'd765; b_exp2 = 10'd133; b_exp3 = 10'd965;
a_sign0 = 4'd4; a_sign1 = 4'd7; a_sign2 = 4'd4; a_sign3 = 4'd2;
b_sign0 = 4'd2; b_sign1 = 4'd6; b_sign2 = 4'd7; b_sign3 = 4'd3;
@(posedge clk_i);
a_mant0 = 8'd251; a_mant1 = 8'd144; a_mant2 = 8'd210; a_mant3 = 8'd194;
b_mant0 = 8'd74; b_mant1 = 8'd104; b_mant2 = 8'd51; b_mant3 = 8'd243;
a_exp0 = 10'd668; a_exp1 = 10'd193; a_exp2 = 10'd179; a_exp3 = 10'd579;
b_exp0 = 10'd898; b_exp1 = 10'd969; b_exp2 = 10'd150; b_exp3 = 10'd20;
a_sign0 = 4'd7; a_sign1 = 4'd1; a_sign2 = 4'd5; a_sign3 = 4'd4;
b_sign0 = 4'd2; b_sign1 = 4'd0; b_sign2 = 4'd1; b_sign3 = 4'd4;
@(posedge clk_i);
a_mant0 = 8'd223; a_mant1 = 8'd151; a_mant2 = 8'd131; a_mant3 = 8'd43;
b_mant0 = 8'd101; b_mant1 = 8'd14; b_mant2 = 8'd127; b_mant3 = 8'd180;
a_exp0 = 10'd234; a_exp1 = 10'd515; a_exp2 = 10'd276; a_exp3 = 10'd142;
b_exp0 = 10'd43; b_exp1 = 10'd417; b_exp2 = 10'd940; b_exp3 = 10'd342;
a_sign0 = 4'd8; a_sign1 = 4'd11; a_sign2 = 4'd4; a_sign3 = 4'd11;
b_sign0 = 4'd2; b_sign1 = 4'd0; b_sign2 = 4'd14; b_sign3 = 4'd8;
@(posedge clk_i);
a_mant0 = 8'd236; a_mant1 = 8'd179; a_mant2 = 8'd193; a_mant3 = 8'd166;
b_mant0 = 8'd23; b_mant1 = 8'd101; b_mant2 = 8'd25; b_mant3 = 8'd120;
a_exp0 = 10'd196; a_exp1 = 10'd912; a_exp2 = 10'd262; a_exp3 = 10'd229;
b_exp0 = 10'd336; b_exp1 = 10'd259; b_exp2 = 10'd644; b_exp3 = 10'd515;
a_sign0 = 4'd16; a_sign1 = 4'd11; a_sign2 = 4'd6; a_sign3 = 4'd10;
b_sign0 = 4'd6; b_sign1 = 4'd7; b_sign2 = 4'd16; b_sign3 = 4'd0;
@(posedge clk_i);
a_mant0 = 8'd197; a_mant1 = 8'd196; a_mant2 = 8'd195; a_mant3 = 8'd17;
b_mant0 = 8'd208; b_mant1 = 8'd194; b_mant2 = 8'd91; b_mant3 = 8'd225;
a_exp0 = 10'd631; a_exp1 = 10'd348; a_exp2 = 10'd41; a_exp3 = 10'd313;
b_exp0 = 10'd31; b_exp1 = 10'd123; b_exp2 = 10'd73; b_exp3 = 10'd479;
a_sign0 = 4'd1; a_sign1 = 4'd6; a_sign2 = 4'd11; a_sign3 = 4'd6;
b_sign0 = 4'd3; b_sign1 = 4'd10; b_sign2 = 4'd6; b_sign3 = 4'd8;
@(posedge clk_i);
a_mant0 = 8'd185; a_mant1 = 8'd147; a_mant2 = 8'd199; a_mant3 = 8'd98;
b_mant0 = 8'd142; b_mant1 = 8'd146; b_mant2 = 8'd119; b_mant3 = 8'd119;
a_exp0 = 10'd302; a_exp1 = 10'd728; a_exp2 = 10'd495; a_exp3 = 10'd927;
b_exp0 = 10'd457; b_exp1 = 10'd278; b_exp2 = 10'd142; b_exp3 = 10'd395;
a_sign0 = 4'd15; a_sign1 = 4'd13; a_sign2 = 4'd1; a_sign3 = 4'd9;
b_sign0 = 4'd12; b_sign1 = 4'd10; b_sign2 = 4'd7; b_sign3 = 4'd5;
@(posedge clk_i);
a_mant0 = 8'd196; a_mant1 = 8'd149; a_mant2 = 8'd45; a_mant3 = 8'd114;
b_mant0 = 8'd21; b_mant1 = 8'd86; b_mant2 = 8'd249; b_mant3 = 8'd47;
a_exp0 = 10'd435; a_exp1 = 10'd743; a_exp2 = 10'd401; a_exp3 = 10'd856;
b_exp0 = 10'd950; b_exp1 = 10'd202; b_exp2 = 10'd223; b_exp3 = 10'd280;
a_sign0 = 4'd10; a_sign1 = 4'd0; a_sign2 = 4'd5; a_sign3 = 4'd3;
b_sign0 = 4'd7; b_sign1 = 4'd2; b_sign2 = 4'd6; b_sign3 = 4'd4;
@(posedge clk_i);
a_mant0 = 8'd59; a_mant1 = 8'd48; a_mant2 = 8'd64; a_mant3 = 8'd254;
b_mant0 = 8'd137; b_mant1 = 8'd26; b_mant2 = 8'd202; b_mant3 = 8'd132;
a_exp0 = 10'd134; a_exp1 = 10'd176; a_exp2 = 10'd427; a_exp3 = 10'd422;
b_exp0 = 10'd409; b_exp1 = 10'd631; b_exp2 = 10'd340; b_exp3 = 10'd29;
a_sign0 = 4'd14; a_sign1 = 4'd16; a_sign2 = 4'd8; a_sign3 = 4'd10;
b_sign0 = 4'd8; b_sign1 = 4'd3; b_sign2 = 4'd8; b_sign3 = 4'd5;
@(posedge clk_i);
shared_exps0 = 8'd115;
shared_exps1 = 8'd113;
a_mant0 = 8'd116; a_mant1 = 8'd111; a_mant2 = 8'd4; a_mant3 = 8'd18;
b_mant0 = 8'd202; b_mant1 = 8'd213; b_mant2 = 8'd192; b_mant3 = 8'd99;
a_exp0 = 10'd1008; a_exp1 = 10'd371; a_exp2 = 10'd772; a_exp3 = 10'd311;
b_exp0 = 10'd412; b_exp1 = 10'd565; b_exp2 = 10'd415; b_exp3 = 10'd992;
a_sign0 = 4'd9; a_sign1 = 4'd5; a_sign2 = 4'd5; a_sign3 = 4'd0;
b_sign0 = 4'd2; b_sign1 = 4'd10; b_sign2 = 4'd3; b_sign3 = 4'd14;
@(posedge clk_i);
a_mant0 = 8'd147; a_mant1 = 8'd127; a_mant2 = 8'd195; a_mant3 = 8'd82;
b_mant0 = 8'd199; b_mant1 = 8'd19; b_mant2 = 8'd245; b_mant3 = 8'd34;
a_exp0 = 10'd84; a_exp1 = 10'd628; a_exp2 = 10'd791; a_exp3 = 10'd186;
b_exp0 = 10'd356; b_exp1 = 10'd819; b_exp2 = 10'd308; b_exp3 = 10'd20;
a_sign0 = 4'd5; a_sign1 = 4'd8; a_sign2 = 4'd15; a_sign3 = 4'd14;
b_sign0 = 4'd1; b_sign1 = 4'd16; b_sign2 = 4'd15; b_sign3 = 4'd14;
@(posedge clk_i);
a_mant0 = 8'd127; a_mant1 = 8'd233; a_mant2 = 8'd246; a_mant3 = 8'd197;
b_mant0 = 8'd221; b_mant1 = 8'd149; b_mant2 = 8'd107; b_mant3 = 8'd87;
a_exp0 = 10'd465; a_exp1 = 10'd138; a_exp2 = 10'd749; a_exp3 = 10'd824;
b_exp0 = 10'd285; b_exp1 = 10'd162; b_exp2 = 10'd617; b_exp3 = 10'd835;
a_sign0 = 4'd11; a_sign1 = 4'd1; a_sign2 = 4'd3; a_sign3 = 4'd8;
b_sign0 = 4'd16; b_sign1 = 4'd3; b_sign2 = 4'd13; b_sign3 = 4'd1;
@(posedge clk_i);
a_mant0 = 8'd172; a_mant1 = 8'd187; a_mant2 = 8'd243; a_mant3 = 8'd213;
b_mant0 = 8'd29; b_mant1 = 8'd61; b_mant2 = 8'd178; b_mant3 = 8'd209;
a_exp0 = 10'd199; a_exp1 = 10'd897; a_exp2 = 10'd264; a_exp3 = 10'd666;
b_exp0 = 10'd120; b_exp1 = 10'd326; b_exp2 = 10'd496; b_exp3 = 10'd65;
a_sign0 = 4'd0; a_sign1 = 4'd12; a_sign2 = 4'd9; a_sign3 = 4'd11;
b_sign0 = 4'd15; b_sign1 = 4'd6; b_sign2 = 4'd12; b_sign3 = 4'd12;
@(posedge clk_i);
a_mant0 = 8'd232; a_mant1 = 8'd88; a_mant2 = 8'd161; a_mant3 = 8'd185;
b_mant0 = 8'd173; b_mant1 = 8'd74; b_mant2 = 8'd98; b_mant3 = 8'd246;
a_exp0 = 10'd930; a_exp1 = 10'd117; a_exp2 = 10'd818; a_exp3 = 10'd586;
b_exp0 = 10'd80; b_exp1 = 10'd362; b_exp2 = 10'd63; b_exp3 = 10'd370;
a_sign0 = 4'd3; a_sign1 = 4'd12; a_sign2 = 4'd15; a_sign3 = 4'd2;
b_sign0 = 4'd0; b_sign1 = 4'd3; b_sign2 = 4'd3; b_sign3 = 4'd16;
@(posedge clk_i);
a_mant0 = 8'd199; a_mant1 = 8'd111; a_mant2 = 8'd118; a_mant3 = 8'd31;
b_mant0 = 8'd100; b_mant1 = 8'd177; b_mant2 = 8'd170; b_mant3 = 8'd170;
a_exp0 = 10'd246; a_exp1 = 10'd50; a_exp2 = 10'd528; a_exp3 = 10'd176;
b_exp0 = 10'd664; b_exp1 = 10'd199; b_exp2 = 10'd980; b_exp3 = 10'd560;
a_sign0 = 4'd12; a_sign1 = 4'd3; a_sign2 = 4'd6; a_sign3 = 4'd5;
b_sign0 = 4'd0; b_sign1 = 4'd1; b_sign2 = 4'd16; b_sign3 = 4'd8;
@(posedge clk_i);
a_mant0 = 8'd205; a_mant1 = 8'd211; a_mant2 = 8'd197; a_mant3 = 8'd26;
b_mant0 = 8'd234; b_mant1 = 8'd220; b_mant2 = 8'd103; b_mant3 = 8'd26;
a_exp0 = 10'd879; a_exp1 = 10'd213; a_exp2 = 10'd554; a_exp3 = 10'd489;
b_exp0 = 10'd973; b_exp1 = 10'd84; b_exp2 = 10'd632; b_exp3 = 10'd694;
a_sign0 = 4'd6; a_sign1 = 4'd3; a_sign2 = 4'd14; a_sign3 = 4'd8;
b_sign0 = 4'd14; b_sign1 = 4'd16; b_sign2 = 4'd6; b_sign3 = 4'd6;
@(posedge clk_i);
a_mant0 = 8'd168; a_mant1 = 8'd136; a_mant2 = 8'd222; a_mant3 = 8'd67;
b_mant0 = 8'd97; b_mant1 = 8'd155; b_mant2 = 8'd234; b_mant3 = 8'd171;
a_exp0 = 10'd1009; a_exp1 = 10'd4; a_exp2 = 10'd501; a_exp3 = 10'd858;
b_exp0 = 10'd21; b_exp1 = 10'd134; b_exp2 = 10'd67; b_exp3 = 10'd204;
a_sign0 = 4'd14; a_sign1 = 4'd3; a_sign2 = 4'd9; a_sign3 = 4'd2;
b_sign0 = 4'd15; b_sign1 = 4'd13; b_sign2 = 4'd7; b_sign3 = 4'd2;
@(posedge clk_i);
shared_exps0 = 8'd115;
shared_exps1 = 8'd163;
a_mant0 = 8'd46; a_mant1 = 8'd207; a_mant2 = 8'd129; a_mant3 = 8'd84;
b_mant0 = 8'd203; b_mant1 = 8'd51; b_mant2 = 8'd89; b_mant3 = 8'd250;
a_exp0 = 10'd329; a_exp1 = 10'd374; a_exp2 = 10'd423; a_exp3 = 10'd860;
b_exp0 = 10'd394; b_exp1 = 10'd342; b_exp2 = 10'd986; b_exp3 = 10'd655;
a_sign0 = 4'd7; a_sign1 = 4'd7; a_sign2 = 4'd5; a_sign3 = 4'd5;
b_sign0 = 4'd16; b_sign1 = 4'd5; b_sign2 = 4'd10; b_sign3 = 4'd5;
@(posedge clk_i);
a_mant0 = 8'd0; a_mant1 = 8'd73; a_mant2 = 8'd190; a_mant3 = 8'd26;
b_mant0 = 8'd76; b_mant1 = 8'd182; b_mant2 = 8'd62; b_mant3 = 8'd103;
a_exp0 = 10'd757; a_exp1 = 10'd81; a_exp2 = 10'd408; a_exp3 = 10'd308;
b_exp0 = 10'd465; b_exp1 = 10'd467; b_exp2 = 10'd229; b_exp3 = 10'd1008;
a_sign0 = 4'd13; a_sign1 = 4'd5; a_sign2 = 4'd1; a_sign3 = 4'd1;
b_sign0 = 4'd6; b_sign1 = 4'd15; b_sign2 = 4'd12; b_sign3 = 4'd14;
@(posedge clk_i);
a_mant0 = 8'd31; a_mant1 = 8'd255; a_mant2 = 8'd28; a_mant3 = 8'd111;
b_mant0 = 8'd16; b_mant1 = 8'd225; b_mant2 = 8'd127; b_mant3 = 8'd104;
a_exp0 = 10'd766; a_exp1 = 10'd700; a_exp2 = 10'd573; a_exp3 = 10'd556;
b_exp0 = 10'd188; b_exp1 = 10'd660; b_exp2 = 10'd167; b_exp3 = 10'd701;
a_sign0 = 4'd15; a_sign1 = 4'd1; a_sign2 = 4'd7; a_sign3 = 4'd15;
b_sign0 = 4'd15; b_sign1 = 4'd6; b_sign2 = 4'd4; b_sign3 = 4'd9;
@(posedge clk_i);
a_mant0 = 8'd207; a_mant1 = 8'd240; a_mant2 = 8'd168; a_mant3 = 8'd34;
b_mant0 = 8'd210; b_mant1 = 8'd194; b_mant2 = 8'd122; b_mant3 = 8'd212;
a_exp0 = 10'd411; a_exp1 = 10'd241; a_exp2 = 10'd829; a_exp3 = 10'd648;
b_exp0 = 10'd842; b_exp1 = 10'd312; b_exp2 = 10'd751; b_exp3 = 10'd8;
a_sign0 = 4'd14; a_sign1 = 4'd12; a_sign2 = 4'd14; a_sign3 = 4'd1;
b_sign0 = 4'd9; b_sign1 = 4'd2; b_sign2 = 4'd14; b_sign3 = 4'd11;
@(posedge clk_i);
a_mant0 = 8'd201; a_mant1 = 8'd8; a_mant2 = 8'd195; a_mant3 = 8'd236;
b_mant0 = 8'd218; b_mant1 = 8'd63; b_mant2 = 8'd56; b_mant3 = 8'd88;
a_exp0 = 10'd310; a_exp1 = 10'd312; a_exp2 = 10'd36; a_exp3 = 10'd2;
b_exp0 = 10'd710; b_exp1 = 10'd928; b_exp2 = 10'd442; b_exp3 = 10'd745;
a_sign0 = 4'd14; a_sign1 = 4'd12; a_sign2 = 4'd3; a_sign3 = 4'd4;
b_sign0 = 4'd8; b_sign1 = 4'd9; b_sign2 = 4'd13; b_sign3 = 4'd12;
@(posedge clk_i);
a_mant0 = 8'd205; a_mant1 = 8'd194; a_mant2 = 8'd89; a_mant3 = 8'd110;
b_mant0 = 8'd234; b_mant1 = 8'd248; b_mant2 = 8'd135; b_mant3 = 8'd122;
a_exp0 = 10'd183; a_exp1 = 10'd990; a_exp2 = 10'd760; a_exp3 = 10'd254;
b_exp0 = 10'd727; b_exp1 = 10'd407; b_exp2 = 10'd750; b_exp3 = 10'd742;
a_sign0 = 4'd11; a_sign1 = 4'd14; a_sign2 = 4'd6; a_sign3 = 4'd15;
b_sign0 = 4'd9; b_sign1 = 4'd0; b_sign2 = 4'd16; b_sign3 = 4'd0;
@(posedge clk_i);
a_mant0 = 8'd217; a_mant1 = 8'd153; a_mant2 = 8'd212; a_mant3 = 8'd29;
b_mant0 = 8'd246; b_mant1 = 8'd182; b_mant2 = 8'd176; b_mant3 = 8'd8;
a_exp0 = 10'd195; a_exp1 = 10'd695; a_exp2 = 10'd944; a_exp3 = 10'd766;
b_exp0 = 10'd1023; b_exp1 = 10'd87; b_exp2 = 10'd780; b_exp3 = 10'd334;
a_sign0 = 4'd2; a_sign1 = 4'd13; a_sign2 = 4'd11; a_sign3 = 4'd16;
b_sign0 = 4'd1; b_sign1 = 4'd4; b_sign2 = 4'd12; b_sign3 = 4'd4;
@(posedge clk_i);
a_mant0 = 8'd227; a_mant1 = 8'd136; a_mant2 = 8'd61; a_mant3 = 8'd102;
b_mant0 = 8'd109; b_mant1 = 8'd104; b_mant2 = 8'd17; b_mant3 = 8'd162;
a_exp0 = 10'd914; a_exp1 = 10'd379; a_exp2 = 10'd30; a_exp3 = 10'd598;
b_exp0 = 10'd849; b_exp1 = 10'd231; b_exp2 = 10'd653; b_exp3 = 10'd366;
a_sign0 = 4'd8; a_sign1 = 4'd10; a_sign2 = 4'd4; a_sign3 = 4'd6;
b_sign0 = 4'd12; b_sign1 = 4'd1; b_sign2 = 4'd7; b_sign3 = 4'd3;
@(posedge clk_i);
shared_exps0 = 8'd140;
shared_exps1 = 8'd113;
rstn = 0;
@(posedge clk_i);
rstn = 1;
a_mant0 = 8'd254; a_mant1 = 8'd32; a_mant2 = 8'd184; a_mant3 = 8'd235;
b_mant0 = 8'd5; b_mant1 = 8'd245; b_mant2 = 8'd165; b_mant3 = 8'd65;
a_exp0 = 10'd395; a_exp1 = 10'd234; a_exp2 = 10'd242; a_exp3 = 10'd763;
b_exp0 = 10'd178; b_exp1 = 10'd322; b_exp2 = 10'd139; b_exp3 = 10'd507;
a_sign0 = 4'd5; a_sign1 = 4'd8; a_sign2 = 4'd2; a_sign3 = 4'd11;
b_sign0 = 4'd4; b_sign1 = 4'd7; b_sign2 = 4'd11; b_sign3 = 4'd5;
@(posedge clk_i);
a_mant0 = 8'd67; a_mant1 = 8'd224; a_mant2 = 8'd67; a_mant3 = 8'd83;
b_mant0 = 8'd39; b_mant1 = 8'd60; b_mant2 = 8'd89; b_mant3 = 8'd6;
a_exp0 = 10'd806; a_exp1 = 10'd720; a_exp2 = 10'd12; a_exp3 = 10'd204;
b_exp0 = 10'd177; b_exp1 = 10'd552; b_exp2 = 10'd300; b_exp3 = 10'd610;
a_sign0 = 4'd4; a_sign1 = 4'd10; a_sign2 = 4'd1; a_sign3 = 4'd4;
b_sign0 = 4'd16; b_sign1 = 4'd11; b_sign2 = 4'd1; b_sign3 = 4'd15;
@(posedge clk_i);
a_mant0 = 8'd72; a_mant1 = 8'd242; a_mant2 = 8'd232; a_mant3 = 8'd141;
b_mant0 = 8'd239; b_mant1 = 8'd169; b_mant2 = 8'd159; b_mant3 = 8'd150;
a_exp0 = 10'd885; a_exp1 = 10'd441; a_exp2 = 10'd57; a_exp3 = 10'd910;
b_exp0 = 10'd636; b_exp1 = 10'd395; b_exp2 = 10'd312; b_exp3 = 10'd365;
a_sign0 = 4'd9; a_sign1 = 4'd7; a_sign2 = 4'd6; a_sign3 = 4'd13;
b_sign0 = 4'd3; b_sign1 = 4'd9; b_sign2 = 4'd13; b_sign3 = 4'd10;
@(posedge clk_i);
a_mant0 = 8'd60; a_mant1 = 8'd143; a_mant2 = 8'd116; a_mant3 = 8'd146;
b_mant0 = 8'd211; b_mant1 = 8'd60; b_mant2 = 8'd178; b_mant3 = 8'd185;
a_exp0 = 10'd433; a_exp1 = 10'd660; a_exp2 = 10'd506; a_exp3 = 10'd176;
b_exp0 = 10'd714; b_exp1 = 10'd214; b_exp2 = 10'd62; b_exp3 = 10'd44;
a_sign0 = 4'd4; a_sign1 = 4'd13; a_sign2 = 4'd10; a_sign3 = 4'd15;
b_sign0 = 4'd16; b_sign1 = 4'd2; b_sign2 = 4'd12; b_sign3 = 4'd4;
@(posedge clk_i);
a_mant0 = 8'd175; a_mant1 = 8'd80; a_mant2 = 8'd68; a_mant3 = 8'd58;
b_mant0 = 8'd177; b_mant1 = 8'd94; b_mant2 = 8'd240; b_mant3 = 8'd7;
a_exp0 = 10'd110; a_exp1 = 10'd1015; a_exp2 = 10'd813; a_exp3 = 10'd869;
b_exp0 = 10'd54; b_exp1 = 10'd1002; b_exp2 = 10'd715; b_exp3 = 10'd469;
a_sign0 = 4'd14; a_sign1 = 4'd8; a_sign2 = 4'd5; a_sign3 = 4'd11;
b_sign0 = 4'd2; b_sign1 = 4'd1; b_sign2 = 4'd1; b_sign3 = 4'd7;
@(posedge clk_i);
a_mant0 = 8'd207; a_mant1 = 8'd154; a_mant2 = 8'd68; a_mant3 = 8'd235;
b_mant0 = 8'd85; b_mant1 = 8'd246; b_mant2 = 8'd185; b_mant3 = 8'd152;
a_exp0 = 10'd97; a_exp1 = 10'd1018; a_exp2 = 10'd322; a_exp3 = 10'd856;
b_exp0 = 10'd781; b_exp1 = 10'd417; b_exp2 = 10'd149; b_exp3 = 10'd131;
a_sign0 = 4'd4; a_sign1 = 4'd9; a_sign2 = 4'd16; a_sign3 = 4'd0;
b_sign0 = 4'd14; b_sign1 = 4'd7; b_sign2 = 4'd5; b_sign3 = 4'd14;
@(posedge clk_i);
a_mant0 = 8'd53; a_mant1 = 8'd112; a_mant2 = 8'd216; a_mant3 = 8'd147;
b_mant0 = 8'd227; b_mant1 = 8'd61; b_mant2 = 8'd233; b_mant3 = 8'd200;
a_exp0 = 10'd832; a_exp1 = 10'd45; a_exp2 = 10'd672; a_exp3 = 10'd245;
b_exp0 = 10'd830; b_exp1 = 10'd831; b_exp2 = 10'd593; b_exp3 = 10'd667;
a_sign0 = 4'd13; a_sign1 = 4'd4; a_sign2 = 4'd9; a_sign3 = 4'd0;
b_sign0 = 4'd3; b_sign1 = 4'd1; b_sign2 = 4'd1; b_sign3 = 4'd2;
@(posedge clk_i);
shared_exps0 = 8'd113;
shared_exps1 = 8'd139;
a_mant0 = 8'd60; a_mant1 = 8'd49; a_mant2 = 8'd213; a_mant3 = 8'd65;
b_mant0 = 8'd50; b_mant1 = 8'd199; b_mant2 = 8'd74; b_mant3 = 8'd95;
a_exp0 = 10'd619; a_exp1 = 10'd1011; a_exp2 = 10'd654; a_exp3 = 10'd759;
b_exp0 = 10'd188; b_exp1 = 10'd524; b_exp2 = 10'd298; b_exp3 = 10'd886;
a_sign0 = 4'd6; a_sign1 = 4'd6; a_sign2 = 4'd16; a_sign3 = 4'd5;
b_sign0 = 4'd14; b_sign1 = 4'd5; b_sign2 = 4'd9; b_sign3 = 4'd9;
@(posedge clk_i);
a_mant0 = 8'd189; a_mant1 = 8'd151; a_mant2 = 8'd129; a_mant3 = 8'd216;
b_mant0 = 8'd153; b_mant1 = 8'd205; b_mant2 = 8'd236; b_mant3 = 8'd223;
a_exp0 = 10'd369; a_exp1 = 10'd148; a_exp2 = 10'd983; a_exp3 = 10'd103;
b_exp0 = 10'd802; b_exp1 = 10'd82; b_exp2 = 10'd391; b_exp3 = 10'd804;
a_sign0 = 4'd1; a_sign1 = 4'd12; a_sign2 = 4'd2; a_sign3 = 4'd13;
b_sign0 = 4'd13; b_sign1 = 4'd9; b_sign2 = 4'd3; b_sign3 = 4'd15;
@(posedge clk_i);
a_mant0 = 8'd75; a_mant1 = 8'd219; a_mant2 = 8'd131; a_mant3 = 8'd150;
b_mant0 = 8'd204; b_mant1 = 8'd15; b_mant2 = 8'd208; b_mant3 = 8'd43;
a_exp0 = 10'd603; a_exp1 = 10'd86; a_exp2 = 10'd182; a_exp3 = 10'd850;
b_exp0 = 10'd648; b_exp1 = 10'd183; b_exp2 = 10'd968; b_exp3 = 10'd480;
a_sign0 = 4'd12; a_sign1 = 4'd3; a_sign2 = 4'd9; a_sign3 = 4'd2;
b_sign0 = 4'd12; b_sign1 = 4'd1; b_sign2 = 4'd3; b_sign3 = 4'd1;
@(posedge clk_i);
a_mant0 = 8'd19; a_mant1 = 8'd69; a_mant2 = 8'd232; a_mant3 = 8'd155;
b_mant0 = 8'd145; b_mant1 = 8'd167; b_mant2 = 8'd246; b_mant3 = 8'd203;
a_exp0 = 10'd512; a_exp1 = 10'd247; a_exp2 = 10'd557; a_exp3 = 10'd108;
b_exp0 = 10'd203; b_exp1 = 10'd915; b_exp2 = 10'd388; b_exp3 = 10'd985;
a_sign0 = 4'd1; a_sign1 = 4'd8; a_sign2 = 4'd16; a_sign3 = 4'd3;
b_sign0 = 4'd14; b_sign1 = 4'd11; b_sign2 = 4'd2; b_sign3 = 4'd4;
@(posedge clk_i);
a_mant0 = 8'd249; a_mant1 = 8'd103; a_mant2 = 8'd72; a_mant3 = 8'd158;
b_mant0 = 8'd64; b_mant1 = 8'd191; b_mant2 = 8'd43; b_mant3 = 8'd80;
a_exp0 = 10'd549; a_exp1 = 10'd968; a_exp2 = 10'd230; a_exp3 = 10'd472;
b_exp0 = 10'd522; b_exp1 = 10'd882; b_exp2 = 10'd957; b_exp3 = 10'd884;
a_sign0 = 4'd9; a_sign1 = 4'd15; a_sign2 = 4'd7; a_sign3 = 4'd12;
b_sign0 = 4'd15; b_sign1 = 4'd8; b_sign2 = 4'd10; b_sign3 = 4'd12;
@(posedge clk_i);
a_mant0 = 8'd165; a_mant1 = 8'd233; a_mant2 = 8'd34; a_mant3 = 8'd66;
b_mant0 = 8'd77; b_mant1 = 8'd91; b_mant2 = 8'd64; b_mant3 = 8'd142;
a_exp0 = 10'd736; a_exp1 = 10'd1006; a_exp2 = 10'd876; a_exp3 = 10'd666;
b_exp0 = 10'd957; b_exp1 = 10'd140; b_exp2 = 10'd668; b_exp3 = 10'd579;
a_sign0 = 4'd3; a_sign1 = 4'd3; a_sign2 = 4'd15; a_sign3 = 4'd9;
b_sign0 = 4'd14; b_sign1 = 4'd1; b_sign2 = 4'd8; b_sign3 = 4'd11;
@(posedge clk_i);
a_mant0 = 8'd147; a_mant1 = 8'd102; a_mant2 = 8'd113; a_mant3 = 8'd80;
b_mant0 = 8'd228; b_mant1 = 8'd253; b_mant2 = 8'd193; b_mant3 = 8'd105;
a_exp0 = 10'd776; a_exp1 = 10'd280; a_exp2 = 10'd105; a_exp3 = 10'd89;
b_exp0 = 10'd392; b_exp1 = 10'd611; b_exp2 = 10'd4; b_exp3 = 10'd45;
a_sign0 = 4'd3; a_sign1 = 4'd10; a_sign2 = 4'd16; a_sign3 = 4'd9;
b_sign0 = 4'd7; b_sign1 = 4'd13; b_sign2 = 4'd5; b_sign3 = 4'd8;
@(posedge clk_i);
a_mant0 = 8'd90; a_mant1 = 8'd114; a_mant2 = 8'd36; a_mant3 = 8'd234;
b_mant0 = 8'd177; b_mant1 = 8'd160; b_mant2 = 8'd77; b_mant3 = 8'd130;
a_exp0 = 10'd144; a_exp1 = 10'd1017; a_exp2 = 10'd761; a_exp3 = 10'd125;
b_exp0 = 10'd605; b_exp1 = 10'd803; b_exp2 = 10'd418; b_exp3 = 10'd178;
a_sign0 = 4'd8; a_sign1 = 4'd14; a_sign2 = 4'd12; a_sign3 = 4'd15;
b_sign0 = 4'd14; b_sign1 = 4'd11; b_sign2 = 4'd7; b_sign3 = 4'd8;
@(posedge clk_i);
shared_exps0 = 8'd135;
shared_exps1 = 8'd132;
a_mant0 = 8'd91; a_mant1 = 8'd57; a_mant2 = 8'd15; a_mant3 = 8'd56;
b_mant0 = 8'd34; b_mant1 = 8'd201; b_mant2 = 8'd234; b_mant3 = 8'd6;
a_exp0 = 10'd861; a_exp1 = 10'd130; a_exp2 = 10'd29; a_exp3 = 10'd113;
b_exp0 = 10'd304; b_exp1 = 10'd264; b_exp2 = 10'd108; b_exp3 = 10'd636;
a_sign0 = 4'd3; a_sign1 = 4'd14; a_sign2 = 4'd11; a_sign3 = 4'd12;
b_sign0 = 4'd4; b_sign1 = 4'd11; b_sign2 = 4'd11; b_sign3 = 4'd3;
@(posedge clk_i);
a_mant0 = 8'd37; a_mant1 = 8'd171; a_mant2 = 8'd254; a_mant3 = 8'd14;
b_mant0 = 8'd32; b_mant1 = 8'd251; b_mant2 = 8'd122; b_mant3 = 8'd207;
a_exp0 = 10'd823; a_exp1 = 10'd22; a_exp2 = 10'd399; a_exp3 = 10'd125;
b_exp0 = 10'd897; b_exp1 = 10'd118; b_exp2 = 10'd187; b_exp3 = 10'd359;
a_sign0 = 4'd12; a_sign1 = 4'd16; a_sign2 = 4'd7; a_sign3 = 4'd12;
b_sign0 = 4'd12; b_sign1 = 4'd11; b_sign2 = 4'd14; b_sign3 = 4'd12;
@(posedge clk_i);
a_mant0 = 8'd121; a_mant1 = 8'd148; a_mant2 = 8'd9; a_mant3 = 8'd59;
b_mant0 = 8'd246; b_mant1 = 8'd66; b_mant2 = 8'd226; b_mant3 = 8'd84;
a_exp0 = 10'd378; a_exp1 = 10'd1009; a_exp2 = 10'd422; a_exp3 = 10'd80;
b_exp0 = 10'd195; b_exp1 = 10'd733; b_exp2 = 10'd804; b_exp3 = 10'd203;
a_sign0 = 4'd2; a_sign1 = 4'd9; a_sign2 = 4'd9; a_sign3 = 4'd0;
b_sign0 = 4'd13; b_sign1 = 4'd13; b_sign2 = 4'd11; b_sign3 = 4'd10;
@(posedge clk_i);
a_mant0 = 8'd129; a_mant1 = 8'd4; a_mant2 = 8'd30; a_mant3 = 8'd87;
b_mant0 = 8'd81; b_mant1 = 8'd157; b_mant2 = 8'd123; b_mant3 = 8'd119;
a_exp0 = 10'd888; a_exp1 = 10'd375; a_exp2 = 10'd641; a_exp3 = 10'd607;
b_exp0 = 10'd713; b_exp1 = 10'd924; b_exp2 = 10'd42; b_exp3 = 10'd42;
a_sign0 = 4'd16; a_sign1 = 4'd7; a_sign2 = 4'd15; a_sign3 = 4'd14;
b_sign0 = 4'd12; b_sign1 = 4'd5; b_sign2 = 4'd11; b_sign3 = 4'd4;
@(posedge clk_i);
a_mant0 = 8'd126; a_mant1 = 8'd220; a_mant2 = 8'd228; a_mant3 = 8'd32;
b_mant0 = 8'd236; b_mant1 = 8'd158; b_mant2 = 8'd251; b_mant3 = 8'd232;
a_exp0 = 10'd63; a_exp1 = 10'd848; a_exp2 = 10'd148; a_exp3 = 10'd883;
b_exp0 = 10'd692; b_exp1 = 10'd864; b_exp2 = 10'd673; b_exp3 = 10'd256;
a_sign0 = 4'd4; a_sign1 = 4'd9; a_sign2 = 4'd13; a_sign3 = 4'd8;
b_sign0 = 4'd6; b_sign1 = 4'd4; b_sign2 = 4'd2; b_sign3 = 4'd11;
@(posedge clk_i);
a_mant0 = 8'd135; a_mant1 = 8'd101; a_mant2 = 8'd122; a_mant3 = 8'd141;
b_mant0 = 8'd75; b_mant1 = 8'd151; b_mant2 = 8'd167; b_mant3 = 8'd194;
a_exp0 = 10'd967; a_exp1 = 10'd309; a_exp2 = 10'd1019; a_exp3 = 10'd528;
b_exp0 = 10'd821; b_exp1 = 10'd201; b_exp2 = 10'd242; b_exp3 = 10'd294;
a_sign0 = 4'd5; a_sign1 = 4'd14; a_sign2 = 4'd15; a_sign3 = 4'd16;
b_sign0 = 4'd6; b_sign1 = 4'd13; b_sign2 = 4'd15; b_sign3 = 4'd6;
@(posedge clk_i);
a_mant0 = 8'd53; a_mant1 = 8'd239; a_mant2 = 8'd68; a_mant3 = 8'd87;
b_mant0 = 8'd134; b_mant1 = 8'd187; b_mant2 = 8'd207; b_mant3 = 8'd230;
a_exp0 = 10'd48; a_exp1 = 10'd908; a_exp2 = 10'd925; a_exp3 = 10'd730;
b_exp0 = 10'd1000; b_exp1 = 10'd263; b_exp2 = 10'd87; b_exp3 = 10'd353;
a_sign0 = 4'd16; a_sign1 = 4'd10; a_sign2 = 4'd12; a_sign3 = 4'd11;
b_sign0 = 4'd1; b_sign1 = 4'd13; b_sign2 = 4'd13; b_sign3 = 4'd1;
@(posedge clk_i);
a_mant0 = 8'd201; a_mant1 = 8'd239; a_mant2 = 8'd216; a_mant3 = 8'd44;
b_mant0 = 8'd31; b_mant1 = 8'd20; b_mant2 = 8'd14; b_mant3 = 8'd117;
a_exp0 = 10'd633; a_exp1 = 10'd127; a_exp2 = 10'd542; a_exp3 = 10'd871;
b_exp0 = 10'd782; b_exp1 = 10'd744; b_exp2 = 10'd953; b_exp3 = 10'd179;
a_sign0 = 4'd1; a_sign1 = 4'd2; a_sign2 = 4'd4; a_sign3 = 4'd3;
b_sign0 = 4'd0; b_sign1 = 4'd16; b_sign2 = 4'd11; b_sign3 = 4'd9;
@(posedge clk_i);
shared_exps0 = 8'd138;
shared_exps1 = 8'd104;
a_mant0 = 8'd54; a_mant1 = 8'd126; a_mant2 = 8'd110; a_mant3 = 8'd215;
b_mant0 = 8'd93; b_mant1 = 8'd105; b_mant2 = 8'd131; b_mant3 = 8'd135;
a_exp0 = 10'd735; a_exp1 = 10'd118; a_exp2 = 10'd588; a_exp3 = 10'd464;
b_exp0 = 10'd986; b_exp1 = 10'd531; b_exp2 = 10'd623; b_exp3 = 10'd577;
a_sign0 = 4'd13; a_sign1 = 4'd11; a_sign2 = 4'd16; a_sign3 = 4'd0;
b_sign0 = 4'd11; b_sign1 = 4'd11; b_sign2 = 4'd2; b_sign3 = 4'd13;
@(posedge clk_i);
a_mant0 = 8'd138; a_mant1 = 8'd166; a_mant2 = 8'd54; a_mant3 = 8'd229;
b_mant0 = 8'd119; b_mant1 = 8'd183; b_mant2 = 8'd63; b_mant3 = 8'd57;
a_exp0 = 10'd930; a_exp1 = 10'd987; a_exp2 = 10'd135; a_exp3 = 10'd392;
b_exp0 = 10'd736; b_exp1 = 10'd861; b_exp2 = 10'd215; b_exp3 = 10'd391;
a_sign0 = 4'd1; a_sign1 = 4'd10; a_sign2 = 4'd10; a_sign3 = 4'd11;
b_sign0 = 4'd5; b_sign1 = 4'd6; b_sign2 = 4'd8; b_sign3 = 4'd13;
@(posedge clk_i);
a_mant0 = 8'd77; a_mant1 = 8'd75; a_mant2 = 8'd227; a_mant3 = 8'd158;
b_mant0 = 8'd196; b_mant1 = 8'd3; b_mant2 = 8'd144; b_mant3 = 8'd43;
a_exp0 = 10'd214; a_exp1 = 10'd737; a_exp2 = 10'd477; a_exp3 = 10'd659;
b_exp0 = 10'd356; b_exp1 = 10'd590; b_exp2 = 10'd151; b_exp3 = 10'd555;
a_sign0 = 4'd7; a_sign1 = 4'd6; a_sign2 = 4'd2; a_sign3 = 4'd8;
b_sign0 = 4'd10; b_sign1 = 4'd3; b_sign2 = 4'd5; b_sign3 = 4'd12;
@(posedge clk_i);
a_mant0 = 8'd25; a_mant1 = 8'd27; a_mant2 = 8'd100; a_mant3 = 8'd31;
b_mant0 = 8'd159; b_mant1 = 8'd181; b_mant2 = 8'd112; b_mant3 = 8'd120;
a_exp0 = 10'd55; a_exp1 = 10'd876; a_exp2 = 10'd797; a_exp3 = 10'd296;
b_exp0 = 10'd170; b_exp1 = 10'd710; b_exp2 = 10'd557; b_exp3 = 10'd2;
a_sign0 = 4'd13; a_sign1 = 4'd10; a_sign2 = 4'd2; a_sign3 = 4'd10;
b_sign0 = 4'd16; b_sign1 = 4'd13; b_sign2 = 4'd15; b_sign3 = 4'd11;
@(posedge clk_i);
a_mant0 = 8'd152; a_mant1 = 8'd134; a_mant2 = 8'd153; a_mant3 = 8'd11;
b_mant0 = 8'd94; b_mant1 = 8'd41; b_mant2 = 8'd128; b_mant3 = 8'd148;
a_exp0 = 10'd829; a_exp1 = 10'd582; a_exp2 = 10'd923; a_exp3 = 10'd492;
b_exp0 = 10'd398; b_exp1 = 10'd318; b_exp2 = 10'd739; b_exp3 = 10'd683;
a_sign0 = 4'd3; a_sign1 = 4'd5; a_sign2 = 4'd12; a_sign3 = 4'd6;
b_sign0 = 4'd12; b_sign1 = 4'd5; b_sign2 = 4'd16; b_sign3 = 4'd8;
@(posedge clk_i);
a_mant0 = 8'd73; a_mant1 = 8'd201; a_mant2 = 8'd63; a_mant3 = 8'd24;
b_mant0 = 8'd228; b_mant1 = 8'd198; b_mant2 = 8'd126; b_mant3 = 8'd184;
a_exp0 = 10'd534; a_exp1 = 10'd502; a_exp2 = 10'd475; a_exp3 = 10'd747;
b_exp0 = 10'd553; b_exp1 = 10'd615; b_exp2 = 10'd821; b_exp3 = 10'd285;
a_sign0 = 4'd2; a_sign1 = 4'd9; a_sign2 = 4'd7; a_sign3 = 4'd15;
b_sign0 = 4'd9; b_sign1 = 4'd10; b_sign2 = 4'd2; b_sign3 = 4'd8;
@(posedge clk_i);
a_mant0 = 8'd180; a_mant1 = 8'd237; a_mant2 = 8'd44; a_mant3 = 8'd38;
b_mant0 = 8'd218; b_mant1 = 8'd171; b_mant2 = 8'd108; b_mant3 = 8'd185;
a_exp0 = 10'd329; a_exp1 = 10'd559; a_exp2 = 10'd1015; a_exp3 = 10'd679;
b_exp0 = 10'd909; b_exp1 = 10'd278; b_exp2 = 10'd64; b_exp3 = 10'd274;
a_sign0 = 4'd6; a_sign1 = 4'd12; a_sign2 = 4'd6; a_sign3 = 4'd7;
b_sign0 = 4'd0; b_sign1 = 4'd9; b_sign2 = 4'd14; b_sign3 = 4'd11;
@(posedge clk_i);
a_mant0 = 8'd119; a_mant1 = 8'd89; a_mant2 = 8'd248; a_mant3 = 8'd20;
b_mant0 = 8'd153; b_mant1 = 8'd79; b_mant2 = 8'd187; b_mant3 = 8'd12;
a_exp0 = 10'd770; a_exp1 = 10'd167; a_exp2 = 10'd634; a_exp3 = 10'd188;
b_exp0 = 10'd483; b_exp1 = 10'd196; b_exp2 = 10'd122; b_exp3 = 10'd825;
a_sign0 = 4'd16; a_sign1 = 4'd14; a_sign2 = 4'd12; a_sign3 = 4'd4;
b_sign0 = 4'd7; b_sign1 = 4'd11; b_sign2 = 4'd3; b_sign3 = 4'd5;
@(posedge clk_i);
shared_exps0 = 8'd102;
shared_exps1 = 8'd137;
rstn = 0;
@(posedge clk_i);
rstn = 1;
a_mant0 = 8'd195; a_mant1 = 8'd53; a_mant2 = 8'd192; a_mant3 = 8'd87;
b_mant0 = 8'd118; b_mant1 = 8'd17; b_mant2 = 8'd235; b_mant3 = 8'd161;
a_exp0 = 10'd67; a_exp1 = 10'd682; a_exp2 = 10'd264; a_exp3 = 10'd978;
b_exp0 = 10'd857; b_exp1 = 10'd585; b_exp2 = 10'd9; b_exp3 = 10'd957;
a_sign0 = 4'd11; a_sign1 = 4'd9; a_sign2 = 4'd10; a_sign3 = 4'd1;
b_sign0 = 4'd8; b_sign1 = 4'd16; b_sign2 = 4'd16; b_sign3 = 4'd13;
@(posedge clk_i);
a_mant0 = 8'd122; a_mant1 = 8'd202; a_mant2 = 8'd24; a_mant3 = 8'd76;
b_mant0 = 8'd56; b_mant1 = 8'd88; b_mant2 = 8'd129; b_mant3 = 8'd61;
a_exp0 = 10'd704; a_exp1 = 10'd554; a_exp2 = 10'd159; a_exp3 = 10'd192;
b_exp0 = 10'd976; b_exp1 = 10'd590; b_exp2 = 10'd606; b_exp3 = 10'd285;
a_sign0 = 4'd8; a_sign1 = 4'd1; a_sign2 = 4'd15; a_sign3 = 4'd12;
b_sign0 = 4'd10; b_sign1 = 4'd11; b_sign2 = 4'd5; b_sign3 = 4'd6;
@(posedge clk_i);
a_mant0 = 8'd20; a_mant1 = 8'd141; a_mant2 = 8'd147; a_mant3 = 8'd59;
b_mant0 = 8'd69; b_mant1 = 8'd105; b_mant2 = 8'd118; b_mant3 = 8'd153;
a_exp0 = 10'd881; a_exp1 = 10'd532; a_exp2 = 10'd505; a_exp3 = 10'd192;
b_exp0 = 10'd17; b_exp1 = 10'd73; b_exp2 = 10'd876; b_exp3 = 10'd242;
a_sign0 = 4'd8; a_sign1 = 4'd7; a_sign2 = 4'd10; a_sign3 = 4'd8;
b_sign0 = 4'd14; b_sign1 = 4'd13; b_sign2 = 4'd7; b_sign3 = 4'd6;
@(posedge clk_i);
a_mant0 = 8'd206; a_mant1 = 8'd253; a_mant2 = 8'd76; a_mant3 = 8'd145;
b_mant0 = 8'd142; b_mant1 = 8'd100; b_mant2 = 8'd6; b_mant3 = 8'd64;
a_exp0 = 10'd857; a_exp1 = 10'd403; a_exp2 = 10'd628; a_exp3 = 10'd878;
b_exp0 = 10'd98; b_exp1 = 10'd161; b_exp2 = 10'd301; b_exp3 = 10'd735;
a_sign0 = 4'd5; a_sign1 = 4'd5; a_sign2 = 4'd7; a_sign3 = 4'd2;
b_sign0 = 4'd8; b_sign1 = 4'd1; b_sign2 = 4'd16; b_sign3 = 4'd12;
@(posedge clk_i);
a_mant0 = 8'd36; a_mant1 = 8'd214; a_mant2 = 8'd48; a_mant3 = 8'd95;
b_mant0 = 8'd141; b_mant1 = 8'd233; b_mant2 = 8'd52; b_mant3 = 8'd14;
a_exp0 = 10'd91; a_exp1 = 10'd649; a_exp2 = 10'd207; a_exp3 = 10'd196;
b_exp0 = 10'd426; b_exp1 = 10'd994; b_exp2 = 10'd193; b_exp3 = 10'd47;
a_sign0 = 4'd1; a_sign1 = 4'd8; a_sign2 = 4'd8; a_sign3 = 4'd0;
b_sign0 = 4'd9; b_sign1 = 4'd3; b_sign2 = 4'd6; b_sign3 = 4'd12;
@(posedge clk_i);
a_mant0 = 8'd15; a_mant1 = 8'd250; a_mant2 = 8'd111; a_mant3 = 8'd111;
b_mant0 = 8'd124; b_mant1 = 8'd199; b_mant2 = 8'd43; b_mant3 = 8'd75;
a_exp0 = 10'd603; a_exp1 = 10'd146; a_exp2 = 10'd606; a_exp3 = 10'd900;
b_exp0 = 10'd961; b_exp1 = 10'd11; b_exp2 = 10'd780; b_exp3 = 10'd364;
a_sign0 = 4'd11; a_sign1 = 4'd8; a_sign2 = 4'd7; a_sign3 = 4'd6;
b_sign0 = 4'd8; b_sign1 = 4'd16; b_sign2 = 4'd5; b_sign3 = 4'd6;
@(posedge clk_i);
a_mant0 = 8'd53; a_mant1 = 8'd228; a_mant2 = 8'd140; a_mant3 = 8'd162;
b_mant0 = 8'd231; b_mant1 = 8'd194; b_mant2 = 8'd12; b_mant3 = 8'd8;
a_exp0 = 10'd395; a_exp1 = 10'd599; a_exp2 = 10'd590; a_exp3 = 10'd956;
b_exp0 = 10'd525; b_exp1 = 10'd35; b_exp2 = 10'd659; b_exp3 = 10'd12;
a_sign0 = 4'd4; a_sign1 = 4'd1; a_sign2 = 4'd3; a_sign3 = 4'd15;
b_sign0 = 4'd13; b_sign1 = 4'd11; b_sign2 = 4'd15; b_sign3 = 4'd7;
@(posedge clk_i);
shared_exps0 = 8'd148;
shared_exps1 = 8'd127;
a_mant0 = 8'd121; a_mant1 = 8'd49; a_mant2 = 8'd120; a_mant3 = 8'd114;
b_mant0 = 8'd31; b_mant1 = 8'd190; b_mant2 = 8'd196; b_mant3 = 8'd48;
a_exp0 = 10'd981; a_exp1 = 10'd751; a_exp2 = 10'd419; a_exp3 = 10'd171;
b_exp0 = 10'd793; b_exp1 = 10'd312; b_exp2 = 10'd789; b_exp3 = 10'd912;
a_sign0 = 4'd9; a_sign1 = 4'd7; a_sign2 = 4'd7; a_sign3 = 4'd2;
b_sign0 = 4'd8; b_sign1 = 4'd3; b_sign2 = 4'd1; b_sign3 = 4'd9;
@(posedge clk_i);
a_mant0 = 8'd13; a_mant1 = 8'd36; a_mant2 = 8'd169; a_mant3 = 8'd101;
b_mant0 = 8'd43; b_mant1 = 8'd39; b_mant2 = 8'd31; b_mant3 = 8'd18;
a_exp0 = 10'd714; a_exp1 = 10'd854; a_exp2 = 10'd330; a_exp3 = 10'd595;
b_exp0 = 10'd789; b_exp1 = 10'd742; b_exp2 = 10'd305; b_exp3 = 10'd784;
a_sign0 = 4'd2; a_sign1 = 4'd9; a_sign2 = 4'd15; a_sign3 = 4'd6;
b_sign0 = 4'd11; b_sign1 = 4'd2; b_sign2 = 4'd8; b_sign3 = 4'd1;
@(posedge clk_i);
a_mant0 = 8'd123; a_mant1 = 8'd34; a_mant2 = 8'd70; a_mant3 = 8'd254;
b_mant0 = 8'd66; b_mant1 = 8'd255; b_mant2 = 8'd198; b_mant3 = 8'd168;
a_exp0 = 10'd722; a_exp1 = 10'd439; a_exp2 = 10'd165; a_exp3 = 10'd567;
b_exp0 = 10'd880; b_exp1 = 10'd304; b_exp2 = 10'd412; b_exp3 = 10'd698;
a_sign0 = 4'd13; a_sign1 = 4'd14; a_sign2 = 4'd2; a_sign3 = 4'd13;
b_sign0 = 4'd2; b_sign1 = 4'd16; b_sign2 = 4'd12; b_sign3 = 4'd16;
@(posedge clk_i);
a_mant0 = 8'd255; a_mant1 = 8'd38; a_mant2 = 8'd209; a_mant3 = 8'd66;
b_mant0 = 8'd31; b_mant1 = 8'd40; b_mant2 = 8'd225; b_mant3 = 8'd132;
a_exp0 = 10'd684; a_exp1 = 10'd671; a_exp2 = 10'd708; a_exp3 = 10'd1010;
b_exp0 = 10'd159; b_exp1 = 10'd566; b_exp2 = 10'd925; b_exp3 = 10'd55;
a_sign0 = 4'd9; a_sign1 = 4'd14; a_sign2 = 4'd1; a_sign3 = 4'd9;
b_sign0 = 4'd9; b_sign1 = 4'd12; b_sign2 = 4'd0; b_sign3 = 4'd11;
@(posedge clk_i);
a_mant0 = 8'd182; a_mant1 = 8'd230; a_mant2 = 8'd98; a_mant3 = 8'd179;
b_mant0 = 8'd223; b_mant1 = 8'd191; b_mant2 = 8'd177; b_mant3 = 8'd191;
a_exp0 = 10'd842; a_exp1 = 10'd376; a_exp2 = 10'd608; a_exp3 = 10'd359;
b_exp0 = 10'd348; b_exp1 = 10'd32; b_exp2 = 10'd208; b_exp3 = 10'd465;
a_sign0 = 4'd1; a_sign1 = 4'd9; a_sign2 = 4'd14; a_sign3 = 4'd2;
b_sign0 = 4'd1; b_sign1 = 4'd0; b_sign2 = 4'd5; b_sign3 = 4'd5;
@(posedge clk_i);
a_mant0 = 8'd23; a_mant1 = 8'd201; a_mant2 = 8'd64; a_mant3 = 8'd225;
b_mant0 = 8'd28; b_mant1 = 8'd172; b_mant2 = 8'd122; b_mant3 = 8'd172;
a_exp0 = 10'd379; a_exp1 = 10'd261; a_exp2 = 10'd653; a_exp3 = 10'd952;
b_exp0 = 10'd736; b_exp1 = 10'd1005; b_exp2 = 10'd950; b_exp3 = 10'd940;
a_sign0 = 4'd11; a_sign1 = 4'd5; a_sign2 = 4'd5; a_sign3 = 4'd15;
b_sign0 = 4'd2; b_sign1 = 4'd15; b_sign2 = 4'd16; b_sign3 = 4'd1;
@(posedge clk_i);
a_mant0 = 8'd215; a_mant1 = 8'd36; a_mant2 = 8'd121; a_mant3 = 8'd134;
b_mant0 = 8'd248; b_mant1 = 8'd143; b_mant2 = 8'd78; b_mant3 = 8'd25;
a_exp0 = 10'd341; a_exp1 = 10'd945; a_exp2 = 10'd660; a_exp3 = 10'd630;
b_exp0 = 10'd367; b_exp1 = 10'd174; b_exp2 = 10'd425; b_exp3 = 10'd985;
a_sign0 = 4'd15; a_sign1 = 4'd0; a_sign2 = 4'd1; a_sign3 = 4'd2;
b_sign0 = 4'd1; b_sign1 = 4'd10; b_sign2 = 4'd0; b_sign3 = 4'd4;
@(posedge clk_i);
a_mant0 = 8'd228; a_mant1 = 8'd98; a_mant2 = 8'd131; a_mant3 = 8'd183;
b_mant0 = 8'd202; b_mant1 = 8'd10; b_mant2 = 8'd82; b_mant3 = 8'd153;
a_exp0 = 10'd438; a_exp1 = 10'd429; a_exp2 = 10'd585; a_exp3 = 10'd150;
b_exp0 = 10'd343; b_exp1 = 10'd887; b_exp2 = 10'd135; b_exp3 = 10'd28;
a_sign0 = 4'd6; a_sign1 = 4'd1; a_sign2 = 4'd7; a_sign3 = 4'd8;
b_sign0 = 4'd9; b_sign1 = 4'd11; b_sign2 = 4'd8; b_sign3 = 4'd15;
@(posedge clk_i);
shared_exps0 = 8'd127;
shared_exps1 = 8'd140;
a_mant0 = 8'd153; a_mant1 = 8'd125; a_mant2 = 8'd204; a_mant3 = 8'd145;
b_mant0 = 8'd129; b_mant1 = 8'd179; b_mant2 = 8'd87; b_mant3 = 8'd168;
a_exp0 = 10'd323; a_exp1 = 10'd404; a_exp2 = 10'd532; a_exp3 = 10'd904;
b_exp0 = 10'd646; b_exp1 = 10'd885; b_exp2 = 10'd893; b_exp3 = 10'd780;
a_sign0 = 4'd6; a_sign1 = 4'd14; a_sign2 = 4'd4; a_sign3 = 4'd10;
b_sign0 = 4'd10; b_sign1 = 4'd14; b_sign2 = 4'd3; b_sign3 = 4'd16;
@(posedge clk_i);
a_mant0 = 8'd151; a_mant1 = 8'd119; a_mant2 = 8'd133; a_mant3 = 8'd163;
b_mant0 = 8'd249; b_mant1 = 8'd236; b_mant2 = 8'd2; b_mant3 = 8'd190;
a_exp0 = 10'd173; a_exp1 = 10'd424; a_exp2 = 10'd740; a_exp3 = 10'd343;
b_exp0 = 10'd906; b_exp1 = 10'd655; b_exp2 = 10'd279; b_exp3 = 10'd195;
a_sign0 = 4'd15; a_sign1 = 4'd1; a_sign2 = 4'd4; a_sign3 = 4'd5;
b_sign0 = 4'd4; b_sign1 = 4'd4; b_sign2 = 4'd8; b_sign3 = 4'd5;
@(posedge clk_i);
a_mant0 = 8'd23; a_mant1 = 8'd240; a_mant2 = 8'd69; a_mant3 = 8'd140;
b_mant0 = 8'd130; b_mant1 = 8'd34; b_mant2 = 8'd59; b_mant3 = 8'd149;
a_exp0 = 10'd1015; a_exp1 = 10'd650; a_exp2 = 10'd880; a_exp3 = 10'd844;
b_exp0 = 10'd773; b_exp1 = 10'd348; b_exp2 = 10'd339; b_exp3 = 10'd517;
a_sign0 = 4'd5; a_sign1 = 4'd3; a_sign2 = 4'd11; a_sign3 = 4'd15;
b_sign0 = 4'd3; b_sign1 = 4'd11; b_sign2 = 4'd0; b_sign3 = 4'd6;
@(posedge clk_i);
a_mant0 = 8'd208; a_mant1 = 8'd154; a_mant2 = 8'd179; a_mant3 = 8'd150;
b_mant0 = 8'd102; b_mant1 = 8'd92; b_mant2 = 8'd218; b_mant3 = 8'd180;
a_exp0 = 10'd134; a_exp1 = 10'd493; a_exp2 = 10'd737; a_exp3 = 10'd731;
b_exp0 = 10'd128; b_exp1 = 10'd100; b_exp2 = 10'd352; b_exp3 = 10'd562;
a_sign0 = 4'd15; a_sign1 = 4'd12; a_sign2 = 4'd0; a_sign3 = 4'd10;
b_sign0 = 4'd3; b_sign1 = 4'd3; b_sign2 = 4'd2; b_sign3 = 4'd3;
@(posedge clk_i);
a_mant0 = 8'd70; a_mant1 = 8'd40; a_mant2 = 8'd53; a_mant3 = 8'd98;
b_mant0 = 8'd91; b_mant1 = 8'd225; b_mant2 = 8'd97; b_mant3 = 8'd126;
a_exp0 = 10'd658; a_exp1 = 10'd626; a_exp2 = 10'd18; a_exp3 = 10'd341;
b_exp0 = 10'd588; b_exp1 = 10'd926; b_exp2 = 10'd80; b_exp3 = 10'd912;
a_sign0 = 4'd13; a_sign1 = 4'd0; a_sign2 = 4'd3; a_sign3 = 4'd13;
b_sign0 = 4'd12; b_sign1 = 4'd9; b_sign2 = 4'd10; b_sign3 = 4'd15;
@(posedge clk_i);
a_mant0 = 8'd199; a_mant1 = 8'd215; a_mant2 = 8'd11; a_mant3 = 8'd180;
b_mant0 = 8'd53; b_mant1 = 8'd191; b_mant2 = 8'd113; b_mant3 = 8'd54;
a_exp0 = 10'd165; a_exp1 = 10'd831; a_exp2 = 10'd586; a_exp3 = 10'd469;
b_exp0 = 10'd914; b_exp1 = 10'd1017; b_exp2 = 10'd893; b_exp3 = 10'd944;
a_sign0 = 4'd5; a_sign1 = 4'd4; a_sign2 = 4'd7; a_sign3 = 4'd10;
b_sign0 = 4'd14; b_sign1 = 4'd2; b_sign2 = 4'd13; b_sign3 = 4'd1;
@(posedge clk_i);
a_mant0 = 8'd74; a_mant1 = 8'd109; a_mant2 = 8'd68; a_mant3 = 8'd194;
b_mant0 = 8'd233; b_mant1 = 8'd32; b_mant2 = 8'd84; b_mant3 = 8'd61;
a_exp0 = 10'd800; a_exp1 = 10'd904; a_exp2 = 10'd983; a_exp3 = 10'd256;
b_exp0 = 10'd827; b_exp1 = 10'd31; b_exp2 = 10'd880; b_exp3 = 10'd960;
a_sign0 = 4'd11; a_sign1 = 4'd3; a_sign2 = 4'd1; a_sign3 = 4'd2;
b_sign0 = 4'd3; b_sign1 = 4'd8; b_sign2 = 4'd16; b_sign3 = 4'd11;
@(posedge clk_i);
a_mant0 = 8'd111; a_mant1 = 8'd153; a_mant2 = 8'd158; a_mant3 = 8'd156;
b_mant0 = 8'd79; b_mant1 = 8'd251; b_mant2 = 8'd206; b_mant3 = 8'd214;
a_exp0 = 10'd601; a_exp1 = 10'd264; a_exp2 = 10'd749; a_exp3 = 10'd990;
b_exp0 = 10'd570; b_exp1 = 10'd116; b_exp2 = 10'd192; b_exp3 = 10'd142;
a_sign0 = 4'd11; a_sign1 = 4'd12; a_sign2 = 4'd12; a_sign3 = 4'd1;
b_sign0 = 4'd3; b_sign1 = 4'd15; b_sign2 = 4'd5; b_sign3 = 4'd12;
@(posedge clk_i);
shared_exps0 = 8'd122;
shared_exps1 = 8'd123;
a_mant0 = 8'd7; a_mant1 = 8'd222; a_mant2 = 8'd45; a_mant3 = 8'd20;
b_mant0 = 8'd146; b_mant1 = 8'd142; b_mant2 = 8'd67; b_mant3 = 8'd133;
a_exp0 = 10'd111; a_exp1 = 10'd158; a_exp2 = 10'd530; a_exp3 = 10'd433;
b_exp0 = 10'd826; b_exp1 = 10'd670; b_exp2 = 10'd1000; b_exp3 = 10'd904;
a_sign0 = 4'd14; a_sign1 = 4'd4; a_sign2 = 4'd16; a_sign3 = 4'd0;
b_sign0 = 4'd7; b_sign1 = 4'd12; b_sign2 = 4'd16; b_sign3 = 4'd11;
@(posedge clk_i);
a_mant0 = 8'd186; a_mant1 = 8'd36; a_mant2 = 8'd150; a_mant3 = 8'd145;
b_mant0 = 8'd57; b_mant1 = 8'd125; b_mant2 = 8'd48; b_mant3 = 8'd104;
a_exp0 = 10'd986; a_exp1 = 10'd830; a_exp2 = 10'd752; a_exp3 = 10'd66;
b_exp0 = 10'd777; b_exp1 = 10'd286; b_exp2 = 10'd52; b_exp3 = 10'd236;
a_sign0 = 4'd8; a_sign1 = 4'd15; a_sign2 = 4'd13; a_sign3 = 4'd8;
b_sign0 = 4'd1; b_sign1 = 4'd2; b_sign2 = 4'd16; b_sign3 = 4'd12;
@(posedge clk_i);
a_mant0 = 8'd3; a_mant1 = 8'd230; a_mant2 = 8'd143; a_mant3 = 8'd179;
b_mant0 = 8'd5; b_mant1 = 8'd58; b_mant2 = 8'd49; b_mant3 = 8'd51;
a_exp0 = 10'd53; a_exp1 = 10'd274; a_exp2 = 10'd673; a_exp3 = 10'd339;
b_exp0 = 10'd317; b_exp1 = 10'd112; b_exp2 = 10'd38; b_exp3 = 10'd381;
a_sign0 = 4'd10; a_sign1 = 4'd7; a_sign2 = 4'd8; a_sign3 = 4'd14;
b_sign0 = 4'd9; b_sign1 = 4'd15; b_sign2 = 4'd5; b_sign3 = 4'd8;
@(posedge clk_i);
a_mant0 = 8'd81; a_mant1 = 8'd230; a_mant2 = 8'd230; a_mant3 = 8'd21;
b_mant0 = 8'd111; b_mant1 = 8'd70; b_mant2 = 8'd197; b_mant3 = 8'd67;
a_exp0 = 10'd438; a_exp1 = 10'd410; a_exp2 = 10'd233; a_exp3 = 10'd549;
b_exp0 = 10'd561; b_exp1 = 10'd723; b_exp2 = 10'd160; b_exp3 = 10'd865;
a_sign0 = 4'd15; a_sign1 = 4'd7; a_sign2 = 4'd2; a_sign3 = 4'd9;
b_sign0 = 4'd5; b_sign1 = 4'd10; b_sign2 = 4'd11; b_sign3 = 4'd15;
@(posedge clk_i);
a_mant0 = 8'd153; a_mant1 = 8'd177; a_mant2 = 8'd193; a_mant3 = 8'd130;
b_mant0 = 8'd166; b_mant1 = 8'd22; b_mant2 = 8'd206; b_mant3 = 8'd95;
a_exp0 = 10'd546; a_exp1 = 10'd156; a_exp2 = 10'd715; a_exp3 = 10'd143;
b_exp0 = 10'd321; b_exp1 = 10'd942; b_exp2 = 10'd189; b_exp3 = 10'd695;
a_sign0 = 4'd15; a_sign1 = 4'd2; a_sign2 = 4'd10; a_sign3 = 4'd1;
b_sign0 = 4'd5; b_sign1 = 4'd5; b_sign2 = 4'd4; b_sign3 = 4'd6;
@(posedge clk_i);
a_mant0 = 8'd75; a_mant1 = 8'd65; a_mant2 = 8'd105; a_mant3 = 8'd106;
b_mant0 = 8'd79; b_mant1 = 8'd254; b_mant2 = 8'd159; b_mant3 = 8'd166;
a_exp0 = 10'd630; a_exp1 = 10'd931; a_exp2 = 10'd592; a_exp3 = 10'd885;
b_exp0 = 10'd270; b_exp1 = 10'd517; b_exp2 = 10'd150; b_exp3 = 10'd981;
a_sign0 = 4'd7; a_sign1 = 4'd9; a_sign2 = 4'd1; a_sign3 = 4'd14;
b_sign0 = 4'd15; b_sign1 = 4'd15; b_sign2 = 4'd15; b_sign3 = 4'd11;
@(posedge clk_i);
a_mant0 = 8'd195; a_mant1 = 8'd118; a_mant2 = 8'd243; a_mant3 = 8'd208;
b_mant0 = 8'd85; b_mant1 = 8'd139; b_mant2 = 8'd111; b_mant3 = 8'd145;
a_exp0 = 10'd865; a_exp1 = 10'd668; a_exp2 = 10'd440; a_exp3 = 10'd990;
b_exp0 = 10'd620; b_exp1 = 10'd372; b_exp2 = 10'd404; b_exp3 = 10'd698;
a_sign0 = 4'd5; a_sign1 = 4'd11; a_sign2 = 4'd15; a_sign3 = 4'd10;
b_sign0 = 4'd13; b_sign1 = 4'd16; b_sign2 = 4'd6; b_sign3 = 4'd0;
@(posedge clk_i);
a_mant0 = 8'd143; a_mant1 = 8'd42; a_mant2 = 8'd82; a_mant3 = 8'd224;
b_mant0 = 8'd217; b_mant1 = 8'd121; b_mant2 = 8'd78; b_mant3 = 8'd171;
a_exp0 = 10'd44; a_exp1 = 10'd959; a_exp2 = 10'd887; a_exp3 = 10'd311;
b_exp0 = 10'd93; b_exp1 = 10'd448; b_exp2 = 10'd861; b_exp3 = 10'd553;
a_sign0 = 4'd0; a_sign1 = 4'd2; a_sign2 = 4'd7; a_sign3 = 4'd15;
b_sign0 = 4'd11; b_sign1 = 4'd2; b_sign2 = 4'd3; b_sign3 = 4'd6;
@(posedge clk_i);
shared_exps0 = 8'd157;
shared_exps1 = 8'd120;
rstn = 0;
@(posedge clk_i);
rstn = 1;
a_mant0 = 8'd129; a_mant1 = 8'd12; a_mant2 = 8'd29; a_mant3 = 8'd97;
b_mant0 = 8'd178; b_mant1 = 8'd151; b_mant2 = 8'd16; b_mant3 = 8'd27;
a_exp0 = 10'd934; a_exp1 = 10'd168; a_exp2 = 10'd949; a_exp3 = 10'd929;
b_exp0 = 10'd237; b_exp1 = 10'd746; b_exp2 = 10'd172; b_exp3 = 10'd467;
a_sign0 = 4'd0; a_sign1 = 4'd0; a_sign2 = 4'd7; a_sign3 = 4'd16;
b_sign0 = 4'd4; b_sign1 = 4'd1; b_sign2 = 4'd3; b_sign3 = 4'd12;
@(posedge clk_i);
a_mant0 = 8'd174; a_mant1 = 8'd59; a_mant2 = 8'd60; a_mant3 = 8'd81;
b_mant0 = 8'd84; b_mant1 = 8'd110; b_mant2 = 8'd180; b_mant3 = 8'd216;
a_exp0 = 10'd477; a_exp1 = 10'd725; a_exp2 = 10'd933; a_exp3 = 10'd513;
b_exp0 = 10'd141; b_exp1 = 10'd120; b_exp2 = 10'd981; b_exp3 = 10'd86;
a_sign0 = 4'd15; a_sign1 = 4'd2; a_sign2 = 4'd3; a_sign3 = 4'd6;
b_sign0 = 4'd5; b_sign1 = 4'd9; b_sign2 = 4'd13; b_sign3 = 4'd7;
@(posedge clk_i);
a_mant0 = 8'd169; a_mant1 = 8'd97; a_mant2 = 8'd81; a_mant3 = 8'd69;
b_mant0 = 8'd165; b_mant1 = 8'd82; b_mant2 = 8'd108; b_mant3 = 8'd140;
a_exp0 = 10'd679; a_exp1 = 10'd332; a_exp2 = 10'd675; a_exp3 = 10'd365;
b_exp0 = 10'd286; b_exp1 = 10'd21; b_exp2 = 10'd21; b_exp3 = 10'd906;
a_sign0 = 4'd0; a_sign1 = 4'd7; a_sign2 = 4'd0; a_sign3 = 4'd14;
b_sign0 = 4'd8; b_sign1 = 4'd5; b_sign2 = 4'd6; b_sign3 = 4'd5;
@(posedge clk_i);
a_mant0 = 8'd2; a_mant1 = 8'd240; a_mant2 = 8'd179; a_mant3 = 8'd155;
b_mant0 = 8'd33; b_mant1 = 8'd21; b_mant2 = 8'd150; b_mant3 = 8'd212;
a_exp0 = 10'd250; a_exp1 = 10'd780; a_exp2 = 10'd98; a_exp3 = 10'd868;
b_exp0 = 10'd97; b_exp1 = 10'd760; b_exp2 = 10'd258; b_exp3 = 10'd492;
a_sign0 = 4'd1; a_sign1 = 4'd4; a_sign2 = 4'd2; a_sign3 = 4'd15;
b_sign0 = 4'd13; b_sign1 = 4'd15; b_sign2 = 4'd15; b_sign3 = 4'd14;
@(posedge clk_i);
a_mant0 = 8'd15; a_mant1 = 8'd240; a_mant2 = 8'd188; a_mant3 = 8'd223;
b_mant0 = 8'd133; b_mant1 = 8'd21; b_mant2 = 8'd40; b_mant3 = 8'd7;
a_exp0 = 10'd683; a_exp1 = 10'd601; a_exp2 = 10'd979; a_exp3 = 10'd503;
b_exp0 = 10'd873; b_exp1 = 10'd723; b_exp2 = 10'd403; b_exp3 = 10'd332;
a_sign0 = 4'd1; a_sign1 = 4'd16; a_sign2 = 4'd8; a_sign3 = 4'd16;
b_sign0 = 4'd4; b_sign1 = 4'd1; b_sign2 = 4'd6; b_sign3 = 4'd2;
@(posedge clk_i);
a_mant0 = 8'd176; a_mant1 = 8'd98; a_mant2 = 8'd226; a_mant3 = 8'd195;
b_mant0 = 8'd105; b_mant1 = 8'd55; b_mant2 = 8'd140; b_mant3 = 8'd185;
a_exp0 = 10'd394; a_exp1 = 10'd329; a_exp2 = 10'd274; a_exp3 = 10'd224;
b_exp0 = 10'd889; b_exp1 = 10'd103; b_exp2 = 10'd807; b_exp3 = 10'd428;
a_sign0 = 4'd15; a_sign1 = 4'd6; a_sign2 = 4'd13; a_sign3 = 4'd11;
b_sign0 = 4'd5; b_sign1 = 4'd16; b_sign2 = 4'd12; b_sign3 = 4'd9;
@(posedge clk_i);
a_mant0 = 8'd87; a_mant1 = 8'd229; a_mant2 = 8'd104; a_mant3 = 8'd242;
b_mant0 = 8'd10; b_mant1 = 8'd230; b_mant2 = 8'd91; b_mant3 = 8'd251;
a_exp0 = 10'd117; a_exp1 = 10'd521; a_exp2 = 10'd90; a_exp3 = 10'd958;
b_exp0 = 10'd996; b_exp1 = 10'd690; b_exp2 = 10'd330; b_exp3 = 10'd707;
a_sign0 = 4'd13; a_sign1 = 4'd9; a_sign2 = 4'd13; a_sign3 = 4'd2;
b_sign0 = 4'd12; b_sign1 = 4'd0; b_sign2 = 4'd6; b_sign3 = 4'd15;
@(posedge clk_i);
shared_exps0 = 8'd115;
shared_exps1 = 8'd135;
a_mant0 = 8'd215; a_mant1 = 8'd109; a_mant2 = 8'd199; a_mant3 = 8'd129;
b_mant0 = 8'd178; b_mant1 = 8'd45; b_mant2 = 8'd28; b_mant3 = 8'd156;
a_exp0 = 10'd972; a_exp1 = 10'd383; a_exp2 = 10'd584; a_exp3 = 10'd768;
b_exp0 = 10'd232; b_exp1 = 10'd343; b_exp2 = 10'd60; b_exp3 = 10'd257;
a_sign0 = 4'd14; a_sign1 = 4'd1; a_sign2 = 4'd10; a_sign3 = 4'd8;
b_sign0 = 4'd2; b_sign1 = 4'd2; b_sign2 = 4'd8; b_sign3 = 4'd15;
@(posedge clk_i);
a_mant0 = 8'd149; a_mant1 = 8'd122; a_mant2 = 8'd193; a_mant3 = 8'd150;
b_mant0 = 8'd227; b_mant1 = 8'd135; b_mant2 = 8'd206; b_mant3 = 8'd96;
a_exp0 = 10'd985; a_exp1 = 10'd69; a_exp2 = 10'd336; a_exp3 = 10'd608;
b_exp0 = 10'd999; b_exp1 = 10'd732; b_exp2 = 10'd604; b_exp3 = 10'd937;
a_sign0 = 4'd12; a_sign1 = 4'd2; a_sign2 = 4'd15; a_sign3 = 4'd7;
b_sign0 = 4'd3; b_sign1 = 4'd7; b_sign2 = 4'd4; b_sign3 = 4'd4;
@(posedge clk_i);
a_mant0 = 8'd191; a_mant1 = 8'd114; a_mant2 = 8'd30; a_mant3 = 8'd241;
b_mant0 = 8'd22; b_mant1 = 8'd69; b_mant2 = 8'd97; b_mant3 = 8'd110;
a_exp0 = 10'd212; a_exp1 = 10'd388; a_exp2 = 10'd722; a_exp3 = 10'd818;
b_exp0 = 10'd194; b_exp1 = 10'd712; b_exp2 = 10'd848; b_exp3 = 10'd1;
a_sign0 = 4'd2; a_sign1 = 4'd8; a_sign2 = 4'd11; a_sign3 = 4'd9;
b_sign0 = 4'd2; b_sign1 = 4'd5; b_sign2 = 4'd14; b_sign3 = 4'd9;
@(posedge clk_i);
a_mant0 = 8'd77; a_mant1 = 8'd74; a_mant2 = 8'd162; a_mant3 = 8'd126;
b_mant0 = 8'd86; b_mant1 = 8'd169; b_mant2 = 8'd204; b_mant3 = 8'd104;
a_exp0 = 10'd930; a_exp1 = 10'd932; a_exp2 = 10'd863; a_exp3 = 10'd5;
b_exp0 = 10'd871; b_exp1 = 10'd334; b_exp2 = 10'd640; b_exp3 = 10'd971;
a_sign0 = 4'd16; a_sign1 = 4'd0; a_sign2 = 4'd2; a_sign3 = 4'd9;
b_sign0 = 4'd3; b_sign1 = 4'd10; b_sign2 = 4'd1; b_sign3 = 4'd3;
@(posedge clk_i);
a_mant0 = 8'd158; a_mant1 = 8'd180; a_mant2 = 8'd178; a_mant3 = 8'd56;
b_mant0 = 8'd59; b_mant1 = 8'd109; b_mant2 = 8'd176; b_mant3 = 8'd238;
a_exp0 = 10'd712; a_exp1 = 10'd671; a_exp2 = 10'd444; a_exp3 = 10'd1014;
b_exp0 = 10'd977; b_exp1 = 10'd600; b_exp2 = 10'd50; b_exp3 = 10'd974;
a_sign0 = 4'd2; a_sign1 = 4'd7; a_sign2 = 4'd16; a_sign3 = 4'd9;
b_sign0 = 4'd3; b_sign1 = 4'd5; b_sign2 = 4'd4; b_sign3 = 4'd6;
@(posedge clk_i);
a_mant0 = 8'd39; a_mant1 = 8'd203; a_mant2 = 8'd113; a_mant3 = 8'd128;
b_mant0 = 8'd22; b_mant1 = 8'd133; b_mant2 = 8'd4; b_mant3 = 8'd228;
a_exp0 = 10'd702; a_exp1 = 10'd206; a_exp2 = 10'd954; a_exp3 = 10'd338;
b_exp0 = 10'd63; b_exp1 = 10'd796; b_exp2 = 10'd50; b_exp3 = 10'd643;
a_sign0 = 4'd14; a_sign1 = 4'd11; a_sign2 = 4'd7; a_sign3 = 4'd6;
b_sign0 = 4'd7; b_sign1 = 4'd8; b_sign2 = 4'd1; b_sign3 = 4'd4;
@(posedge clk_i);
a_mant0 = 8'd158; a_mant1 = 8'd1; a_mant2 = 8'd90; a_mant3 = 8'd22;
b_mant0 = 8'd148; b_mant1 = 8'd51; b_mant2 = 8'd183; b_mant3 = 8'd6;
a_exp0 = 10'd735; a_exp1 = 10'd915; a_exp2 = 10'd118; a_exp3 = 10'd1012;
b_exp0 = 10'd901; b_exp1 = 10'd896; b_exp2 = 10'd613; b_exp3 = 10'd161;
a_sign0 = 4'd15; a_sign1 = 4'd9; a_sign2 = 4'd13; a_sign3 = 4'd0;
b_sign0 = 4'd10; b_sign1 = 4'd8; b_sign2 = 4'd13; b_sign3 = 4'd16;
@(posedge clk_i);
a_mant0 = 8'd102; a_mant1 = 8'd107; a_mant2 = 8'd40; a_mant3 = 8'd59;
b_mant0 = 8'd106; b_mant1 = 8'd85; b_mant2 = 8'd109; b_mant3 = 8'd154;
a_exp0 = 10'd81; a_exp1 = 10'd552; a_exp2 = 10'd904; a_exp3 = 10'd985;
b_exp0 = 10'd104; b_exp1 = 10'd158; b_exp2 = 10'd179; b_exp3 = 10'd549;
a_sign0 = 4'd9; a_sign1 = 4'd14; a_sign2 = 4'd11; a_sign3 = 4'd3;
b_sign0 = 4'd0; b_sign1 = 4'd7; b_sign2 = 4'd5; b_sign3 = 4'd15;
@(posedge clk_i);
shared_exps0 = 8'd131;
shared_exps1 = 8'd107;
a_mant0 = 8'd97; a_mant1 = 8'd126; a_mant2 = 8'd93; a_mant3 = 8'd109;
b_mant0 = 8'd163; b_mant1 = 8'd135; b_mant2 = 8'd104; b_mant3 = 8'd39;
a_exp0 = 10'd59; a_exp1 = 10'd874; a_exp2 = 10'd650; a_exp3 = 10'd435;
b_exp0 = 10'd742; b_exp1 = 10'd193; b_exp2 = 10'd1021; b_exp3 = 10'd502;
a_sign0 = 4'd3; a_sign1 = 4'd4; a_sign2 = 4'd0; a_sign3 = 4'd6;
b_sign0 = 4'd12; b_sign1 = 4'd13; b_sign2 = 4'd0; b_sign3 = 4'd10;
@(posedge clk_i);
a_mant0 = 8'd162; a_mant1 = 8'd182; a_mant2 = 8'd177; a_mant3 = 8'd237;
b_mant0 = 8'd168; b_mant1 = 8'd95; b_mant2 = 8'd219; b_mant3 = 8'd118;
a_exp0 = 10'd985; a_exp1 = 10'd73; a_exp2 = 10'd500; a_exp3 = 10'd883;
b_exp0 = 10'd607; b_exp1 = 10'd918; b_exp2 = 10'd865; b_exp3 = 10'd84;
a_sign0 = 4'd6; a_sign1 = 4'd3; a_sign2 = 4'd6; a_sign3 = 4'd16;
b_sign0 = 4'd4; b_sign1 = 4'd13; b_sign2 = 4'd13; b_sign3 = 4'd1;
@(posedge clk_i);
a_mant0 = 8'd194; a_mant1 = 8'd11; a_mant2 = 8'd143; a_mant3 = 8'd141;
b_mant0 = 8'd165; b_mant1 = 8'd56; b_mant2 = 8'd93; b_mant3 = 8'd46;
a_exp0 = 10'd753; a_exp1 = 10'd769; a_exp2 = 10'd826; a_exp3 = 10'd916;
b_exp0 = 10'd753; b_exp1 = 10'd892; b_exp2 = 10'd83; b_exp3 = 10'd776;
a_sign0 = 4'd6; a_sign1 = 4'd15; a_sign2 = 4'd6; a_sign3 = 4'd15;
b_sign0 = 4'd6; b_sign1 = 4'd1; b_sign2 = 4'd11; b_sign3 = 4'd7;
@(posedge clk_i);
a_mant0 = 8'd44; a_mant1 = 8'd70; a_mant2 = 8'd125; a_mant3 = 8'd215;
b_mant0 = 8'd17; b_mant1 = 8'd134; b_mant2 = 8'd124; b_mant3 = 8'd121;
a_exp0 = 10'd550; a_exp1 = 10'd258; a_exp2 = 10'd291; a_exp3 = 10'd397;
b_exp0 = 10'd138; b_exp1 = 10'd437; b_exp2 = 10'd192; b_exp3 = 10'd230;
a_sign0 = 4'd7; a_sign1 = 4'd15; a_sign2 = 4'd10; a_sign3 = 4'd2;
b_sign0 = 4'd8; b_sign1 = 4'd9; b_sign2 = 4'd12; b_sign3 = 4'd6;
@(posedge clk_i);
a_mant0 = 8'd206; a_mant1 = 8'd56; a_mant2 = 8'd217; a_mant3 = 8'd161;
b_mant0 = 8'd54; b_mant1 = 8'd90; b_mant2 = 8'd176; b_mant3 = 8'd205;
a_exp0 = 10'd787; a_exp1 = 10'd458; a_exp2 = 10'd953; a_exp3 = 10'd300;
b_exp0 = 10'd648; b_exp1 = 10'd159; b_exp2 = 10'd342; b_exp3 = 10'd850;
a_sign0 = 4'd0; a_sign1 = 4'd15; a_sign2 = 4'd13; a_sign3 = 4'd1;
b_sign0 = 4'd15; b_sign1 = 4'd10; b_sign2 = 4'd1; b_sign3 = 4'd6;
@(posedge clk_i);
a_mant0 = 8'd180; a_mant1 = 8'd75; a_mant2 = 8'd168; a_mant3 = 8'd208;
b_mant0 = 8'd233; b_mant1 = 8'd92; b_mant2 = 8'd110; b_mant3 = 8'd31;
a_exp0 = 10'd406; a_exp1 = 10'd360; a_exp2 = 10'd204; a_exp3 = 10'd109;
b_exp0 = 10'd412; b_exp1 = 10'd371; b_exp2 = 10'd809; b_exp3 = 10'd678;
a_sign0 = 4'd0; a_sign1 = 4'd3; a_sign2 = 4'd12; a_sign3 = 4'd9;
b_sign0 = 4'd2; b_sign1 = 4'd5; b_sign2 = 4'd14; b_sign3 = 4'd7;
@(posedge clk_i);
a_mant0 = 8'd25; a_mant1 = 8'd9; a_mant2 = 8'd210; a_mant3 = 8'd184;
b_mant0 = 8'd243; b_mant1 = 8'd18; b_mant2 = 8'd233; b_mant3 = 8'd78;
a_exp0 = 10'd69; a_exp1 = 10'd951; a_exp2 = 10'd961; a_exp3 = 10'd37;
b_exp0 = 10'd905; b_exp1 = 10'd916; b_exp2 = 10'd634; b_exp3 = 10'd416;
a_sign0 = 4'd13; a_sign1 = 4'd9; a_sign2 = 4'd11; a_sign3 = 4'd12;
b_sign0 = 4'd0; b_sign1 = 4'd13; b_sign2 = 4'd0; b_sign3 = 4'd13;
@(posedge clk_i);
a_mant0 = 8'd188; a_mant1 = 8'd118; a_mant2 = 8'd126; a_mant3 = 8'd41;
b_mant0 = 8'd179; b_mant1 = 8'd20; b_mant2 = 8'd254; b_mant3 = 8'd0;
a_exp0 = 10'd224; a_exp1 = 10'd6; a_exp2 = 10'd50; a_exp3 = 10'd327;
b_exp0 = 10'd868; b_exp1 = 10'd392; b_exp2 = 10'd274; b_exp3 = 10'd416;
a_sign0 = 4'd15; a_sign1 = 4'd2; a_sign2 = 4'd5; a_sign3 = 4'd6;
b_sign0 = 4'd13; b_sign1 = 4'd9; b_sign2 = 4'd11; b_sign3 = 4'd7;
@(posedge clk_i);
shared_exps0 = 8'd103;
shared_exps1 = 8'd133;
a_mant0 = 8'd189; a_mant1 = 8'd148; a_mant2 = 8'd104; a_mant3 = 8'd112;
b_mant0 = 8'd52; b_mant1 = 8'd221; b_mant2 = 8'd168; b_mant3 = 8'd75;
a_exp0 = 10'd272; a_exp1 = 10'd248; a_exp2 = 10'd72; a_exp3 = 10'd766;
b_exp0 = 10'd166; b_exp1 = 10'd534; b_exp2 = 10'd259; b_exp3 = 10'd41;
a_sign0 = 4'd13; a_sign1 = 4'd4; a_sign2 = 4'd16; a_sign3 = 4'd12;
b_sign0 = 4'd16; b_sign1 = 4'd5; b_sign2 = 4'd2; b_sign3 = 4'd2;
@(posedge clk_i);
a_mant0 = 8'd130; a_mant1 = 8'd183; a_mant2 = 8'd48; a_mant3 = 8'd179;
b_mant0 = 8'd156; b_mant1 = 8'd72; b_mant2 = 8'd245; b_mant3 = 8'd150;
a_exp0 = 10'd465; a_exp1 = 10'd635; a_exp2 = 10'd466; a_exp3 = 10'd340;
b_exp0 = 10'd813; b_exp1 = 10'd241; b_exp2 = 10'd798; b_exp3 = 10'd422;
a_sign0 = 4'd9; a_sign1 = 4'd11; a_sign2 = 4'd4; a_sign3 = 4'd12;
b_sign0 = 4'd16; b_sign1 = 4'd16; b_sign2 = 4'd14; b_sign3 = 4'd16;
@(posedge clk_i);
a_mant0 = 8'd80; a_mant1 = 8'd92; a_mant2 = 8'd63; a_mant3 = 8'd135;
b_mant0 = 8'd180; b_mant1 = 8'd56; b_mant2 = 8'd43; b_mant3 = 8'd41;
a_exp0 = 10'd843; a_exp1 = 10'd55; a_exp2 = 10'd414; a_exp3 = 10'd447;
b_exp0 = 10'd451; b_exp1 = 10'd765; b_exp2 = 10'd373; b_exp3 = 10'd671;
a_sign0 = 4'd7; a_sign1 = 4'd9; a_sign2 = 4'd6; a_sign3 = 4'd11;
b_sign0 = 4'd10; b_sign1 = 4'd7; b_sign2 = 4'd5; b_sign3 = 4'd7;
@(posedge clk_i);
a_mant0 = 8'd164; a_mant1 = 8'd149; a_mant2 = 8'd54; a_mant3 = 8'd54;
b_mant0 = 8'd45; b_mant1 = 8'd108; b_mant2 = 8'd81; b_mant3 = 8'd4;
a_exp0 = 10'd322; a_exp1 = 10'd835; a_exp2 = 10'd367; a_exp3 = 10'd332;
b_exp0 = 10'd476; b_exp1 = 10'd824; b_exp2 = 10'd6; b_exp3 = 10'd916;
a_sign0 = 4'd4; a_sign1 = 4'd7; a_sign2 = 4'd1; a_sign3 = 4'd12;
b_sign0 = 4'd13; b_sign1 = 4'd11; b_sign2 = 4'd7; b_sign3 = 4'd13;
@(posedge clk_i);
a_mant0 = 8'd12; a_mant1 = 8'd122; a_mant2 = 8'd36; a_mant3 = 8'd159;
b_mant0 = 8'd217; b_mant1 = 8'd253; b_mant2 = 8'd67; b_mant3 = 8'd178;
a_exp0 = 10'd155; a_exp1 = 10'd82; a_exp2 = 10'd429; a_exp3 = 10'd971;
b_exp0 = 10'd498; b_exp1 = 10'd750; b_exp2 = 10'd444; b_exp3 = 10'd498;
a_sign0 = 4'd10; a_sign1 = 4'd15; a_sign2 = 4'd14; a_sign3 = 4'd1;
b_sign0 = 4'd9; b_sign1 = 4'd3; b_sign2 = 4'd13; b_sign3 = 4'd10;
@(posedge clk_i);
a_mant0 = 8'd245; a_mant1 = 8'd230; a_mant2 = 8'd149; a_mant3 = 8'd72;
b_mant0 = 8'd32; b_mant1 = 8'd61; b_mant2 = 8'd106; b_mant3 = 8'd21;
a_exp0 = 10'd502; a_exp1 = 10'd59; a_exp2 = 10'd32; a_exp3 = 10'd320;
b_exp0 = 10'd852; b_exp1 = 10'd703; b_exp2 = 10'd131; b_exp3 = 10'd26;
a_sign0 = 4'd8; a_sign1 = 4'd14; a_sign2 = 4'd10; a_sign3 = 4'd3;
b_sign0 = 4'd6; b_sign1 = 4'd11; b_sign2 = 4'd13; b_sign3 = 4'd0;
@(posedge clk_i);
a_mant0 = 8'd74; a_mant1 = 8'd153; a_mant2 = 8'd54; a_mant3 = 8'd185;
b_mant0 = 8'd159; b_mant1 = 8'd169; b_mant2 = 8'd6; b_mant3 = 8'd159;
a_exp0 = 10'd88; a_exp1 = 10'd100; a_exp2 = 10'd977; a_exp3 = 10'd283;
b_exp0 = 10'd392; b_exp1 = 10'd741; b_exp2 = 10'd283; b_exp3 = 10'd601;
a_sign0 = 4'd6; a_sign1 = 4'd13; a_sign2 = 4'd1; a_sign3 = 4'd13;
b_sign0 = 4'd16; b_sign1 = 4'd9; b_sign2 = 4'd1; b_sign3 = 4'd14;
@(posedge clk_i);
a_mant0 = 8'd193; a_mant1 = 8'd240; a_mant2 = 8'd23; a_mant3 = 8'd150;
b_mant0 = 8'd167; b_mant1 = 8'd43; b_mant2 = 8'd69; b_mant3 = 8'd6;
a_exp0 = 10'd194; a_exp1 = 10'd200; a_exp2 = 10'd926; a_exp3 = 10'd794;
b_exp0 = 10'd163; b_exp1 = 10'd623; b_exp2 = 10'd738; b_exp3 = 10'd458;
a_sign0 = 4'd0; a_sign1 = 4'd1; a_sign2 = 4'd2; a_sign3 = 4'd13;
b_sign0 = 4'd4; b_sign1 = 4'd12; b_sign2 = 4'd12; b_sign3 = 4'd13;
@(posedge clk_i);
shared_exps0 = 8'd146;
shared_exps1 = 8'd134;
rstn = 0;
@(posedge clk_i);
rstn = 1;
a_mant0 = 8'd13; a_mant1 = 8'd17; a_mant2 = 8'd204; a_mant3 = 8'd120;
b_mant0 = 8'd136; b_mant1 = 8'd124; b_mant2 = 8'd3; b_mant3 = 8'd48;
a_exp0 = 10'd501; a_exp1 = 10'd155; a_exp2 = 10'd897; a_exp3 = 10'd89;
b_exp0 = 10'd729; b_exp1 = 10'd593; b_exp2 = 10'd190; b_exp3 = 10'd935;
a_sign0 = 4'd8; a_sign1 = 4'd5; a_sign2 = 4'd5; a_sign3 = 4'd1;
b_sign0 = 4'd2; b_sign1 = 4'd8; b_sign2 = 4'd2; b_sign3 = 4'd13;
@(posedge clk_i);
a_mant0 = 8'd64; a_mant1 = 8'd170; a_mant2 = 8'd245; a_mant3 = 8'd179;
b_mant0 = 8'd59; b_mant1 = 8'd157; b_mant2 = 8'd140; b_mant3 = 8'd167;
a_exp0 = 10'd679; a_exp1 = 10'd211; a_exp2 = 10'd888; a_exp3 = 10'd625;
b_exp0 = 10'd210; b_exp1 = 10'd807; b_exp2 = 10'd567; b_exp3 = 10'd214;
a_sign0 = 4'd12; a_sign1 = 4'd1; a_sign2 = 4'd7; a_sign3 = 4'd10;
b_sign0 = 4'd10; b_sign1 = 4'd8; b_sign2 = 4'd5; b_sign3 = 4'd10;
@(posedge clk_i);
a_mant0 = 8'd250; a_mant1 = 8'd19; a_mant2 = 8'd29; a_mant3 = 8'd212;
b_mant0 = 8'd26; b_mant1 = 8'd128; b_mant2 = 8'd178; b_mant3 = 8'd133;
a_exp0 = 10'd201; a_exp1 = 10'd211; a_exp2 = 10'd872; a_exp3 = 10'd355;
b_exp0 = 10'd245; b_exp1 = 10'd729; b_exp2 = 10'd622; b_exp3 = 10'd958;
a_sign0 = 4'd0; a_sign1 = 4'd15; a_sign2 = 4'd9; a_sign3 = 4'd10;
b_sign0 = 4'd9; b_sign1 = 4'd15; b_sign2 = 4'd12; b_sign3 = 4'd16;
@(posedge clk_i);
a_mant0 = 8'd225; a_mant1 = 8'd220; a_mant2 = 8'd209; a_mant3 = 8'd112;
b_mant0 = 8'd4; b_mant1 = 8'd25; b_mant2 = 8'd122; b_mant3 = 8'd18;
a_exp0 = 10'd13; a_exp1 = 10'd267; a_exp2 = 10'd780; a_exp3 = 10'd798;
b_exp0 = 10'd824; b_exp1 = 10'd638; b_exp2 = 10'd22; b_exp3 = 10'd1001;
a_sign0 = 4'd0; a_sign1 = 4'd1; a_sign2 = 4'd5; a_sign3 = 4'd10;
b_sign0 = 4'd10; b_sign1 = 4'd13; b_sign2 = 4'd9; b_sign3 = 4'd2;
@(posedge clk_i);
a_mant0 = 8'd243; a_mant1 = 8'd212; a_mant2 = 8'd181; a_mant3 = 8'd145;
b_mant0 = 8'd202; b_mant1 = 8'd165; b_mant2 = 8'd185; b_mant3 = 8'd112;
a_exp0 = 10'd415; a_exp1 = 10'd340; a_exp2 = 10'd203; a_exp3 = 10'd798;
b_exp0 = 10'd721; b_exp1 = 10'd323; b_exp2 = 10'd52; b_exp3 = 10'd134;
a_sign0 = 4'd15; a_sign1 = 4'd16; a_sign2 = 4'd7; a_sign3 = 4'd2;
b_sign0 = 4'd8; b_sign1 = 4'd7; b_sign2 = 4'd16; b_sign3 = 4'd12;
@(posedge clk_i);
a_mant0 = 8'd140; a_mant1 = 8'd63; a_mant2 = 8'd9; a_mant3 = 8'd57;
b_mant0 = 8'd156; b_mant1 = 8'd4; b_mant2 = 8'd11; b_mant3 = 8'd189;
a_exp0 = 10'd141; a_exp1 = 10'd858; a_exp2 = 10'd560; a_exp3 = 10'd267;
b_exp0 = 10'd747; b_exp1 = 10'd649; b_exp2 = 10'd334; b_exp3 = 10'd979;
a_sign0 = 4'd15; a_sign1 = 4'd1; a_sign2 = 4'd5; a_sign3 = 4'd15;
b_sign0 = 4'd2; b_sign1 = 4'd15; b_sign2 = 4'd6; b_sign3 = 4'd6;
@(posedge clk_i);
a_mant0 = 8'd100; a_mant1 = 8'd143; a_mant2 = 8'd23; a_mant3 = 8'd206;
b_mant0 = 8'd14; b_mant1 = 8'd229; b_mant2 = 8'd30; b_mant3 = 8'd201;
a_exp0 = 10'd692; a_exp1 = 10'd742; a_exp2 = 10'd637; a_exp3 = 10'd917;
b_exp0 = 10'd1002; b_exp1 = 10'd552; b_exp2 = 10'd1020; b_exp3 = 10'd350;
a_sign0 = 4'd0; a_sign1 = 4'd16; a_sign2 = 4'd16; a_sign3 = 4'd1;
b_sign0 = 4'd11; b_sign1 = 4'd7; b_sign2 = 4'd13; b_sign3 = 4'd4;
@(posedge clk_i);
shared_exps0 = 8'd133;
shared_exps1 = 8'd114;
a_mant0 = 8'd108; a_mant1 = 8'd110; a_mant2 = 8'd144; a_mant3 = 8'd180;
b_mant0 = 8'd41; b_mant1 = 8'd166; b_mant2 = 8'd117; b_mant3 = 8'd78;
a_exp0 = 10'd566; a_exp1 = 10'd679; a_exp2 = 10'd374; a_exp3 = 10'd312;
b_exp0 = 10'd529; b_exp1 = 10'd337; b_exp2 = 10'd217; b_exp3 = 10'd45;
a_sign0 = 4'd6; a_sign1 = 4'd2; a_sign2 = 4'd1; a_sign3 = 4'd10;
b_sign0 = 4'd8; b_sign1 = 4'd15; b_sign2 = 4'd16; b_sign3 = 4'd1;
@(posedge clk_i);
a_mant0 = 8'd242; a_mant1 = 8'd229; a_mant2 = 8'd209; a_mant3 = 8'd223;
b_mant0 = 8'd196; b_mant1 = 8'd115; b_mant2 = 8'd252; b_mant3 = 8'd63;
a_exp0 = 10'd566; a_exp1 = 10'd794; a_exp2 = 10'd463; a_exp3 = 10'd14;
b_exp0 = 10'd14; b_exp1 = 10'd481; b_exp2 = 10'd553; b_exp3 = 10'd576;
a_sign0 = 4'd3; a_sign1 = 4'd8; a_sign2 = 4'd9; a_sign3 = 4'd0;
b_sign0 = 4'd7; b_sign1 = 4'd7; b_sign2 = 4'd12; b_sign3 = 4'd16;
@(posedge clk_i);
a_mant0 = 8'd57; a_mant1 = 8'd191; a_mant2 = 8'd194; a_mant3 = 8'd243;
b_mant0 = 8'd9; b_mant1 = 8'd61; b_mant2 = 8'd152; b_mant3 = 8'd27;
a_exp0 = 10'd781; a_exp1 = 10'd547; a_exp2 = 10'd262; a_exp3 = 10'd437;
b_exp0 = 10'd253; b_exp1 = 10'd628; b_exp2 = 10'd713; b_exp3 = 10'd349;
a_sign0 = 4'd16; a_sign1 = 4'd11; a_sign2 = 4'd14; a_sign3 = 4'd10;
b_sign0 = 4'd3; b_sign1 = 4'd2; b_sign2 = 4'd7; b_sign3 = 4'd2;
@(posedge clk_i);
a_mant0 = 8'd200; a_mant1 = 8'd53; a_mant2 = 8'd126; a_mant3 = 8'd106;
b_mant0 = 8'd230; b_mant1 = 8'd47; b_mant2 = 8'd162; b_mant3 = 8'd70;
a_exp0 = 10'd208; a_exp1 = 10'd14; a_exp2 = 10'd14; a_exp3 = 10'd249;
b_exp0 = 10'd271; b_exp1 = 10'd175; b_exp2 = 10'd166; b_exp3 = 10'd504;
a_sign0 = 4'd2; a_sign1 = 4'd5; a_sign2 = 4'd15; a_sign3 = 4'd2;
b_sign0 = 4'd3; b_sign1 = 4'd16; b_sign2 = 4'd12; b_sign3 = 4'd14;
@(posedge clk_i);
a_mant0 = 8'd195; a_mant1 = 8'd77; a_mant2 = 8'd109; a_mant3 = 8'd58;
b_mant0 = 8'd223; b_mant1 = 8'd51; b_mant2 = 8'd26; b_mant3 = 8'd51;
a_exp0 = 10'd514; a_exp1 = 10'd45; a_exp2 = 10'd467; a_exp3 = 10'd1014;
b_exp0 = 10'd368; b_exp1 = 10'd559; b_exp2 = 10'd510; b_exp3 = 10'd793;
a_sign0 = 4'd14; a_sign1 = 4'd12; a_sign2 = 4'd14; a_sign3 = 4'd10;
b_sign0 = 4'd8; b_sign1 = 4'd15; b_sign2 = 4'd6; b_sign3 = 4'd12;
@(posedge clk_i);
a_mant0 = 8'd149; a_mant1 = 8'd128; a_mant2 = 8'd36; a_mant3 = 8'd251;
b_mant0 = 8'd24; b_mant1 = 8'd243; b_mant2 = 8'd47; b_mant3 = 8'd81;
a_exp0 = 10'd453; a_exp1 = 10'd990; a_exp2 = 10'd528; a_exp3 = 10'd31;
b_exp0 = 10'd516; b_exp1 = 10'd432; b_exp2 = 10'd116; b_exp3 = 10'd532;
a_sign0 = 4'd16; a_sign1 = 4'd4; a_sign2 = 4'd8; a_sign3 = 4'd15;
b_sign0 = 4'd6; b_sign1 = 4'd8; b_sign2 = 4'd15; b_sign3 = 4'd8;
@(posedge clk_i);
a_mant0 = 8'd195; a_mant1 = 8'd229; a_mant2 = 8'd172; a_mant3 = 8'd142;
b_mant0 = 8'd84; b_mant1 = 8'd170; b_mant2 = 8'd173; b_mant3 = 8'd193;
a_exp0 = 10'd68; a_exp1 = 10'd428; a_exp2 = 10'd957; a_exp3 = 10'd839;
b_exp0 = 10'd308; b_exp1 = 10'd233; b_exp2 = 10'd805; b_exp3 = 10'd641;
a_sign0 = 4'd4; a_sign1 = 4'd1; a_sign2 = 4'd12; a_sign3 = 4'd8;
b_sign0 = 4'd14; b_sign1 = 4'd3; b_sign2 = 4'd7; b_sign3 = 4'd10;
@(posedge clk_i);
a_mant0 = 8'd31; a_mant1 = 8'd82; a_mant2 = 8'd199; a_mant3 = 8'd165;
b_mant0 = 8'd245; b_mant1 = 8'd69; b_mant2 = 8'd15; b_mant3 = 8'd106;
a_exp0 = 10'd930; a_exp1 = 10'd629; a_exp2 = 10'd806; a_exp3 = 10'd717;
b_exp0 = 10'd73; b_exp1 = 10'd761; b_exp2 = 10'd221; b_exp3 = 10'd5;
a_sign0 = 4'd8; a_sign1 = 4'd14; a_sign2 = 4'd12; a_sign3 = 4'd12;
b_sign0 = 4'd4; b_sign1 = 4'd12; b_sign2 = 4'd5; b_sign3 = 4'd1;
@(posedge clk_i);
shared_exps0 = 8'd117;
shared_exps1 = 8'd155;
a_mant0 = 8'd54; a_mant1 = 8'd115; a_mant2 = 8'd72; a_mant3 = 8'd158;
b_mant0 = 8'd74; b_mant1 = 8'd136; b_mant2 = 8'd155; b_mant3 = 8'd141;
a_exp0 = 10'd906; a_exp1 = 10'd352; a_exp2 = 10'd55; a_exp3 = 10'd554;
b_exp0 = 10'd996; b_exp1 = 10'd931; b_exp2 = 10'd453; b_exp3 = 10'd116;
a_sign0 = 4'd3; a_sign1 = 4'd5; a_sign2 = 4'd5; a_sign3 = 4'd13;
b_sign0 = 4'd11; b_sign1 = 4'd8; b_sign2 = 4'd15; b_sign3 = 4'd13;
@(posedge clk_i);
a_mant0 = 8'd115; a_mant1 = 8'd232; a_mant2 = 8'd122; a_mant3 = 8'd192;
b_mant0 = 8'd86; b_mant1 = 8'd210; b_mant2 = 8'd179; b_mant3 = 8'd79;
a_exp0 = 10'd113; a_exp1 = 10'd342; a_exp2 = 10'd399; a_exp3 = 10'd438;
b_exp0 = 10'd350; b_exp1 = 10'd367; b_exp2 = 10'd123; b_exp3 = 10'd295;
a_sign0 = 4'd13; a_sign1 = 4'd7; a_sign2 = 4'd6; a_sign3 = 4'd16;
b_sign0 = 4'd16; b_sign1 = 4'd4; b_sign2 = 4'd9; b_sign3 = 4'd6;
@(posedge clk_i);
a_mant0 = 8'd176; a_mant1 = 8'd91; a_mant2 = 8'd188; a_mant3 = 8'd119;
b_mant0 = 8'd35; b_mant1 = 8'd205; b_mant2 = 8'd129; b_mant3 = 8'd174;
a_exp0 = 10'd875; a_exp1 = 10'd24; a_exp2 = 10'd787; a_exp3 = 10'd955;
b_exp0 = 10'd932; b_exp1 = 10'd531; b_exp2 = 10'd474; b_exp3 = 10'd823;
a_sign0 = 4'd12; a_sign1 = 4'd5; a_sign2 = 4'd15; a_sign3 = 4'd0;
b_sign0 = 4'd1; b_sign1 = 4'd3; b_sign2 = 4'd8; b_sign3 = 4'd7;
@(posedge clk_i);
a_mant0 = 8'd229; a_mant1 = 8'd122; a_mant2 = 8'd117; a_mant3 = 8'd49;
b_mant0 = 8'd119; b_mant1 = 8'd194; b_mant2 = 8'd36; b_mant3 = 8'd211;
a_exp0 = 10'd280; a_exp1 = 10'd646; a_exp2 = 10'd860; a_exp3 = 10'd920;
b_exp0 = 10'd223; b_exp1 = 10'd976; b_exp2 = 10'd275; b_exp3 = 10'd46;
a_sign0 = 4'd1; a_sign1 = 4'd15; a_sign2 = 4'd8; a_sign3 = 4'd11;
b_sign0 = 4'd16; b_sign1 = 4'd9; b_sign2 = 4'd14; b_sign3 = 4'd11;
@(posedge clk_i);
a_mant0 = 8'd81; a_mant1 = 8'd236; a_mant2 = 8'd17; a_mant3 = 8'd113;
b_mant0 = 8'd53; b_mant1 = 8'd146; b_mant2 = 8'd4; b_mant3 = 8'd224;
a_exp0 = 10'd1013; a_exp1 = 10'd603; a_exp2 = 10'd203; a_exp3 = 10'd647;
b_exp0 = 10'd952; b_exp1 = 10'd806; b_exp2 = 10'd632; b_exp3 = 10'd770;
a_sign0 = 4'd1; a_sign1 = 4'd12; a_sign2 = 4'd0; a_sign3 = 4'd14;
b_sign0 = 4'd15; b_sign1 = 4'd13; b_sign2 = 4'd8; b_sign3 = 4'd16;
@(posedge clk_i);
a_mant0 = 8'd59; a_mant1 = 8'd165; a_mant2 = 8'd202; a_mant3 = 8'd215;
b_mant0 = 8'd71; b_mant1 = 8'd103; b_mant2 = 8'd237; b_mant3 = 8'd41;
a_exp0 = 10'd258; a_exp1 = 10'd437; a_exp2 = 10'd848; a_exp3 = 10'd446;
b_exp0 = 10'd915; b_exp1 = 10'd511; b_exp2 = 10'd854; b_exp3 = 10'd749;
a_sign0 = 4'd16; a_sign1 = 4'd9; a_sign2 = 4'd0; a_sign3 = 4'd14;
b_sign0 = 4'd14; b_sign1 = 4'd3; b_sign2 = 4'd8; b_sign3 = 4'd6;
@(posedge clk_i);
a_mant0 = 8'd35; a_mant1 = 8'd57; a_mant2 = 8'd105; a_mant3 = 8'd185;
b_mant0 = 8'd100; b_mant1 = 8'd8; b_mant2 = 8'd105; b_mant3 = 8'd111;
a_exp0 = 10'd107; a_exp1 = 10'd1004; a_exp2 = 10'd54; a_exp3 = 10'd607;
b_exp0 = 10'd668; b_exp1 = 10'd492; b_exp2 = 10'd183; b_exp3 = 10'd771;
a_sign0 = 4'd5; a_sign1 = 4'd3; a_sign2 = 4'd8; a_sign3 = 4'd1;
b_sign0 = 4'd12; b_sign1 = 4'd8; b_sign2 = 4'd1; b_sign3 = 4'd11;
@(posedge clk_i);
a_mant0 = 8'd242; a_mant1 = 8'd173; a_mant2 = 8'd149; a_mant3 = 8'd50;
b_mant0 = 8'd77; b_mant1 = 8'd152; b_mant2 = 8'd149; b_mant3 = 8'd207;
a_exp0 = 10'd154; a_exp1 = 10'd2; a_exp2 = 10'd453; a_exp3 = 10'd651;
b_exp0 = 10'd354; b_exp1 = 10'd620; b_exp2 = 10'd260; b_exp3 = 10'd214;
a_sign0 = 4'd8; a_sign1 = 4'd16; a_sign2 = 4'd16; a_sign3 = 4'd5;
b_sign0 = 4'd3; b_sign1 = 4'd12; b_sign2 = 4'd8; b_sign3 = 4'd13;
@(posedge clk_i);
shared_exps0 = 8'd122;
shared_exps1 = 8'd100;
a_mant0 = 8'd220; a_mant1 = 8'd215; a_mant2 = 8'd84; a_mant3 = 8'd206;
b_mant0 = 8'd52; b_mant1 = 8'd82; b_mant2 = 8'd37; b_mant3 = 8'd31;
a_exp0 = 10'd333; a_exp1 = 10'd637; a_exp2 = 10'd382; a_exp3 = 10'd200;
b_exp0 = 10'd306; b_exp1 = 10'd673; b_exp2 = 10'd727; b_exp3 = 10'd810;
a_sign0 = 4'd9; a_sign1 = 4'd11; a_sign2 = 4'd1; a_sign3 = 4'd16;
b_sign0 = 4'd14; b_sign1 = 4'd15; b_sign2 = 4'd14; b_sign3 = 4'd8;
@(posedge clk_i);
a_mant0 = 8'd208; a_mant1 = 8'd21; a_mant2 = 8'd200; a_mant3 = 8'd106;
b_mant0 = 8'd158; b_mant1 = 8'd121; b_mant2 = 8'd241; b_mant3 = 8'd125;
a_exp0 = 10'd945; a_exp1 = 10'd432; a_exp2 = 10'd150; a_exp3 = 10'd41;
b_exp0 = 10'd158; b_exp1 = 10'd585; b_exp2 = 10'd7; b_exp3 = 10'd752;
a_sign0 = 4'd12; a_sign1 = 4'd11; a_sign2 = 4'd4; a_sign3 = 4'd16;
b_sign0 = 4'd1; b_sign1 = 4'd11; b_sign2 = 4'd0; b_sign3 = 4'd16;
@(posedge clk_i);
a_mant0 = 8'd251; a_mant1 = 8'd130; a_mant2 = 8'd227; a_mant3 = 8'd234;
b_mant0 = 8'd73; b_mant1 = 8'd34; b_mant2 = 8'd45; b_mant3 = 8'd108;
a_exp0 = 10'd752; a_exp1 = 10'd401; a_exp2 = 10'd428; a_exp3 = 10'd963;
b_exp0 = 10'd747; b_exp1 = 10'd897; b_exp2 = 10'd963; b_exp3 = 10'd191;
a_sign0 = 4'd6; a_sign1 = 4'd11; a_sign2 = 4'd8; a_sign3 = 4'd15;
b_sign0 = 4'd9; b_sign1 = 4'd16; b_sign2 = 4'd13; b_sign3 = 4'd2;
@(posedge clk_i);
a_mant0 = 8'd167; a_mant1 = 8'd168; a_mant2 = 8'd174; a_mant3 = 8'd8;
b_mant0 = 8'd104; b_mant1 = 8'd201; b_mant2 = 8'd134; b_mant3 = 8'd255;
a_exp0 = 10'd205; a_exp1 = 10'd39; a_exp2 = 10'd482; a_exp3 = 10'd833;
b_exp0 = 10'd7; b_exp1 = 10'd338; b_exp2 = 10'd855; b_exp3 = 10'd1011;
a_sign0 = 4'd12; a_sign1 = 4'd9; a_sign2 = 4'd11; a_sign3 = 4'd1;
b_sign0 = 4'd11; b_sign1 = 4'd11; b_sign2 = 4'd3; b_sign3 = 4'd5;
@(posedge clk_i);
a_mant0 = 8'd106; a_mant1 = 8'd251; a_mant2 = 8'd215; a_mant3 = 8'd167;
b_mant0 = 8'd163; b_mant1 = 8'd177; b_mant2 = 8'd42; b_mant3 = 8'd52;
a_exp0 = 10'd894; a_exp1 = 10'd134; a_exp2 = 10'd464; a_exp3 = 10'd425;
b_exp0 = 10'd677; b_exp1 = 10'd142; b_exp2 = 10'd520; b_exp3 = 10'd972;
a_sign0 = 4'd9; a_sign1 = 4'd4; a_sign2 = 4'd5; a_sign3 = 4'd15;
b_sign0 = 4'd12; b_sign1 = 4'd8; b_sign2 = 4'd4; b_sign3 = 4'd11;
@(posedge clk_i);
a_mant0 = 8'd5; a_mant1 = 8'd53; a_mant2 = 8'd116; a_mant3 = 8'd50;
b_mant0 = 8'd97; b_mant1 = 8'd159; b_mant2 = 8'd219; b_mant3 = 8'd1;
a_exp0 = 10'd989; a_exp1 = 10'd688; a_exp2 = 10'd820; a_exp3 = 10'd582;
b_exp0 = 10'd498; b_exp1 = 10'd928; b_exp2 = 10'd77; b_exp3 = 10'd499;
a_sign0 = 4'd4; a_sign1 = 4'd14; a_sign2 = 4'd14; a_sign3 = 4'd11;
b_sign0 = 4'd8; b_sign1 = 4'd1; b_sign2 = 4'd14; b_sign3 = 4'd8;
@(posedge clk_i);
a_mant0 = 8'd172; a_mant1 = 8'd244; a_mant2 = 8'd206; a_mant3 = 8'd134;
b_mant0 = 8'd125; b_mant1 = 8'd20; b_mant2 = 8'd189; b_mant3 = 8'd190;
a_exp0 = 10'd140; a_exp1 = 10'd225; a_exp2 = 10'd48; a_exp3 = 10'd743;
b_exp0 = 10'd70; b_exp1 = 10'd648; b_exp2 = 10'd668; b_exp3 = 10'd601;
a_sign0 = 4'd16; a_sign1 = 4'd2; a_sign2 = 4'd4; a_sign3 = 4'd15;
b_sign0 = 4'd3; b_sign1 = 4'd9; b_sign2 = 4'd14; b_sign3 = 4'd0;
@(posedge clk_i);
a_mant0 = 8'd148; a_mant1 = 8'd34; a_mant2 = 8'd162; a_mant3 = 8'd186;
b_mant0 = 8'd97; b_mant1 = 8'd113; b_mant2 = 8'd1; b_mant3 = 8'd98;
a_exp0 = 10'd751; a_exp1 = 10'd452; a_exp2 = 10'd47; a_exp3 = 10'd1006;
b_exp0 = 10'd480; b_exp1 = 10'd436; b_exp2 = 10'd778; b_exp3 = 10'd463;
a_sign0 = 4'd12; a_sign1 = 4'd10; a_sign2 = 4'd12; a_sign3 = 4'd9;
b_sign0 = 4'd2; b_sign1 = 4'd10; b_sign2 = 4'd15; b_sign3 = 4'd15;
@(posedge clk_i);
shared_exps0 = 8'd165;
shared_exps1 = 8'd119;
rstn = 0;
@(posedge clk_i);
rstn = 1;
a_mant0 = 8'd45; a_mant1 = 8'd238; a_mant2 = 8'd116; a_mant3 = 8'd122;
b_mant0 = 8'd93; b_mant1 = 8'd19; b_mant2 = 8'd118; b_mant3 = 8'd77;
a_exp0 = 10'd900; a_exp1 = 10'd104; a_exp2 = 10'd70; a_exp3 = 10'd157;
b_exp0 = 10'd182; b_exp1 = 10'd429; b_exp2 = 10'd89; b_exp3 = 10'd424;
a_sign0 = 4'd6; a_sign1 = 4'd0; a_sign2 = 4'd12; a_sign3 = 4'd14;
b_sign0 = 4'd8; b_sign1 = 4'd3; b_sign2 = 4'd8; b_sign3 = 4'd12;
@(posedge clk_i);
a_mant0 = 8'd151; a_mant1 = 8'd193; a_mant2 = 8'd200; a_mant3 = 8'd185;
b_mant0 = 8'd90; b_mant1 = 8'd50; b_mant2 = 8'd89; b_mant3 = 8'd104;
a_exp0 = 10'd157; a_exp1 = 10'd987; a_exp2 = 10'd290; a_exp3 = 10'd319;
b_exp0 = 10'd154; b_exp1 = 10'd178; b_exp2 = 10'd342; b_exp3 = 10'd211;
a_sign0 = 4'd16; a_sign1 = 4'd7; a_sign2 = 4'd10; a_sign3 = 4'd1;
b_sign0 = 4'd16; b_sign1 = 4'd8; b_sign2 = 4'd11; b_sign3 = 4'd9;
@(posedge clk_i);
a_mant0 = 8'd97; a_mant1 = 8'd46; a_mant2 = 8'd236; a_mant3 = 8'd136;
b_mant0 = 8'd217; b_mant1 = 8'd99; b_mant2 = 8'd185; b_mant3 = 8'd0;
a_exp0 = 10'd575; a_exp1 = 10'd645; a_exp2 = 10'd446; a_exp3 = 10'd157;
b_exp0 = 10'd754; b_exp1 = 10'd822; b_exp2 = 10'd895; b_exp3 = 10'd972;
a_sign0 = 4'd3; a_sign1 = 4'd12; a_sign2 = 4'd11; a_sign3 = 4'd14;
b_sign0 = 4'd4; b_sign1 = 4'd5; b_sign2 = 4'd9; b_sign3 = 4'd6;
@(posedge clk_i);
a_mant0 = 8'd231; a_mant1 = 8'd219; a_mant2 = 8'd118; a_mant3 = 8'd221;
b_mant0 = 8'd61; b_mant1 = 8'd67; b_mant2 = 8'd184; b_mant3 = 8'd108;
a_exp0 = 10'd409; a_exp1 = 10'd300; a_exp2 = 10'd524; a_exp3 = 10'd571;
b_exp0 = 10'd473; b_exp1 = 10'd337; b_exp2 = 10'd1019; b_exp3 = 10'd384;
a_sign0 = 4'd13; a_sign1 = 4'd8; a_sign2 = 4'd3; a_sign3 = 4'd9;
b_sign0 = 4'd2; b_sign1 = 4'd2; b_sign2 = 4'd7; b_sign3 = 4'd15;
@(posedge clk_i);
a_mant0 = 8'd237; a_mant1 = 8'd87; a_mant2 = 8'd148; a_mant3 = 8'd1;
b_mant0 = 8'd111; b_mant1 = 8'd155; b_mant2 = 8'd203; b_mant3 = 8'd3;
a_exp0 = 10'd799; a_exp1 = 10'd798; a_exp2 = 10'd381; a_exp3 = 10'd762;
b_exp0 = 10'd478; b_exp1 = 10'd227; b_exp2 = 10'd313; b_exp3 = 10'd869;
a_sign0 = 4'd5; a_sign1 = 4'd8; a_sign2 = 4'd15; a_sign3 = 4'd9;
b_sign0 = 4'd11; b_sign1 = 4'd10; b_sign2 = 4'd9; b_sign3 = 4'd0;
@(posedge clk_i);
a_mant0 = 8'd207; a_mant1 = 8'd79; a_mant2 = 8'd185; a_mant3 = 8'd190;
b_mant0 = 8'd193; b_mant1 = 8'd43; b_mant2 = 8'd157; b_mant3 = 8'd12;
a_exp0 = 10'd348; a_exp1 = 10'd736; a_exp2 = 10'd464; a_exp3 = 10'd767;
b_exp0 = 10'd641; b_exp1 = 10'd867; b_exp2 = 10'd259; b_exp3 = 10'd857;
a_sign0 = 4'd12; a_sign1 = 4'd0; a_sign2 = 4'd10; a_sign3 = 4'd9;
b_sign0 = 4'd11; b_sign1 = 4'd3; b_sign2 = 4'd11; b_sign3 = 4'd13;
@(posedge clk_i);
a_mant0 = 8'd251; a_mant1 = 8'd162; a_mant2 = 8'd71; a_mant3 = 8'd149;
b_mant0 = 8'd114; b_mant1 = 8'd42; b_mant2 = 8'd211; b_mant3 = 8'd45;
a_exp0 = 10'd910; a_exp1 = 10'd596; a_exp2 = 10'd624; a_exp3 = 10'd18;
b_exp0 = 10'd440; b_exp1 = 10'd259; b_exp2 = 10'd92; b_exp3 = 10'd669;
a_sign0 = 4'd14; a_sign1 = 4'd3; a_sign2 = 4'd7; a_sign3 = 4'd6;
b_sign0 = 4'd0; b_sign1 = 4'd7; b_sign2 = 4'd4; b_sign3 = 4'd3;
@(posedge clk_i);
shared_exps0 = 8'd115;
shared_exps1 = 8'd101;
a_mant0 = 8'd68; a_mant1 = 8'd239; a_mant2 = 8'd96; a_mant3 = 8'd218;
b_mant0 = 8'd93; b_mant1 = 8'd30; b_mant2 = 8'd21; b_mant3 = 8'd255;
a_exp0 = 10'd886; a_exp1 = 10'd39; a_exp2 = 10'd835; a_exp3 = 10'd269;
b_exp0 = 10'd285; b_exp1 = 10'd848; b_exp2 = 10'd243; b_exp3 = 10'd210;
a_sign0 = 4'd11; a_sign1 = 4'd8; a_sign2 = 4'd15; a_sign3 = 4'd13;
b_sign0 = 4'd2; b_sign1 = 4'd6; b_sign2 = 4'd14; b_sign3 = 4'd0;
@(posedge clk_i);
a_mant0 = 8'd138; a_mant1 = 8'd205; a_mant2 = 8'd220; a_mant3 = 8'd239;
b_mant0 = 8'd108; b_mant1 = 8'd238; b_mant2 = 8'd96; b_mant3 = 8'd245;
a_exp0 = 10'd746; a_exp1 = 10'd134; a_exp2 = 10'd602; a_exp3 = 10'd167;
b_exp0 = 10'd791; b_exp1 = 10'd380; b_exp2 = 10'd680; b_exp3 = 10'd470;
a_sign0 = 4'd11; a_sign1 = 4'd14; a_sign2 = 4'd9; a_sign3 = 4'd1;
b_sign0 = 4'd12; b_sign1 = 4'd0; b_sign2 = 4'd14; b_sign3 = 4'd9;
@(posedge clk_i);
a_mant0 = 8'd210; a_mant1 = 8'd3; a_mant2 = 8'd33; a_mant3 = 8'd34;
b_mant0 = 8'd123; b_mant1 = 8'd57; b_mant2 = 8'd28; b_mant3 = 8'd207;
a_exp0 = 10'd41; a_exp1 = 10'd526; a_exp2 = 10'd73; a_exp3 = 10'd626;
b_exp0 = 10'd270; b_exp1 = 10'd234; b_exp2 = 10'd122; b_exp3 = 10'd101;
a_sign0 = 4'd6; a_sign1 = 4'd1; a_sign2 = 4'd16; a_sign3 = 4'd3;
b_sign0 = 4'd16; b_sign1 = 4'd8; b_sign2 = 4'd9; b_sign3 = 4'd0;
@(posedge clk_i);
a_mant0 = 8'd36; a_mant1 = 8'd12; a_mant2 = 8'd203; a_mant3 = 8'd238;
b_mant0 = 8'd215; b_mant1 = 8'd139; b_mant2 = 8'd51; b_mant3 = 8'd108;
a_exp0 = 10'd925; a_exp1 = 10'd528; a_exp2 = 10'd514; a_exp3 = 10'd380;
b_exp0 = 10'd347; b_exp1 = 10'd902; b_exp2 = 10'd127; b_exp3 = 10'd769;
a_sign0 = 4'd13; a_sign1 = 4'd14; a_sign2 = 4'd6; a_sign3 = 4'd16;
b_sign0 = 4'd5; b_sign1 = 4'd2; b_sign2 = 4'd9; b_sign3 = 4'd9;
@(posedge clk_i);
a_mant0 = 8'd44; a_mant1 = 8'd221; a_mant2 = 8'd48; a_mant3 = 8'd225;
b_mant0 = 8'd85; b_mant1 = 8'd57; b_mant2 = 8'd103; b_mant3 = 8'd129;
a_exp0 = 10'd569; a_exp1 = 10'd842; a_exp2 = 10'd930; a_exp3 = 10'd457;
b_exp0 = 10'd241; b_exp1 = 10'd460; b_exp2 = 10'd216; b_exp3 = 10'd572;
a_sign0 = 4'd13; a_sign1 = 4'd14; a_sign2 = 4'd4; a_sign3 = 4'd0;
b_sign0 = 4'd12; b_sign1 = 4'd9; b_sign2 = 4'd7; b_sign3 = 4'd11;
@(posedge clk_i);
a_mant0 = 8'd193; a_mant1 = 8'd187; a_mant2 = 8'd208; a_mant3 = 8'd95;
b_mant0 = 8'd223; b_mant1 = 8'd146; b_mant2 = 8'd54; b_mant3 = 8'd36;
a_exp0 = 10'd239; a_exp1 = 10'd936; a_exp2 = 10'd845; a_exp3 = 10'd708;
b_exp0 = 10'd969; b_exp1 = 10'd834; b_exp2 = 10'd802; b_exp3 = 10'd269;
a_sign0 = 4'd7; a_sign1 = 4'd3; a_sign2 = 4'd7; a_sign3 = 4'd11;
b_sign0 = 4'd2; b_sign1 = 4'd3; b_sign2 = 4'd1; b_sign3 = 4'd1;
@(posedge clk_i);
a_mant0 = 8'd178; a_mant1 = 8'd242; a_mant2 = 8'd17; a_mant3 = 8'd29;
b_mant0 = 8'd157; b_mant1 = 8'd80; b_mant2 = 8'd158; b_mant3 = 8'd129;
a_exp0 = 10'd347; a_exp1 = 10'd936; a_exp2 = 10'd668; a_exp3 = 10'd534;
b_exp0 = 10'd422; b_exp1 = 10'd548; b_exp2 = 10'd241; b_exp3 = 10'd312;
a_sign0 = 4'd14; a_sign1 = 4'd4; a_sign2 = 4'd1; a_sign3 = 4'd9;
b_sign0 = 4'd1; b_sign1 = 4'd3; b_sign2 = 4'd2; b_sign3 = 4'd0;
@(posedge clk_i);
a_mant0 = 8'd240; a_mant1 = 8'd91; a_mant2 = 8'd236; a_mant3 = 8'd52;
b_mant0 = 8'd201; b_mant1 = 8'd252; b_mant2 = 8'd166; b_mant3 = 8'd140;
a_exp0 = 10'd311; a_exp1 = 10'd109; a_exp2 = 10'd161; a_exp3 = 10'd277;
b_exp0 = 10'd3; b_exp1 = 10'd470; b_exp2 = 10'd835; b_exp3 = 10'd624;
a_sign0 = 4'd2; a_sign1 = 4'd3; a_sign2 = 4'd11; a_sign3 = 4'd5;
b_sign0 = 4'd1; b_sign1 = 4'd3; b_sign2 = 4'd0; b_sign3 = 4'd7;
@(posedge clk_i);
shared_exps0 = 8'd123;
shared_exps1 = 8'd137;
a_mant0 = 8'd23; a_mant1 = 8'd59; a_mant2 = 8'd1; a_mant3 = 8'd200;
b_mant0 = 8'd69; b_mant1 = 8'd24; b_mant2 = 8'd47; b_mant3 = 8'd200;
a_exp0 = 10'd103; a_exp1 = 10'd604; a_exp2 = 10'd39; a_exp3 = 10'd837;
b_exp0 = 10'd964; b_exp1 = 10'd235; b_exp2 = 10'd240; b_exp3 = 10'd773;
a_sign0 = 4'd9; a_sign1 = 4'd4; a_sign2 = 4'd1; a_sign3 = 4'd11;
b_sign0 = 4'd14; b_sign1 = 4'd1; b_sign2 = 4'd1; b_sign3 = 4'd15;
@(posedge clk_i);
a_mant0 = 8'd248; a_mant1 = 8'd122; a_mant2 = 8'd216; a_mant3 = 8'd157;
b_mant0 = 8'd120; b_mant1 = 8'd224; b_mant2 = 8'd56; b_mant3 = 8'd15;
a_exp0 = 10'd639; a_exp1 = 10'd297; a_exp2 = 10'd266; a_exp3 = 10'd601;
b_exp0 = 10'd172; b_exp1 = 10'd892; b_exp2 = 10'd52; b_exp3 = 10'd198;
a_sign0 = 4'd7; a_sign1 = 4'd8; a_sign2 = 4'd3; a_sign3 = 4'd13;
b_sign0 = 4'd0; b_sign1 = 4'd15; b_sign2 = 4'd16; b_sign3 = 4'd1;
@(posedge clk_i);
a_mant0 = 8'd16; a_mant1 = 8'd105; a_mant2 = 8'd27; a_mant3 = 8'd70;
b_mant0 = 8'd246; b_mant1 = 8'd228; b_mant2 = 8'd192; b_mant3 = 8'd53;
a_exp0 = 10'd994; a_exp1 = 10'd749; a_exp2 = 10'd61; a_exp3 = 10'd45;
b_exp0 = 10'd963; b_exp1 = 10'd803; b_exp2 = 10'd82; b_exp3 = 10'd58;
a_sign0 = 4'd14; a_sign1 = 4'd14; a_sign2 = 4'd3; a_sign3 = 4'd13;
b_sign0 = 4'd16; b_sign1 = 4'd2; b_sign2 = 4'd8; b_sign3 = 4'd0;
@(posedge clk_i);
a_mant0 = 8'd84; a_mant1 = 8'd249; a_mant2 = 8'd42; a_mant3 = 8'd13;
b_mant0 = 8'd190; b_mant1 = 8'd106; b_mant2 = 8'd147; b_mant3 = 8'd55;
a_exp0 = 10'd306; a_exp1 = 10'd97; a_exp2 = 10'd511; a_exp3 = 10'd80;
b_exp0 = 10'd802; b_exp1 = 10'd783; b_exp2 = 10'd917; b_exp3 = 10'd432;
a_sign0 = 4'd13; a_sign1 = 4'd4; a_sign2 = 4'd14; a_sign3 = 4'd14;
b_sign0 = 4'd14; b_sign1 = 4'd14; b_sign2 = 4'd9; b_sign3 = 4'd12;
@(posedge clk_i);
a_mant0 = 8'd201; a_mant1 = 8'd248; a_mant2 = 8'd94; a_mant3 = 8'd102;
b_mant0 = 8'd171; b_mant1 = 8'd162; b_mant2 = 8'd86; b_mant3 = 8'd233;
a_exp0 = 10'd816; a_exp1 = 10'd309; a_exp2 = 10'd888; a_exp3 = 10'd607;
b_exp0 = 10'd902; b_exp1 = 10'd46; b_exp2 = 10'd154; b_exp3 = 10'd73;
a_sign0 = 4'd14; a_sign1 = 4'd16; a_sign2 = 4'd8; a_sign3 = 4'd5;
b_sign0 = 4'd15; b_sign1 = 4'd14; b_sign2 = 4'd12; b_sign3 = 4'd11;
@(posedge clk_i);
a_mant0 = 8'd76; a_mant1 = 8'd0; a_mant2 = 8'd187; a_mant3 = 8'd100;
b_mant0 = 8'd200; b_mant1 = 8'd122; b_mant2 = 8'd96; b_mant3 = 8'd127;
a_exp0 = 10'd875; a_exp1 = 10'd944; a_exp2 = 10'd690; a_exp3 = 10'd638;
b_exp0 = 10'd845; b_exp1 = 10'd14; b_exp2 = 10'd899; b_exp3 = 10'd466;
a_sign0 = 4'd14; a_sign1 = 4'd1; a_sign2 = 4'd14; a_sign3 = 4'd12;
b_sign0 = 4'd13; b_sign1 = 4'd5; b_sign2 = 4'd12; b_sign3 = 4'd7;
@(posedge clk_i);
a_mant0 = 8'd37; a_mant1 = 8'd206; a_mant2 = 8'd199; a_mant3 = 8'd151;
b_mant0 = 8'd130; b_mant1 = 8'd82; b_mant2 = 8'd180; b_mant3 = 8'd228;
a_exp0 = 10'd468; a_exp1 = 10'd578; a_exp2 = 10'd469; a_exp3 = 10'd357;
b_exp0 = 10'd457; b_exp1 = 10'd642; b_exp2 = 10'd967; b_exp3 = 10'd982;
a_sign0 = 4'd11; a_sign1 = 4'd15; a_sign2 = 4'd13; a_sign3 = 4'd6;
b_sign0 = 4'd15; b_sign1 = 4'd2; b_sign2 = 4'd14; b_sign3 = 4'd1;
@(posedge clk_i);
a_mant0 = 8'd154; a_mant1 = 8'd163; a_mant2 = 8'd0; a_mant3 = 8'd167;
b_mant0 = 8'd56; b_mant1 = 8'd103; b_mant2 = 8'd23; b_mant3 = 8'd139;
a_exp0 = 10'd300; a_exp1 = 10'd593; a_exp2 = 10'd13; a_exp3 = 10'd799;
b_exp0 = 10'd390; b_exp1 = 10'd174; b_exp2 = 10'd535; b_exp3 = 10'd28;
a_sign0 = 4'd0; a_sign1 = 4'd12; a_sign2 = 4'd14; a_sign3 = 4'd4;
b_sign0 = 4'd4; b_sign1 = 4'd9; b_sign2 = 4'd7; b_sign3 = 4'd16;
@(posedge clk_i);
shared_exps0 = 8'd119;
shared_exps1 = 8'd112;
a_mant0 = 8'd146; a_mant1 = 8'd121; a_mant2 = 8'd126; a_mant3 = 8'd197;
b_mant0 = 8'd32; b_mant1 = 8'd184; b_mant2 = 8'd113; b_mant3 = 8'd247;
a_exp0 = 10'd146; a_exp1 = 10'd931; a_exp2 = 10'd275; a_exp3 = 10'd226;
b_exp0 = 10'd198; b_exp1 = 10'd846; b_exp2 = 10'd269; b_exp3 = 10'd745;
a_sign0 = 4'd9; a_sign1 = 4'd5; a_sign2 = 4'd9; a_sign3 = 4'd6;
b_sign0 = 4'd0; b_sign1 = 4'd0; b_sign2 = 4'd10; b_sign3 = 4'd15;
@(posedge clk_i);
a_mant0 = 8'd75; a_mant1 = 8'd183; a_mant2 = 8'd158; a_mant3 = 8'd194;
b_mant0 = 8'd84; b_mant1 = 8'd99; b_mant2 = 8'd38; b_mant3 = 8'd250;
a_exp0 = 10'd89; a_exp1 = 10'd491; a_exp2 = 10'd688; a_exp3 = 10'd57;
b_exp0 = 10'd347; b_exp1 = 10'd854; b_exp2 = 10'd1010; b_exp3 = 10'd441;
a_sign0 = 4'd8; a_sign1 = 4'd1; a_sign2 = 4'd6; a_sign3 = 4'd3;
b_sign0 = 4'd11; b_sign1 = 4'd9; b_sign2 = 4'd12; b_sign3 = 4'd6;
@(posedge clk_i);
a_mant0 = 8'd182; a_mant1 = 8'd228; a_mant2 = 8'd61; a_mant3 = 8'd104;
b_mant0 = 8'd97; b_mant1 = 8'd121; b_mant2 = 8'd36; b_mant3 = 8'd136;
a_exp0 = 10'd379; a_exp1 = 10'd778; a_exp2 = 10'd847; a_exp3 = 10'd13;
b_exp0 = 10'd414; b_exp1 = 10'd840; b_exp2 = 10'd458; b_exp3 = 10'd869;
a_sign0 = 4'd11; a_sign1 = 4'd5; a_sign2 = 4'd13; a_sign3 = 4'd15;
b_sign0 = 4'd9; b_sign1 = 4'd2; b_sign2 = 4'd11; b_sign3 = 4'd10;
@(posedge clk_i);
a_mant0 = 8'd248; a_mant1 = 8'd190; a_mant2 = 8'd86; a_mant3 = 8'd245;
b_mant0 = 8'd201; b_mant1 = 8'd219; b_mant2 = 8'd143; b_mant3 = 8'd220;
a_exp0 = 10'd928; a_exp1 = 10'd222; a_exp2 = 10'd125; a_exp3 = 10'd475;
b_exp0 = 10'd78; b_exp1 = 10'd762; b_exp2 = 10'd295; b_exp3 = 10'd299;
a_sign0 = 4'd10; a_sign1 = 4'd5; a_sign2 = 4'd5; a_sign3 = 4'd8;
b_sign0 = 4'd10; b_sign1 = 4'd14; b_sign2 = 4'd4; b_sign3 = 4'd9;
@(posedge clk_i);
a_mant0 = 8'd246; a_mant1 = 8'd113; a_mant2 = 8'd46; a_mant3 = 8'd94;
b_mant0 = 8'd1; b_mant1 = 8'd172; b_mant2 = 8'd236; b_mant3 = 8'd58;
a_exp0 = 10'd600; a_exp1 = 10'd322; a_exp2 = 10'd548; a_exp3 = 10'd465;
b_exp0 = 10'd370; b_exp1 = 10'd693; b_exp2 = 10'd715; b_exp3 = 10'd666;
a_sign0 = 4'd10; a_sign1 = 4'd15; a_sign2 = 4'd13; a_sign3 = 4'd8;
b_sign0 = 4'd8; b_sign1 = 4'd4; b_sign2 = 4'd1; b_sign3 = 4'd14;
@(posedge clk_i);
a_mant0 = 8'd65; a_mant1 = 8'd204; a_mant2 = 8'd17; a_mant3 = 8'd102;
b_mant0 = 8'd120; b_mant1 = 8'd114; b_mant2 = 8'd238; b_mant3 = 8'd57;
a_exp0 = 10'd338; a_exp1 = 10'd339; a_exp2 = 10'd505; a_exp3 = 10'd399;
b_exp0 = 10'd909; b_exp1 = 10'd311; b_exp2 = 10'd469; b_exp3 = 10'd614;
a_sign0 = 4'd6; a_sign1 = 4'd6; a_sign2 = 4'd14; a_sign3 = 4'd3;
b_sign0 = 4'd8; b_sign1 = 4'd10; b_sign2 = 4'd3; b_sign3 = 4'd1;
@(posedge clk_i);
a_mant0 = 8'd86; a_mant1 = 8'd87; a_mant2 = 8'd212; a_mant3 = 8'd102;
b_mant0 = 8'd93; b_mant1 = 8'd55; b_mant2 = 8'd71; b_mant3 = 8'd166;
a_exp0 = 10'd552; a_exp1 = 10'd572; a_exp2 = 10'd771; a_exp3 = 10'd395;
b_exp0 = 10'd269; b_exp1 = 10'd31; b_exp2 = 10'd741; b_exp3 = 10'd106;
a_sign0 = 4'd7; a_sign1 = 4'd10; a_sign2 = 4'd2; a_sign3 = 4'd13;
b_sign0 = 4'd7; b_sign1 = 4'd9; b_sign2 = 4'd14; b_sign3 = 4'd3;
@(posedge clk_i);
a_mant0 = 8'd121; a_mant1 = 8'd76; a_mant2 = 8'd81; a_mant3 = 8'd26;
b_mant0 = 8'd213; b_mant1 = 8'd87; b_mant2 = 8'd187; b_mant3 = 8'd125;
a_exp0 = 10'd774; a_exp1 = 10'd261; a_exp2 = 10'd183; a_exp3 = 10'd233;
b_exp0 = 10'd408; b_exp1 = 10'd913; b_exp2 = 10'd64; b_exp3 = 10'd826;
a_sign0 = 4'd11; a_sign1 = 4'd5; a_sign2 = 4'd11; a_sign3 = 4'd11;
b_sign0 = 4'd13; b_sign1 = 4'd0; b_sign2 = 4'd10; b_sign3 = 4'd5;
@(posedge clk_i);
shared_exps0 = 8'd134;
shared_exps1 = 8'd106;
rstn = 0;
@(posedge clk_i);
rstn = 1;
a_mant0 = 8'd234; a_mant1 = 8'd52; a_mant2 = 8'd84; a_mant3 = 8'd165;
b_mant0 = 8'd157; b_mant1 = 8'd155; b_mant2 = 8'd212; b_mant3 = 8'd206;
a_exp0 = 10'd486; a_exp1 = 10'd907; a_exp2 = 10'd970; a_exp3 = 10'd214;
b_exp0 = 10'd50; b_exp1 = 10'd552; b_exp2 = 10'd857; b_exp3 = 10'd472;
a_sign0 = 4'd4; a_sign1 = 4'd7; a_sign2 = 4'd11; a_sign3 = 4'd10;
b_sign0 = 4'd2; b_sign1 = 4'd14; b_sign2 = 4'd14; b_sign3 = 4'd2;
@(posedge clk_i);
a_mant0 = 8'd227; a_mant1 = 8'd227; a_mant2 = 8'd56; a_mant3 = 8'd30;
b_mant0 = 8'd179; b_mant1 = 8'd18; b_mant2 = 8'd242; b_mant3 = 8'd202;
a_exp0 = 10'd562; a_exp1 = 10'd944; a_exp2 = 10'd941; a_exp3 = 10'd409;
b_exp0 = 10'd519; b_exp1 = 10'd396; b_exp2 = 10'd782; b_exp3 = 10'd1014;
a_sign0 = 4'd0; a_sign1 = 4'd12; a_sign2 = 4'd14; a_sign3 = 4'd0;
b_sign0 = 4'd4; b_sign1 = 4'd10; b_sign2 = 4'd7; b_sign3 = 4'd16;
@(posedge clk_i);
a_mant0 = 8'd26; a_mant1 = 8'd61; a_mant2 = 8'd206; a_mant3 = 8'd109;
b_mant0 = 8'd244; b_mant1 = 8'd64; b_mant2 = 8'd163; b_mant3 = 8'd20;
a_exp0 = 10'd4; a_exp1 = 10'd7; a_exp2 = 10'd566; a_exp3 = 10'd875;
b_exp0 = 10'd768; b_exp1 = 10'd790; b_exp2 = 10'd228; b_exp3 = 10'd587;
a_sign0 = 4'd4; a_sign1 = 4'd0; a_sign2 = 4'd9; a_sign3 = 4'd9;
b_sign0 = 4'd4; b_sign1 = 4'd15; b_sign2 = 4'd1; b_sign3 = 4'd7;
@(posedge clk_i);
a_mant0 = 8'd175; a_mant1 = 8'd126; a_mant2 = 8'd30; a_mant3 = 8'd22;
b_mant0 = 8'd30; b_mant1 = 8'd150; b_mant2 = 8'd35; b_mant3 = 8'd33;
a_exp0 = 10'd223; a_exp1 = 10'd459; a_exp2 = 10'd13; a_exp3 = 10'd396;
b_exp0 = 10'd259; b_exp1 = 10'd389; b_exp2 = 10'd173; b_exp3 = 10'd796;
a_sign0 = 4'd7; a_sign1 = 4'd2; a_sign2 = 4'd4; a_sign3 = 4'd1;
b_sign0 = 4'd1; b_sign1 = 4'd11; b_sign2 = 4'd0; b_sign3 = 4'd16;
@(posedge clk_i);
a_mant0 = 8'd3; a_mant1 = 8'd150; a_mant2 = 8'd175; a_mant3 = 8'd171;
b_mant0 = 8'd249; b_mant1 = 8'd203; b_mant2 = 8'd125; b_mant3 = 8'd216;
a_exp0 = 10'd305; a_exp1 = 10'd663; a_exp2 = 10'd836; a_exp3 = 10'd288;
b_exp0 = 10'd99; b_exp1 = 10'd197; b_exp2 = 10'd918; b_exp3 = 10'd29;
a_sign0 = 4'd4; a_sign1 = 4'd5; a_sign2 = 4'd8; a_sign3 = 4'd13;
b_sign0 = 4'd1; b_sign1 = 4'd1; b_sign2 = 4'd11; b_sign3 = 4'd9;
@(posedge clk_i);
a_mant0 = 8'd23; a_mant1 = 8'd48; a_mant2 = 8'd123; a_mant3 = 8'd186;
b_mant0 = 8'd207; b_mant1 = 8'd42; b_mant2 = 8'd130; b_mant3 = 8'd74;
a_exp0 = 10'd1007; a_exp1 = 10'd580; a_exp2 = 10'd812; a_exp3 = 10'd36;
b_exp0 = 10'd396; b_exp1 = 10'd789; b_exp2 = 10'd125; b_exp3 = 10'd968;
a_sign0 = 4'd5; a_sign1 = 4'd9; a_sign2 = 4'd10; a_sign3 = 4'd12;
b_sign0 = 4'd10; b_sign1 = 4'd1; b_sign2 = 4'd12; b_sign3 = 4'd16;
@(posedge clk_i);
a_mant0 = 8'd57; a_mant1 = 8'd139; a_mant2 = 8'd19; a_mant3 = 8'd14;
b_mant0 = 8'd133; b_mant1 = 8'd72; b_mant2 = 8'd254; b_mant3 = 8'd37;
a_exp0 = 10'd53; a_exp1 = 10'd544; a_exp2 = 10'd760; a_exp3 = 10'd353;
b_exp0 = 10'd660; b_exp1 = 10'd523; b_exp2 = 10'd693; b_exp3 = 10'd991;
a_sign0 = 4'd15; a_sign1 = 4'd12; a_sign2 = 4'd16; a_sign3 = 4'd8;
b_sign0 = 4'd1; b_sign1 = 4'd2; b_sign2 = 4'd5; b_sign3 = 4'd0;
@(posedge clk_i);
shared_exps0 = 8'd134;
shared_exps1 = 8'd98;
a_mant0 = 8'd235; a_mant1 = 8'd135; a_mant2 = 8'd52; a_mant3 = 8'd241;
b_mant0 = 8'd102; b_mant1 = 8'd19; b_mant2 = 8'd60; b_mant3 = 8'd210;
a_exp0 = 10'd896; a_exp1 = 10'd1021; a_exp2 = 10'd638; a_exp3 = 10'd43;
b_exp0 = 10'd269; b_exp1 = 10'd729; b_exp2 = 10'd563; b_exp3 = 10'd393;
a_sign0 = 4'd8; a_sign1 = 4'd7; a_sign2 = 4'd15; a_sign3 = 4'd3;
b_sign0 = 4'd16; b_sign1 = 4'd9; b_sign2 = 4'd8; b_sign3 = 4'd11;
@(posedge clk_i);
a_mant0 = 8'd117; a_mant1 = 8'd7; a_mant2 = 8'd126; a_mant3 = 8'd181;
b_mant0 = 8'd206; b_mant1 = 8'd28; b_mant2 = 8'd234; b_mant3 = 8'd34;
a_exp0 = 10'd395; a_exp1 = 10'd720; a_exp2 = 10'd961; a_exp3 = 10'd456;
b_exp0 = 10'd844; b_exp1 = 10'd469; b_exp2 = 10'd825; b_exp3 = 10'd340;
a_sign0 = 4'd14; a_sign1 = 4'd15; a_sign2 = 4'd16; a_sign3 = 4'd10;
b_sign0 = 4'd5; b_sign1 = 4'd15; b_sign2 = 4'd10; b_sign3 = 4'd6;
@(posedge clk_i);
a_mant0 = 8'd46; a_mant1 = 8'd144; a_mant2 = 8'd203; a_mant3 = 8'd135;
b_mant0 = 8'd38; b_mant1 = 8'd141; b_mant2 = 8'd237; b_mant3 = 8'd89;
a_exp0 = 10'd995; a_exp1 = 10'd645; a_exp2 = 10'd572; a_exp3 = 10'd55;
b_exp0 = 10'd661; b_exp1 = 10'd297; b_exp2 = 10'd375; b_exp3 = 10'd126;
a_sign0 = 4'd1; a_sign1 = 4'd1; a_sign2 = 4'd16; a_sign3 = 4'd0;
b_sign0 = 4'd1; b_sign1 = 4'd14; b_sign2 = 4'd16; b_sign3 = 4'd9;
@(posedge clk_i);
a_mant0 = 8'd35; a_mant1 = 8'd124; a_mant2 = 8'd200; a_mant3 = 8'd135;
b_mant0 = 8'd170; b_mant1 = 8'd41; b_mant2 = 8'd168; b_mant3 = 8'd39;
a_exp0 = 10'd395; a_exp1 = 10'd224; a_exp2 = 10'd425; a_exp3 = 10'd240;
b_exp0 = 10'd732; b_exp1 = 10'd643; b_exp2 = 10'd714; b_exp3 = 10'd691;
a_sign0 = 4'd11; a_sign1 = 4'd6; a_sign2 = 4'd8; a_sign3 = 4'd0;
b_sign0 = 4'd6; b_sign1 = 4'd4; b_sign2 = 4'd13; b_sign3 = 4'd11;
@(posedge clk_i);
a_mant0 = 8'd51; a_mant1 = 8'd189; a_mant2 = 8'd50; a_mant3 = 8'd101;
b_mant0 = 8'd162; b_mant1 = 8'd216; b_mant2 = 8'd172; b_mant3 = 8'd28;
a_exp0 = 10'd585; a_exp1 = 10'd478; a_exp2 = 10'd386; a_exp3 = 10'd107;
b_exp0 = 10'd777; b_exp1 = 10'd40; b_exp2 = 10'd278; b_exp3 = 10'd440;
a_sign0 = 4'd6; a_sign1 = 4'd11; a_sign2 = 4'd12; a_sign3 = 4'd14;
b_sign0 = 4'd14; b_sign1 = 4'd12; b_sign2 = 4'd3; b_sign3 = 4'd6;
@(posedge clk_i);
a_mant0 = 8'd32; a_mant1 = 8'd210; a_mant2 = 8'd40; a_mant3 = 8'd70;
b_mant0 = 8'd196; b_mant1 = 8'd168; b_mant2 = 8'd25; b_mant3 = 8'd172;
a_exp0 = 10'd594; a_exp1 = 10'd587; a_exp2 = 10'd572; a_exp3 = 10'd25;
b_exp0 = 10'd152; b_exp1 = 10'd215; b_exp2 = 10'd81; b_exp3 = 10'd859;
a_sign0 = 4'd13; a_sign1 = 4'd2; a_sign2 = 4'd12; a_sign3 = 4'd11;
b_sign0 = 4'd16; b_sign1 = 4'd14; b_sign2 = 4'd11; b_sign3 = 4'd5;
@(posedge clk_i);
a_mant0 = 8'd247; a_mant1 = 8'd60; a_mant2 = 8'd181; a_mant3 = 8'd29;
b_mant0 = 8'd76; b_mant1 = 8'd213; b_mant2 = 8'd170; b_mant3 = 8'd171;
a_exp0 = 10'd1003; a_exp1 = 10'd642; a_exp2 = 10'd887; a_exp3 = 10'd802;
b_exp0 = 10'd289; b_exp1 = 10'd527; b_exp2 = 10'd847; b_exp3 = 10'd927;
a_sign0 = 4'd9; a_sign1 = 4'd2; a_sign2 = 4'd0; a_sign3 = 4'd6;
b_sign0 = 4'd1; b_sign1 = 4'd0; b_sign2 = 4'd2; b_sign3 = 4'd14;
@(posedge clk_i);
a_mant0 = 8'd222; a_mant1 = 8'd40; a_mant2 = 8'd71; a_mant3 = 8'd211;
b_mant0 = 8'd188; b_mant1 = 8'd224; b_mant2 = 8'd193; b_mant3 = 8'd160;
a_exp0 = 10'd848; a_exp1 = 10'd651; a_exp2 = 10'd42; a_exp3 = 10'd877;
b_exp0 = 10'd765; b_exp1 = 10'd250; b_exp2 = 10'd239; b_exp3 = 10'd998;
a_sign0 = 4'd10; a_sign1 = 4'd13; a_sign2 = 4'd5; a_sign3 = 4'd14;
b_sign0 = 4'd3; b_sign1 = 4'd13; b_sign2 = 4'd9; b_sign3 = 4'd6;
@(posedge clk_i);
shared_exps0 = 8'd150;
shared_exps1 = 8'd141;
a_mant0 = 8'd239; a_mant1 = 8'd241; a_mant2 = 8'd6; a_mant3 = 8'd41;
b_mant0 = 8'd96; b_mant1 = 8'd221; b_mant2 = 8'd127; b_mant3 = 8'd182;
a_exp0 = 10'd768; a_exp1 = 10'd33; a_exp2 = 10'd340; a_exp3 = 10'd23;
b_exp0 = 10'd637; b_exp1 = 10'd436; b_exp2 = 10'd829; b_exp3 = 10'd194;
a_sign0 = 4'd0; a_sign1 = 4'd0; a_sign2 = 4'd7; a_sign3 = 4'd14;
b_sign0 = 4'd13; b_sign1 = 4'd2; b_sign2 = 4'd9; b_sign3 = 4'd15;
@(posedge clk_i);
a_mant0 = 8'd192; a_mant1 = 8'd127; a_mant2 = 8'd161; a_mant3 = 8'd86;
b_mant0 = 8'd238; b_mant1 = 8'd117; b_mant2 = 8'd133; b_mant3 = 8'd163;
a_exp0 = 10'd812; a_exp1 = 10'd900; a_exp2 = 10'd509; a_exp3 = 10'd596;
b_exp0 = 10'd1009; b_exp1 = 10'd524; b_exp2 = 10'd579; b_exp3 = 10'd175;
a_sign0 = 4'd9; a_sign1 = 4'd13; a_sign2 = 4'd3; a_sign3 = 4'd10;
b_sign0 = 4'd6; b_sign1 = 4'd4; b_sign2 = 4'd2; b_sign3 = 4'd12;
@(posedge clk_i);
a_mant0 = 8'd1; a_mant1 = 8'd140; a_mant2 = 8'd3; a_mant3 = 8'd85;
b_mant0 = 8'd163; b_mant1 = 8'd33; b_mant2 = 8'd170; b_mant3 = 8'd8;
a_exp0 = 10'd364; a_exp1 = 10'd1019; a_exp2 = 10'd242; a_exp3 = 10'd860;
b_exp0 = 10'd291; b_exp1 = 10'd612; b_exp2 = 10'd902; b_exp3 = 10'd871;
a_sign0 = 4'd13; a_sign1 = 4'd6; a_sign2 = 4'd1; a_sign3 = 4'd9;
b_sign0 = 4'd14; b_sign1 = 4'd2; b_sign2 = 4'd12; b_sign3 = 4'd14;
@(posedge clk_i);
a_mant0 = 8'd131; a_mant1 = 8'd191; a_mant2 = 8'd196; a_mant3 = 8'd222;
b_mant0 = 8'd223; b_mant1 = 8'd67; b_mant2 = 8'd135; b_mant3 = 8'd104;
a_exp0 = 10'd334; a_exp1 = 10'd841; a_exp2 = 10'd908; a_exp3 = 10'd577;
b_exp0 = 10'd912; b_exp1 = 10'd882; b_exp2 = 10'd995; b_exp3 = 10'd180;
a_sign0 = 4'd0; a_sign1 = 4'd12; a_sign2 = 4'd7; a_sign3 = 4'd11;
b_sign0 = 4'd3; b_sign1 = 4'd13; b_sign2 = 4'd15; b_sign3 = 4'd3;
@(posedge clk_i);
a_mant0 = 8'd237; a_mant1 = 8'd76; a_mant2 = 8'd43; a_mant3 = 8'd175;
b_mant0 = 8'd204; b_mant1 = 8'd194; b_mant2 = 8'd143; b_mant3 = 8'd16;
a_exp0 = 10'd476; a_exp1 = 10'd493; a_exp2 = 10'd349; a_exp3 = 10'd360;
b_exp0 = 10'd70; b_exp1 = 10'd73; b_exp2 = 10'd126; b_exp3 = 10'd321;
a_sign0 = 4'd14; a_sign1 = 4'd14; a_sign2 = 4'd4; a_sign3 = 4'd8;
b_sign0 = 4'd14; b_sign1 = 4'd7; b_sign2 = 4'd1; b_sign3 = 4'd11;
@(posedge clk_i);
a_mant0 = 8'd250; a_mant1 = 8'd67; a_mant2 = 8'd115; a_mant3 = 8'd255;
b_mant0 = 8'd216; b_mant1 = 8'd190; b_mant2 = 8'd192; b_mant3 = 8'd136;
a_exp0 = 10'd303; a_exp1 = 10'd963; a_exp2 = 10'd803; a_exp3 = 10'd730;
b_exp0 = 10'd673; b_exp1 = 10'd570; b_exp2 = 10'd668; b_exp3 = 10'd693;
a_sign0 = 4'd6; a_sign1 = 4'd13; a_sign2 = 4'd8; a_sign3 = 4'd2;
b_sign0 = 4'd5; b_sign1 = 4'd9; b_sign2 = 4'd12; b_sign3 = 4'd7;
@(posedge clk_i);
a_mant0 = 8'd109; a_mant1 = 8'd207; a_mant2 = 8'd217; a_mant3 = 8'd102;
b_mant0 = 8'd125; b_mant1 = 8'd217; b_mant2 = 8'd22; b_mant3 = 8'd47;
a_exp0 = 10'd161; a_exp1 = 10'd186; a_exp2 = 10'd220; a_exp3 = 10'd392;
b_exp0 = 10'd382; b_exp1 = 10'd1018; b_exp2 = 10'd963; b_exp3 = 10'd96;
a_sign0 = 4'd5; a_sign1 = 4'd5; a_sign2 = 4'd12; a_sign3 = 4'd9;
b_sign0 = 4'd11; b_sign1 = 4'd13; b_sign2 = 4'd6; b_sign3 = 4'd3;
@(posedge clk_i);
a_mant0 = 8'd60; a_mant1 = 8'd29; a_mant2 = 8'd227; a_mant3 = 8'd162;
b_mant0 = 8'd168; b_mant1 = 8'd122; b_mant2 = 8'd111; b_mant3 = 8'd83;
a_exp0 = 10'd213; a_exp1 = 10'd128; a_exp2 = 10'd60; a_exp3 = 10'd488;
b_exp0 = 10'd713; b_exp1 = 10'd61; b_exp2 = 10'd872; b_exp3 = 10'd488;
a_sign0 = 4'd3; a_sign1 = 4'd16; a_sign2 = 4'd3; a_sign3 = 4'd1;
b_sign0 = 4'd2; b_sign1 = 4'd12; b_sign2 = 4'd15; b_sign3 = 4'd4;
@(posedge clk_i);
shared_exps0 = 8'd118;
shared_exps1 = 8'd144;
a_mant0 = 8'd209; a_mant1 = 8'd157; a_mant2 = 8'd79; a_mant3 = 8'd128;
b_mant0 = 8'd68; b_mant1 = 8'd125; b_mant2 = 8'd36; b_mant3 = 8'd235;
a_exp0 = 10'd71; a_exp1 = 10'd442; a_exp2 = 10'd803; a_exp3 = 10'd533;
b_exp0 = 10'd917; b_exp1 = 10'd501; b_exp2 = 10'd850; b_exp3 = 10'd486;
a_sign0 = 4'd4; a_sign1 = 4'd3; a_sign2 = 4'd6; a_sign3 = 4'd7;
b_sign0 = 4'd14; b_sign1 = 4'd11; b_sign2 = 4'd6; b_sign3 = 4'd12;
@(posedge clk_i);
a_mant0 = 8'd17; a_mant1 = 8'd220; a_mant2 = 8'd172; a_mant3 = 8'd25;
b_mant0 = 8'd57; b_mant1 = 8'd85; b_mant2 = 8'd131; b_mant3 = 8'd167;
a_exp0 = 10'd766; a_exp1 = 10'd112; a_exp2 = 10'd603; a_exp3 = 10'd930;
b_exp0 = 10'd913; b_exp1 = 10'd706; b_exp2 = 10'd165; b_exp3 = 10'd880;
a_sign0 = 4'd12; a_sign1 = 4'd2; a_sign2 = 4'd7; a_sign3 = 4'd5;
b_sign0 = 4'd0; b_sign1 = 4'd6; b_sign2 = 4'd16; b_sign3 = 4'd1;
@(posedge clk_i);
a_mant0 = 8'd79; a_mant1 = 8'd54; a_mant2 = 8'd208; a_mant3 = 8'd231;
b_mant0 = 8'd218; b_mant1 = 8'd103; b_mant2 = 8'd178; b_mant3 = 8'd58;
a_exp0 = 10'd409; a_exp1 = 10'd530; a_exp2 = 10'd224; a_exp3 = 10'd573;
b_exp0 = 10'd645; b_exp1 = 10'd1019; b_exp2 = 10'd541; b_exp3 = 10'd225;
a_sign0 = 4'd16; a_sign1 = 4'd11; a_sign2 = 4'd10; a_sign3 = 4'd5;
b_sign0 = 4'd9; b_sign1 = 4'd10; b_sign2 = 4'd14; b_sign3 = 4'd7;
@(posedge clk_i);
a_mant0 = 8'd35; a_mant1 = 8'd208; a_mant2 = 8'd171; a_mant3 = 8'd183;
b_mant0 = 8'd140; b_mant1 = 8'd8; b_mant2 = 8'd35; b_mant3 = 8'd67;
a_exp0 = 10'd225; a_exp1 = 10'd938; a_exp2 = 10'd201; a_exp3 = 10'd275;
b_exp0 = 10'd418; b_exp1 = 10'd289; b_exp2 = 10'd653; b_exp3 = 10'd412;
a_sign0 = 4'd3; a_sign1 = 4'd9; a_sign2 = 4'd16; a_sign3 = 4'd8;
b_sign0 = 4'd6; b_sign1 = 4'd15; b_sign2 = 4'd14; b_sign3 = 4'd7;
@(posedge clk_i);
a_mant0 = 8'd215; a_mant1 = 8'd185; a_mant2 = 8'd70; a_mant3 = 8'd88;
b_mant0 = 8'd132; b_mant1 = 8'd237; b_mant2 = 8'd219; b_mant3 = 8'd47;
a_exp0 = 10'd287; a_exp1 = 10'd640; a_exp2 = 10'd822; a_exp3 = 10'd862;
b_exp0 = 10'd21; b_exp1 = 10'd643; b_exp2 = 10'd139; b_exp3 = 10'd127;
a_sign0 = 4'd10; a_sign1 = 4'd12; a_sign2 = 4'd11; a_sign3 = 4'd14;
b_sign0 = 4'd16; b_sign1 = 4'd11; b_sign2 = 4'd4; b_sign3 = 4'd4;
@(posedge clk_i);
a_mant0 = 8'd162; a_mant1 = 8'd133; a_mant2 = 8'd59; a_mant3 = 8'd65;
b_mant0 = 8'd48; b_mant1 = 8'd124; b_mant2 = 8'd242; b_mant3 = 8'd200;
a_exp0 = 10'd528; a_exp1 = 10'd391; a_exp2 = 10'd402; a_exp3 = 10'd13;
b_exp0 = 10'd840; b_exp1 = 10'd652; b_exp2 = 10'd210; b_exp3 = 10'd893;
a_sign0 = 4'd12; a_sign1 = 4'd12; a_sign2 = 4'd12; a_sign3 = 4'd12;
b_sign0 = 4'd6; b_sign1 = 4'd2; b_sign2 = 4'd2; b_sign3 = 4'd13;
@(posedge clk_i);
a_mant0 = 8'd45; a_mant1 = 8'd68; a_mant2 = 8'd145; a_mant3 = 8'd113;
b_mant0 = 8'd244; b_mant1 = 8'd145; b_mant2 = 8'd28; b_mant3 = 8'd86;
a_exp0 = 10'd646; a_exp1 = 10'd676; a_exp2 = 10'd494; a_exp3 = 10'd559;
b_exp0 = 10'd478; b_exp1 = 10'd456; b_exp2 = 10'd773; b_exp3 = 10'd287;
a_sign0 = 4'd5; a_sign1 = 4'd2; a_sign2 = 4'd15; a_sign3 = 4'd7;
b_sign0 = 4'd10; b_sign1 = 4'd14; b_sign2 = 4'd16; b_sign3 = 4'd13;
@(posedge clk_i);
a_mant0 = 8'd135; a_mant1 = 8'd83; a_mant2 = 8'd88; a_mant3 = 8'd156;
b_mant0 = 8'd8; b_mant1 = 8'd145; b_mant2 = 8'd238; b_mant3 = 8'd56;
a_exp0 = 10'd947; a_exp1 = 10'd443; a_exp2 = 10'd148; a_exp3 = 10'd353;
b_exp0 = 10'd455; b_exp1 = 10'd720; b_exp2 = 10'd655; b_exp3 = 10'd638;
a_sign0 = 4'd11; a_sign1 = 4'd13; a_sign2 = 4'd11; a_sign3 = 4'd9;
b_sign0 = 4'd0; b_sign1 = 4'd16; b_sign2 = 4'd5; b_sign3 = 4'd1;
@(posedge clk_i);
shared_exps0 = 8'd122;
shared_exps1 = 8'd119;
rstn = 0;
@(posedge clk_i);
rstn = 1;
a_mant0 = 8'd39; a_mant1 = 8'd171; a_mant2 = 8'd98; a_mant3 = 8'd210;
b_mant0 = 8'd209; b_mant1 = 8'd40; b_mant2 = 8'd182; b_mant3 = 8'd132;
a_exp0 = 10'd977; a_exp1 = 10'd689; a_exp2 = 10'd654; a_exp3 = 10'd38;
b_exp0 = 10'd53; b_exp1 = 10'd809; b_exp2 = 10'd193; b_exp3 = 10'd551;
a_sign0 = 4'd0; a_sign1 = 4'd1; a_sign2 = 4'd14; a_sign3 = 4'd8;
b_sign0 = 4'd14; b_sign1 = 4'd10; b_sign2 = 4'd3; b_sign3 = 4'd6;
@(posedge clk_i);
a_mant0 = 8'd249; a_mant1 = 8'd28; a_mant2 = 8'd157; a_mant3 = 8'd86;
b_mant0 = 8'd30; b_mant1 = 8'd178; b_mant2 = 8'd155; b_mant3 = 8'd120;
a_exp0 = 10'd229; a_exp1 = 10'd212; a_exp2 = 10'd512; a_exp3 = 10'd875;
b_exp0 = 10'd930; b_exp1 = 10'd228; b_exp2 = 10'd207; b_exp3 = 10'd1007;
a_sign0 = 4'd8; a_sign1 = 4'd8; a_sign2 = 4'd9; a_sign3 = 4'd8;
b_sign0 = 4'd0; b_sign1 = 4'd5; b_sign2 = 4'd2; b_sign3 = 4'd6;
@(posedge clk_i);
a_mant0 = 8'd107; a_mant1 = 8'd28; a_mant2 = 8'd63; a_mant3 = 8'd4;
b_mant0 = 8'd233; b_mant1 = 8'd52; b_mant2 = 8'd80; b_mant3 = 8'd4;
a_exp0 = 10'd99; a_exp1 = 10'd642; a_exp2 = 10'd952; a_exp3 = 10'd407;
b_exp0 = 10'd670; b_exp1 = 10'd419; b_exp2 = 10'd510; b_exp3 = 10'd384;
a_sign0 = 4'd12; a_sign1 = 4'd3; a_sign2 = 4'd8; a_sign3 = 4'd1;
b_sign0 = 4'd1; b_sign1 = 4'd3; b_sign2 = 4'd16; b_sign3 = 4'd11;
@(posedge clk_i);
a_mant0 = 8'd38; a_mant1 = 8'd102; a_mant2 = 8'd233; a_mant3 = 8'd139;
b_mant0 = 8'd177; b_mant1 = 8'd70; b_mant2 = 8'd178; b_mant3 = 8'd215;
a_exp0 = 10'd723; a_exp1 = 10'd505; a_exp2 = 10'd569; a_exp3 = 10'd594;
b_exp0 = 10'd60; b_exp1 = 10'd295; b_exp2 = 10'd68; b_exp3 = 10'd47;
a_sign0 = 4'd16; a_sign1 = 4'd12; a_sign2 = 4'd2; a_sign3 = 4'd13;
b_sign0 = 4'd13; b_sign1 = 4'd13; b_sign2 = 4'd1; b_sign3 = 4'd0;
@(posedge clk_i);
a_mant0 = 8'd44; a_mant1 = 8'd62; a_mant2 = 8'd139; a_mant3 = 8'd183;
b_mant0 = 8'd2; b_mant1 = 8'd246; b_mant2 = 8'd58; b_mant3 = 8'd123;
a_exp0 = 10'd818; a_exp1 = 10'd153; a_exp2 = 10'd478; a_exp3 = 10'd742;
b_exp0 = 10'd154; b_exp1 = 10'd263; b_exp2 = 10'd983; b_exp3 = 10'd640;
a_sign0 = 4'd14; a_sign1 = 4'd13; a_sign2 = 4'd11; a_sign3 = 4'd0;
b_sign0 = 4'd13; b_sign1 = 4'd6; b_sign2 = 4'd7; b_sign3 = 4'd6;
@(posedge clk_i);
a_mant0 = 8'd214; a_mant1 = 8'd60; a_mant2 = 8'd80; a_mant3 = 8'd31;
b_mant0 = 8'd156; b_mant1 = 8'd105; b_mant2 = 8'd130; b_mant3 = 8'd77;
a_exp0 = 10'd314; a_exp1 = 10'd899; a_exp2 = 10'd52; a_exp3 = 10'd285;
b_exp0 = 10'd975; b_exp1 = 10'd683; b_exp2 = 10'd895; b_exp3 = 10'd753;
a_sign0 = 4'd11; a_sign1 = 4'd15; a_sign2 = 4'd15; a_sign3 = 4'd9;
b_sign0 = 4'd16; b_sign1 = 4'd11; b_sign2 = 4'd16; b_sign3 = 4'd0;
@(posedge clk_i);
a_mant0 = 8'd198; a_mant1 = 8'd233; a_mant2 = 8'd222; a_mant3 = 8'd150;
b_mant0 = 8'd240; b_mant1 = 8'd144; b_mant2 = 8'd28; b_mant3 = 8'd176;
a_exp0 = 10'd705; a_exp1 = 10'd257; a_exp2 = 10'd89; a_exp3 = 10'd321;
b_exp0 = 10'd744; b_exp1 = 10'd290; b_exp2 = 10'd503; b_exp3 = 10'd561;
a_sign0 = 4'd7; a_sign1 = 4'd8; a_sign2 = 4'd1; a_sign3 = 4'd16;
b_sign0 = 4'd10; b_sign1 = 4'd4; b_sign2 = 4'd1; b_sign3 = 4'd15;
@(posedge clk_i);
shared_exps0 = 8'd136;
shared_exps1 = 8'd119;
a_mant0 = 8'd172; a_mant1 = 8'd66; a_mant2 = 8'd200; a_mant3 = 8'd178;
b_mant0 = 8'd200; b_mant1 = 8'd203; b_mant2 = 8'd252; b_mant3 = 8'd108;
a_exp0 = 10'd477; a_exp1 = 10'd174; a_exp2 = 10'd109; a_exp3 = 10'd754;
b_exp0 = 10'd352; b_exp1 = 10'd320; b_exp2 = 10'd499; b_exp3 = 10'd913;
a_sign0 = 4'd5; a_sign1 = 4'd7; a_sign2 = 4'd10; a_sign3 = 4'd1;
b_sign0 = 4'd7; b_sign1 = 4'd8; b_sign2 = 4'd10; b_sign3 = 4'd2;
@(posedge clk_i);
a_mant0 = 8'd119; a_mant1 = 8'd144; a_mant2 = 8'd10; a_mant3 = 8'd242;
b_mant0 = 8'd246; b_mant1 = 8'd88; b_mant2 = 8'd229; b_mant3 = 8'd97;
a_exp0 = 10'd247; a_exp1 = 10'd365; a_exp2 = 10'd211; a_exp3 = 10'd719;
b_exp0 = 10'd382; b_exp1 = 10'd607; b_exp2 = 10'd504; b_exp3 = 10'd506;
a_sign0 = 4'd8; a_sign1 = 4'd6; a_sign2 = 4'd15; a_sign3 = 4'd7;
b_sign0 = 4'd7; b_sign1 = 4'd11; b_sign2 = 4'd5; b_sign3 = 4'd2;
@(posedge clk_i);
a_mant0 = 8'd162; a_mant1 = 8'd200; a_mant2 = 8'd73; a_mant3 = 8'd131;
b_mant0 = 8'd36; b_mant1 = 8'd4; b_mant2 = 8'd213; b_mant3 = 8'd220;
a_exp0 = 10'd865; a_exp1 = 10'd986; a_exp2 = 10'd528; a_exp3 = 10'd86;
b_exp0 = 10'd481; b_exp1 = 10'd86; b_exp2 = 10'd261; b_exp3 = 10'd170;
a_sign0 = 4'd14; a_sign1 = 4'd7; a_sign2 = 4'd3; a_sign3 = 4'd6;
b_sign0 = 4'd12; b_sign1 = 4'd5; b_sign2 = 4'd4; b_sign3 = 4'd10;
@(posedge clk_i);
a_mant0 = 8'd199; a_mant1 = 8'd68; a_mant2 = 8'd34; a_mant3 = 8'd86;
b_mant0 = 8'd61; b_mant1 = 8'd146; b_mant2 = 8'd96; b_mant3 = 8'd82;
a_exp0 = 10'd705; a_exp1 = 10'd992; a_exp2 = 10'd658; a_exp3 = 10'd724;
b_exp0 = 10'd778; b_exp1 = 10'd341; b_exp2 = 10'd900; b_exp3 = 10'd939;
a_sign0 = 4'd4; a_sign1 = 4'd2; a_sign2 = 4'd16; a_sign3 = 4'd11;
b_sign0 = 4'd2; b_sign1 = 4'd15; b_sign2 = 4'd15; b_sign3 = 4'd6;
@(posedge clk_i);
a_mant0 = 8'd181; a_mant1 = 8'd198; a_mant2 = 8'd234; a_mant3 = 8'd190;
b_mant0 = 8'd73; b_mant1 = 8'd42; b_mant2 = 8'd154; b_mant3 = 8'd225;
a_exp0 = 10'd1002; a_exp1 = 10'd916; a_exp2 = 10'd60; a_exp3 = 10'd645;
b_exp0 = 10'd200; b_exp1 = 10'd765; b_exp2 = 10'd254; b_exp3 = 10'd760;
a_sign0 = 4'd0; a_sign1 = 4'd1; a_sign2 = 4'd16; a_sign3 = 4'd2;
b_sign0 = 4'd4; b_sign1 = 4'd4; b_sign2 = 4'd9; b_sign3 = 4'd0;
@(posedge clk_i);
a_mant0 = 8'd250; a_mant1 = 8'd71; a_mant2 = 8'd178; a_mant3 = 8'd67;
b_mant0 = 8'd27; b_mant1 = 8'd81; b_mant2 = 8'd233; b_mant3 = 8'd100;
a_exp0 = 10'd815; a_exp1 = 10'd574; a_exp2 = 10'd111; a_exp3 = 10'd969;
b_exp0 = 10'd732; b_exp1 = 10'd59; b_exp2 = 10'd643; b_exp3 = 10'd893;
a_sign0 = 4'd11; a_sign1 = 4'd4; a_sign2 = 4'd4; a_sign3 = 4'd5;
b_sign0 = 4'd1; b_sign1 = 4'd2; b_sign2 = 4'd1; b_sign3 = 4'd8;
@(posedge clk_i);
a_mant0 = 8'd116; a_mant1 = 8'd112; a_mant2 = 8'd80; a_mant3 = 8'd76;
b_mant0 = 8'd103; b_mant1 = 8'd167; b_mant2 = 8'd23; b_mant3 = 8'd168;
a_exp0 = 10'd685; a_exp1 = 10'd652; a_exp2 = 10'd60; a_exp3 = 10'd1016;
b_exp0 = 10'd64; b_exp1 = 10'd817; b_exp2 = 10'd70; b_exp3 = 10'd562;
a_sign0 = 4'd5; a_sign1 = 4'd11; a_sign2 = 4'd11; a_sign3 = 4'd14;
b_sign0 = 4'd4; b_sign1 = 4'd4; b_sign2 = 4'd4; b_sign3 = 4'd16;
@(posedge clk_i);
a_mant0 = 8'd191; a_mant1 = 8'd246; a_mant2 = 8'd46; a_mant3 = 8'd179;
b_mant0 = 8'd77; b_mant1 = 8'd175; b_mant2 = 8'd218; b_mant3 = 8'd40;
a_exp0 = 10'd949; a_exp1 = 10'd305; a_exp2 = 10'd979; a_exp3 = 10'd59;
b_exp0 = 10'd587; b_exp1 = 10'd898; b_exp2 = 10'd1006; b_exp3 = 10'd1013;
a_sign0 = 4'd10; a_sign1 = 4'd11; a_sign2 = 4'd3; a_sign3 = 4'd9;
b_sign0 = 4'd2; b_sign1 = 4'd3; b_sign2 = 4'd5; b_sign3 = 4'd1;
@(posedge clk_i);
shared_exps0 = 8'd118;
shared_exps1 = 8'd140;
a_mant0 = 8'd182; a_mant1 = 8'd116; a_mant2 = 8'd2; a_mant3 = 8'd101;
b_mant0 = 8'd114; b_mant1 = 8'd39; b_mant2 = 8'd107; b_mant3 = 8'd151;
a_exp0 = 10'd647; a_exp1 = 10'd60; a_exp2 = 10'd854; a_exp3 = 10'd792;
b_exp0 = 10'd873; b_exp1 = 10'd315; b_exp2 = 10'd426; b_exp3 = 10'd229;
a_sign0 = 4'd12; a_sign1 = 4'd2; a_sign2 = 4'd12; a_sign3 = 4'd7;
b_sign0 = 4'd1; b_sign1 = 4'd11; b_sign2 = 4'd7; b_sign3 = 4'd14;
@(posedge clk_i);
a_mant0 = 8'd13; a_mant1 = 8'd247; a_mant2 = 8'd178; a_mant3 = 8'd1;
b_mant0 = 8'd208; b_mant1 = 8'd243; b_mant2 = 8'd249; b_mant3 = 8'd79;
a_exp0 = 10'd582; a_exp1 = 10'd661; a_exp2 = 10'd658; a_exp3 = 10'd444;
b_exp0 = 10'd343; b_exp1 = 10'd986; b_exp2 = 10'd436; b_exp3 = 10'd788;
a_sign0 = 4'd4; a_sign1 = 4'd10; a_sign2 = 4'd15; a_sign3 = 4'd9;
b_sign0 = 4'd7; b_sign1 = 4'd4; b_sign2 = 4'd14; b_sign3 = 4'd7;
@(posedge clk_i);
a_mant0 = 8'd84; a_mant1 = 8'd34; a_mant2 = 8'd116; a_mant3 = 8'd86;
b_mant0 = 8'd204; b_mant1 = 8'd140; b_mant2 = 8'd45; b_mant3 = 8'd103;
a_exp0 = 10'd542; a_exp1 = 10'd715; a_exp2 = 10'd623; a_exp3 = 10'd634;
b_exp0 = 10'd730; b_exp1 = 10'd613; b_exp2 = 10'd197; b_exp3 = 10'd80;
a_sign0 = 4'd0; a_sign1 = 4'd4; a_sign2 = 4'd4; a_sign3 = 4'd3;
b_sign0 = 4'd15; b_sign1 = 4'd14; b_sign2 = 4'd13; b_sign3 = 4'd7;
@(posedge clk_i);
a_mant0 = 8'd212; a_mant1 = 8'd236; a_mant2 = 8'd113; a_mant3 = 8'd131;
b_mant0 = 8'd222; b_mant1 = 8'd41; b_mant2 = 8'd212; b_mant3 = 8'd241;
a_exp0 = 10'd638; a_exp1 = 10'd277; a_exp2 = 10'd685; a_exp3 = 10'd762;
b_exp0 = 10'd106; b_exp1 = 10'd432; b_exp2 = 10'd693; b_exp3 = 10'd723;
a_sign0 = 4'd10; a_sign1 = 4'd0; a_sign2 = 4'd14; a_sign3 = 4'd12;
b_sign0 = 4'd16; b_sign1 = 4'd8; b_sign2 = 4'd4; b_sign3 = 4'd3;
@(posedge clk_i);
a_mant0 = 8'd124; a_mant1 = 8'd46; a_mant2 = 8'd8; a_mant3 = 8'd3;
b_mant0 = 8'd79; b_mant1 = 8'd148; b_mant2 = 8'd149; b_mant3 = 8'd180;
a_exp0 = 10'd335; a_exp1 = 10'd59; a_exp2 = 10'd260; a_exp3 = 10'd77;
b_exp0 = 10'd401; b_exp1 = 10'd186; b_exp2 = 10'd862; b_exp3 = 10'd911;
a_sign0 = 4'd1; a_sign1 = 4'd2; a_sign2 = 4'd2; a_sign3 = 4'd13;
b_sign0 = 4'd15; b_sign1 = 4'd1; b_sign2 = 4'd8; b_sign3 = 4'd10;
@(posedge clk_i);
a_mant0 = 8'd248; a_mant1 = 8'd36; a_mant2 = 8'd132; a_mant3 = 8'd136;
b_mant0 = 8'd117; b_mant1 = 8'd69; b_mant2 = 8'd179; b_mant3 = 8'd211;
a_exp0 = 10'd969; a_exp1 = 10'd325; a_exp2 = 10'd544; a_exp3 = 10'd758;
b_exp0 = 10'd213; b_exp1 = 10'd426; b_exp2 = 10'd247; b_exp3 = 10'd924;
a_sign0 = 4'd5; a_sign1 = 4'd5; a_sign2 = 4'd14; a_sign3 = 4'd3;
b_sign0 = 4'd4; b_sign1 = 4'd3; b_sign2 = 4'd0; b_sign3 = 4'd6;
@(posedge clk_i);
a_mant0 = 8'd26; a_mant1 = 8'd207; a_mant2 = 8'd173; a_mant3 = 8'd33;
b_mant0 = 8'd118; b_mant1 = 8'd69; b_mant2 = 8'd70; b_mant3 = 8'd228;
a_exp0 = 10'd584; a_exp1 = 10'd376; a_exp2 = 10'd341; a_exp3 = 10'd729;
b_exp0 = 10'd288; b_exp1 = 10'd489; b_exp2 = 10'd738; b_exp3 = 10'd712;
a_sign0 = 4'd13; a_sign1 = 4'd2; a_sign2 = 4'd15; a_sign3 = 4'd7;
b_sign0 = 4'd3; b_sign1 = 4'd1; b_sign2 = 4'd8; b_sign3 = 4'd15;
@(posedge clk_i);
a_mant0 = 8'd214; a_mant1 = 8'd158; a_mant2 = 8'd57; a_mant3 = 8'd107;
b_mant0 = 8'd183; b_mant1 = 8'd44; b_mant2 = 8'd148; b_mant3 = 8'd36;
a_exp0 = 10'd154; a_exp1 = 10'd255; a_exp2 = 10'd176; a_exp3 = 10'd536;
b_exp0 = 10'd180; b_exp1 = 10'd163; b_exp2 = 10'd870; b_exp3 = 10'd616;
a_sign0 = 4'd13; a_sign1 = 4'd2; a_sign2 = 4'd1; a_sign3 = 4'd11;
b_sign0 = 4'd5; b_sign1 = 4'd7; b_sign2 = 4'd15; b_sign3 = 4'd10;
@(posedge clk_i);
shared_exps0 = 8'd136;
shared_exps1 = 8'd126;
a_mant0 = 8'd85; a_mant1 = 8'd231; a_mant2 = 8'd131; a_mant3 = 8'd7;
b_mant0 = 8'd53; b_mant1 = 8'd131; b_mant2 = 8'd193; b_mant3 = 8'd25;
a_exp0 = 10'd292; a_exp1 = 10'd341; a_exp2 = 10'd747; a_exp3 = 10'd478;
b_exp0 = 10'd25; b_exp1 = 10'd142; b_exp2 = 10'd977; b_exp3 = 10'd395;
a_sign0 = 4'd3; a_sign1 = 4'd13; a_sign2 = 4'd8; a_sign3 = 4'd8;
b_sign0 = 4'd3; b_sign1 = 4'd12; b_sign2 = 4'd15; b_sign3 = 4'd8;
@(posedge clk_i);
a_mant0 = 8'd216; a_mant1 = 8'd8; a_mant2 = 8'd32; a_mant3 = 8'd175;
b_mant0 = 8'd3; b_mant1 = 8'd134; b_mant2 = 8'd32; b_mant3 = 8'd110;
a_exp0 = 10'd582; a_exp1 = 10'd515; a_exp2 = 10'd624; a_exp3 = 10'd141;
b_exp0 = 10'd1000; b_exp1 = 10'd371; b_exp2 = 10'd764; b_exp3 = 10'd525;
a_sign0 = 4'd12; a_sign1 = 4'd7; a_sign2 = 4'd6; a_sign3 = 4'd9;
b_sign0 = 4'd10; b_sign1 = 4'd4; b_sign2 = 4'd15; b_sign3 = 4'd10;
@(posedge clk_i);
a_mant0 = 8'd163; a_mant1 = 8'd12; a_mant2 = 8'd139; a_mant3 = 8'd48;
b_mant0 = 8'd93; b_mant1 = 8'd117; b_mant2 = 8'd227; b_mant3 = 8'd84;
a_exp0 = 10'd341; a_exp1 = 10'd428; a_exp2 = 10'd514; a_exp3 = 10'd699;
b_exp0 = 10'd257; b_exp1 = 10'd491; b_exp2 = 10'd843; b_exp3 = 10'd1005;
a_sign0 = 4'd6; a_sign1 = 4'd14; a_sign2 = 4'd13; a_sign3 = 4'd14;
b_sign0 = 4'd2; b_sign1 = 4'd6; b_sign2 = 4'd7; b_sign3 = 4'd1;
@(posedge clk_i);
a_mant0 = 8'd80; a_mant1 = 8'd224; a_mant2 = 8'd106; a_mant3 = 8'd196;
b_mant0 = 8'd43; b_mant1 = 8'd73; b_mant2 = 8'd76; b_mant3 = 8'd85;
a_exp0 = 10'd90; a_exp1 = 10'd383; a_exp2 = 10'd444; a_exp3 = 10'd1009;
b_exp0 = 10'd922; b_exp1 = 10'd450; b_exp2 = 10'd541; b_exp3 = 10'd426;
a_sign0 = 4'd7; a_sign1 = 4'd15; a_sign2 = 4'd1; a_sign3 = 4'd5;
b_sign0 = 4'd14; b_sign1 = 4'd9; b_sign2 = 4'd14; b_sign3 = 4'd2;
@(posedge clk_i);
a_mant0 = 8'd107; a_mant1 = 8'd208; a_mant2 = 8'd45; a_mant3 = 8'd50;
b_mant0 = 8'd187; b_mant1 = 8'd15; b_mant2 = 8'd10; b_mant3 = 8'd92;
a_exp0 = 10'd907; a_exp1 = 10'd580; a_exp2 = 10'd70; a_exp3 = 10'd489;
b_exp0 = 10'd81; b_exp1 = 10'd374; b_exp2 = 10'd609; b_exp3 = 10'd1019;
a_sign0 = 4'd8; a_sign1 = 4'd15; a_sign2 = 4'd10; a_sign3 = 4'd3;
b_sign0 = 4'd15; b_sign1 = 4'd11; b_sign2 = 4'd5; b_sign3 = 4'd11;
@(posedge clk_i);
a_mant0 = 8'd42; a_mant1 = 8'd56; a_mant2 = 8'd147; a_mant3 = 8'd5;
b_mant0 = 8'd124; b_mant1 = 8'd170; b_mant2 = 8'd47; b_mant3 = 8'd93;
a_exp0 = 10'd173; a_exp1 = 10'd267; a_exp2 = 10'd715; a_exp3 = 10'd761;
b_exp0 = 10'd698; b_exp1 = 10'd125; b_exp2 = 10'd64; b_exp3 = 10'd485;
a_sign0 = 4'd2; a_sign1 = 4'd3; a_sign2 = 4'd12; a_sign3 = 4'd7;
b_sign0 = 4'd13; b_sign1 = 4'd8; b_sign2 = 4'd2; b_sign3 = 4'd11;
@(posedge clk_i);
a_mant0 = 8'd199; a_mant1 = 8'd234; a_mant2 = 8'd208; a_mant3 = 8'd94;
b_mant0 = 8'd153; b_mant1 = 8'd150; b_mant2 = 8'd46; b_mant3 = 8'd52;
a_exp0 = 10'd852; a_exp1 = 10'd620; a_exp2 = 10'd157; a_exp3 = 10'd32;
b_exp0 = 10'd743; b_exp1 = 10'd665; b_exp2 = 10'd741; b_exp3 = 10'd6;
a_sign0 = 4'd11; a_sign1 = 4'd7; a_sign2 = 4'd13; a_sign3 = 4'd16;
b_sign0 = 4'd16; b_sign1 = 4'd7; b_sign2 = 4'd5; b_sign3 = 4'd11;
@(posedge clk_i);
a_mant0 = 8'd164; a_mant1 = 8'd54; a_mant2 = 8'd30; a_mant3 = 8'd179;
b_mant0 = 8'd214; b_mant1 = 8'd21; b_mant2 = 8'd146; b_mant3 = 8'd114;
a_exp0 = 10'd120; a_exp1 = 10'd640; a_exp2 = 10'd856; a_exp3 = 10'd506;
b_exp0 = 10'd362; b_exp1 = 10'd514; b_exp2 = 10'd257; b_exp3 = 10'd364;
a_sign0 = 4'd3; a_sign1 = 4'd0; a_sign2 = 4'd4; a_sign3 = 4'd2;
b_sign0 = 4'd6; b_sign1 = 4'd8; b_sign2 = 4'd5; b_sign3 = 4'd8;
@(posedge clk_i);
shared_exps0 = 8'd146;
shared_exps1 = 8'd128;
rstn = 0;
@(posedge clk_i);
rstn = 1;
a_mant0 = 8'd57; a_mant1 = 8'd56; a_mant2 = 8'd169; a_mant3 = 8'd19;
b_mant0 = 8'd93; b_mant1 = 8'd193; b_mant2 = 8'd18; b_mant3 = 8'd55;
a_exp0 = 10'd756; a_exp1 = 10'd993; a_exp2 = 10'd100; a_exp3 = 10'd190;
b_exp0 = 10'd266; b_exp1 = 10'd647; b_exp2 = 10'd647; b_exp3 = 10'd409;
a_sign0 = 4'd15; a_sign1 = 4'd0; a_sign2 = 4'd2; a_sign3 = 4'd16;
b_sign0 = 4'd8; b_sign1 = 4'd16; b_sign2 = 4'd8; b_sign3 = 4'd11;
@(posedge clk_i);
a_mant0 = 8'd157; a_mant1 = 8'd145; a_mant2 = 8'd129; a_mant3 = 8'd3;
b_mant0 = 8'd205; b_mant1 = 8'd225; b_mant2 = 8'd198; b_mant3 = 8'd1;
a_exp0 = 10'd1023; a_exp1 = 10'd986; a_exp2 = 10'd323; a_exp3 = 10'd916;
b_exp0 = 10'd740; b_exp1 = 10'd755; b_exp2 = 10'd108; b_exp3 = 10'd78;
a_sign0 = 4'd5; a_sign1 = 4'd6; a_sign2 = 4'd16; a_sign3 = 4'd12;
b_sign0 = 4'd0; b_sign1 = 4'd15; b_sign2 = 4'd7; b_sign3 = 4'd16;
@(posedge clk_i);
a_mant0 = 8'd44; a_mant1 = 8'd230; a_mant2 = 8'd178; a_mant3 = 8'd58;
b_mant0 = 8'd33; b_mant1 = 8'd38; b_mant2 = 8'd84; b_mant3 = 8'd161;
a_exp0 = 10'd983; a_exp1 = 10'd766; a_exp2 = 10'd428; a_exp3 = 10'd11;
b_exp0 = 10'd269; b_exp1 = 10'd266; b_exp2 = 10'd434; b_exp3 = 10'd538;
a_sign0 = 4'd12; a_sign1 = 4'd10; a_sign2 = 4'd0; a_sign3 = 4'd1;
b_sign0 = 4'd15; b_sign1 = 4'd16; b_sign2 = 4'd16; b_sign3 = 4'd0;
@(posedge clk_i);
a_mant0 = 8'd173; a_mant1 = 8'd238; a_mant2 = 8'd55; a_mant3 = 8'd75;
b_mant0 = 8'd97; b_mant1 = 8'd192; b_mant2 = 8'd153; b_mant3 = 8'd112;
a_exp0 = 10'd148; a_exp1 = 10'd337; a_exp2 = 10'd571; a_exp3 = 10'd904;
b_exp0 = 10'd299; b_exp1 = 10'd230; b_exp2 = 10'd117; b_exp3 = 10'd944;
a_sign0 = 4'd16; a_sign1 = 4'd10; a_sign2 = 4'd7; a_sign3 = 4'd15;
b_sign0 = 4'd1; b_sign1 = 4'd15; b_sign2 = 4'd0; b_sign3 = 4'd2;
@(posedge clk_i);
a_mant0 = 8'd253; a_mant1 = 8'd84; a_mant2 = 8'd187; a_mant3 = 8'd123;
b_mant0 = 8'd4; b_mant1 = 8'd1; b_mant2 = 8'd6; b_mant3 = 8'd79;
a_exp0 = 10'd192; a_exp1 = 10'd376; a_exp2 = 10'd304; a_exp3 = 10'd173;
b_exp0 = 10'd104; b_exp1 = 10'd324; b_exp2 = 10'd501; b_exp3 = 10'd106;
a_sign0 = 4'd3; a_sign1 = 4'd12; a_sign2 = 4'd4; a_sign3 = 4'd5;
b_sign0 = 4'd2; b_sign1 = 4'd7; b_sign2 = 4'd2; b_sign3 = 4'd15;
@(posedge clk_i);
a_mant0 = 8'd187; a_mant1 = 8'd243; a_mant2 = 8'd52; a_mant3 = 8'd118;
b_mant0 = 8'd90; b_mant1 = 8'd225; b_mant2 = 8'd26; b_mant3 = 8'd91;
a_exp0 = 10'd355; a_exp1 = 10'd218; a_exp2 = 10'd954; a_exp3 = 10'd416;
b_exp0 = 10'd738; b_exp1 = 10'd589; b_exp2 = 10'd586; b_exp3 = 10'd747;
a_sign0 = 4'd6; a_sign1 = 4'd8; a_sign2 = 4'd16; a_sign3 = 4'd1;
b_sign0 = 4'd3; b_sign1 = 4'd3; b_sign2 = 4'd13; b_sign3 = 4'd12;
@(posedge clk_i);
a_mant0 = 8'd55; a_mant1 = 8'd214; a_mant2 = 8'd253; a_mant3 = 8'd101;
b_mant0 = 8'd243; b_mant1 = 8'd66; b_mant2 = 8'd94; b_mant3 = 8'd33;
a_exp0 = 10'd912; a_exp1 = 10'd590; a_exp2 = 10'd315; a_exp3 = 10'd897;
b_exp0 = 10'd685; b_exp1 = 10'd513; b_exp2 = 10'd685; b_exp3 = 10'd862;
a_sign0 = 4'd3; a_sign1 = 4'd6; a_sign2 = 4'd7; a_sign3 = 4'd16;
b_sign0 = 4'd14; b_sign1 = 4'd3; b_sign2 = 4'd16; b_sign3 = 4'd2;
@(posedge clk_i);
shared_exps0 = 8'd122;
shared_exps1 = 8'd102;
a_mant0 = 8'd236; a_mant1 = 8'd102; a_mant2 = 8'd241; a_mant3 = 8'd234;
b_mant0 = 8'd52; b_mant1 = 8'd152; b_mant2 = 8'd249; b_mant3 = 8'd197;
a_exp0 = 10'd634; a_exp1 = 10'd60; a_exp2 = 10'd84; a_exp3 = 10'd262;
b_exp0 = 10'd342; b_exp1 = 10'd552; b_exp2 = 10'd282; b_exp3 = 10'd331;
a_sign0 = 4'd7; a_sign1 = 4'd4; a_sign2 = 4'd12; a_sign3 = 4'd0;
b_sign0 = 4'd6; b_sign1 = 4'd5; b_sign2 = 4'd0; b_sign3 = 4'd0;
@(posedge clk_i);
a_mant0 = 8'd165; a_mant1 = 8'd5; a_mant2 = 8'd102; a_mant3 = 8'd176;
b_mant0 = 8'd72; b_mant1 = 8'd202; b_mant2 = 8'd151; b_mant3 = 8'd215;
a_exp0 = 10'd414; a_exp1 = 10'd448; a_exp2 = 10'd632; a_exp3 = 10'd1015;
b_exp0 = 10'd829; b_exp1 = 10'd395; b_exp2 = 10'd631; b_exp3 = 10'd1009;
a_sign0 = 4'd2; a_sign1 = 4'd1; a_sign2 = 4'd5; a_sign3 = 4'd4;
b_sign0 = 4'd1; b_sign1 = 4'd3; b_sign2 = 4'd13; b_sign3 = 4'd10;
@(posedge clk_i);
a_mant0 = 8'd246; a_mant1 = 8'd86; a_mant2 = 8'd172; a_mant3 = 8'd250;
b_mant0 = 8'd73; b_mant1 = 8'd125; b_mant2 = 8'd214; b_mant3 = 8'd192;
a_exp0 = 10'd713; a_exp1 = 10'd250; a_exp2 = 10'd332; a_exp3 = 10'd415;
b_exp0 = 10'd409; b_exp1 = 10'd306; b_exp2 = 10'd262; b_exp3 = 10'd300;
a_sign0 = 4'd1; a_sign1 = 4'd1; a_sign2 = 4'd11; a_sign3 = 4'd3;
b_sign0 = 4'd16; b_sign1 = 4'd5; b_sign2 = 4'd3; b_sign3 = 4'd15;
@(posedge clk_i);
a_mant0 = 8'd197; a_mant1 = 8'd114; a_mant2 = 8'd77; a_mant3 = 8'd228;
b_mant0 = 8'd98; b_mant1 = 8'd5; b_mant2 = 8'd151; b_mant3 = 8'd168;
a_exp0 = 10'd79; a_exp1 = 10'd632; a_exp2 = 10'd262; a_exp3 = 10'd272;
b_exp0 = 10'd672; b_exp1 = 10'd743; b_exp2 = 10'd241; b_exp3 = 10'd128;
a_sign0 = 4'd0; a_sign1 = 4'd7; a_sign2 = 4'd5; a_sign3 = 4'd6;
b_sign0 = 4'd1; b_sign1 = 4'd16; b_sign2 = 4'd8; b_sign3 = 4'd10;
@(posedge clk_i);
a_mant0 = 8'd165; a_mant1 = 8'd70; a_mant2 = 8'd99; a_mant3 = 8'd154;
b_mant0 = 8'd36; b_mant1 = 8'd152; b_mant2 = 8'd49; b_mant3 = 8'd174;
a_exp0 = 10'd891; a_exp1 = 10'd96; a_exp2 = 10'd650; a_exp3 = 10'd199;
b_exp0 = 10'd111; b_exp1 = 10'd0; b_exp2 = 10'd207; b_exp3 = 10'd100;
a_sign0 = 4'd4; a_sign1 = 4'd12; a_sign2 = 4'd10; a_sign3 = 4'd11;
b_sign0 = 4'd3; b_sign1 = 4'd3; b_sign2 = 4'd2; b_sign3 = 4'd8;
@(posedge clk_i);
a_mant0 = 8'd114; a_mant1 = 8'd35; a_mant2 = 8'd221; a_mant3 = 8'd251;
b_mant0 = 8'd142; b_mant1 = 8'd5; b_mant2 = 8'd144; b_mant3 = 8'd106;
a_exp0 = 10'd160; a_exp1 = 10'd155; a_exp2 = 10'd888; a_exp3 = 10'd300;
b_exp0 = 10'd546; b_exp1 = 10'd188; b_exp2 = 10'd234; b_exp3 = 10'd617;
a_sign0 = 4'd12; a_sign1 = 4'd11; a_sign2 = 4'd5; a_sign3 = 4'd14;
b_sign0 = 4'd13; b_sign1 = 4'd4; b_sign2 = 4'd7; b_sign3 = 4'd9;
@(posedge clk_i);
a_mant0 = 8'd64; a_mant1 = 8'd93; a_mant2 = 8'd34; a_mant3 = 8'd91;
b_mant0 = 8'd80; b_mant1 = 8'd188; b_mant2 = 8'd238; b_mant3 = 8'd143;
a_exp0 = 10'd958; a_exp1 = 10'd752; a_exp2 = 10'd959; a_exp3 = 10'd917;
b_exp0 = 10'd532; b_exp1 = 10'd165; b_exp2 = 10'd347; b_exp3 = 10'd776;
a_sign0 = 4'd11; a_sign1 = 4'd10; a_sign2 = 4'd13; a_sign3 = 4'd8;
b_sign0 = 4'd9; b_sign1 = 4'd8; b_sign2 = 4'd14; b_sign3 = 4'd2;
@(posedge clk_i);
a_mant0 = 8'd95; a_mant1 = 8'd6; a_mant2 = 8'd221; a_mant3 = 8'd254;
b_mant0 = 8'd130; b_mant1 = 8'd138; b_mant2 = 8'd89; b_mant3 = 8'd1;
a_exp0 = 10'd347; a_exp1 = 10'd530; a_exp2 = 10'd735; a_exp3 = 10'd255;
b_exp0 = 10'd276; b_exp1 = 10'd343; b_exp2 = 10'd651; b_exp3 = 10'd245;
a_sign0 = 4'd3; a_sign1 = 4'd11; a_sign2 = 4'd8; a_sign3 = 4'd5;
b_sign0 = 4'd4; b_sign1 = 4'd7; b_sign2 = 4'd1; b_sign3 = 4'd12;
@(posedge clk_i);
shared_exps0 = 8'd117;
shared_exps1 = 8'd148;
a_mant0 = 8'd200; a_mant1 = 8'd190; a_mant2 = 8'd124; a_mant3 = 8'd157;
b_mant0 = 8'd116; b_mant1 = 8'd196; b_mant2 = 8'd227; b_mant3 = 8'd77;
a_exp0 = 10'd498; a_exp1 = 10'd706; a_exp2 = 10'd825; a_exp3 = 10'd877;
b_exp0 = 10'd780; b_exp1 = 10'd505; b_exp2 = 10'd348; b_exp3 = 10'd586;
a_sign0 = 4'd8; a_sign1 = 4'd16; a_sign2 = 4'd5; a_sign3 = 4'd14;
b_sign0 = 4'd8; b_sign1 = 4'd11; b_sign2 = 4'd2; b_sign3 = 4'd5;
@(posedge clk_i);
a_mant0 = 8'd183; a_mant1 = 8'd11; a_mant2 = 8'd169; a_mant3 = 8'd196;
b_mant0 = 8'd98; b_mant1 = 8'd193; b_mant2 = 8'd110; b_mant3 = 8'd99;
a_exp0 = 10'd695; a_exp1 = 10'd302; a_exp2 = 10'd198; a_exp3 = 10'd252;
b_exp0 = 10'd599; b_exp1 = 10'd1021; b_exp2 = 10'd670; b_exp3 = 10'd904;
a_sign0 = 4'd13; a_sign1 = 4'd4; a_sign2 = 4'd3; a_sign3 = 4'd11;
b_sign0 = 4'd4; b_sign1 = 4'd16; b_sign2 = 4'd6; b_sign3 = 4'd13;
@(posedge clk_i);
a_mant0 = 8'd69; a_mant1 = 8'd122; a_mant2 = 8'd165; a_mant3 = 8'd221;
b_mant0 = 8'd121; b_mant1 = 8'd105; b_mant2 = 8'd132; b_mant3 = 8'd177;
a_exp0 = 10'd123; a_exp1 = 10'd437; a_exp2 = 10'd107; a_exp3 = 10'd841;
b_exp0 = 10'd122; b_exp1 = 10'd739; b_exp2 = 10'd592; b_exp3 = 10'd943;
a_sign0 = 4'd6; a_sign1 = 4'd6; a_sign2 = 4'd7; a_sign3 = 4'd16;
b_sign0 = 4'd9; b_sign1 = 4'd1; b_sign2 = 4'd5; b_sign3 = 4'd16;
@(posedge clk_i);
a_mant0 = 8'd55; a_mant1 = 8'd4; a_mant2 = 8'd211; a_mant3 = 8'd113;
b_mant0 = 8'd129; b_mant1 = 8'd55; b_mant2 = 8'd224; b_mant3 = 8'd183;
a_exp0 = 10'd151; a_exp1 = 10'd237; a_exp2 = 10'd957; a_exp3 = 10'd445;
b_exp0 = 10'd408; b_exp1 = 10'd535; b_exp2 = 10'd919; b_exp3 = 10'd83;
a_sign0 = 4'd13; a_sign1 = 4'd7; a_sign2 = 4'd10; a_sign3 = 4'd3;
b_sign0 = 4'd7; b_sign1 = 4'd3; b_sign2 = 4'd11; b_sign3 = 4'd7;
@(posedge clk_i);
a_mant0 = 8'd226; a_mant1 = 8'd68; a_mant2 = 8'd149; a_mant3 = 8'd240;
b_mant0 = 8'd43; b_mant1 = 8'd0; b_mant2 = 8'd176; b_mant3 = 8'd58;
a_exp0 = 10'd657; a_exp1 = 10'd595; a_exp2 = 10'd988; a_exp3 = 10'd264;
b_exp0 = 10'd872; b_exp1 = 10'd409; b_exp2 = 10'd458; b_exp3 = 10'd740;
a_sign0 = 4'd16; a_sign1 = 4'd11; a_sign2 = 4'd16; a_sign3 = 4'd1;
b_sign0 = 4'd9; b_sign1 = 4'd14; b_sign2 = 4'd0; b_sign3 = 4'd4;
@(posedge clk_i);
a_mant0 = 8'd87; a_mant1 = 8'd151; a_mant2 = 8'd185; a_mant3 = 8'd112;
b_mant0 = 8'd231; b_mant1 = 8'd237; b_mant2 = 8'd70; b_mant3 = 8'd30;
a_exp0 = 10'd126; a_exp1 = 10'd38; a_exp2 = 10'd351; a_exp3 = 10'd957;
b_exp0 = 10'd404; b_exp1 = 10'd734; b_exp2 = 10'd65; b_exp3 = 10'd852;
a_sign0 = 4'd8; a_sign1 = 4'd10; a_sign2 = 4'd13; a_sign3 = 4'd15;
b_sign0 = 4'd7; b_sign1 = 4'd2; b_sign2 = 4'd7; b_sign3 = 4'd0;
@(posedge clk_i);
a_mant0 = 8'd73; a_mant1 = 8'd91; a_mant2 = 8'd57; a_mant3 = 8'd57;
b_mant0 = 8'd62; b_mant1 = 8'd246; b_mant2 = 8'd203; b_mant3 = 8'd56;
a_exp0 = 10'd896; a_exp1 = 10'd665; a_exp2 = 10'd68; a_exp3 = 10'd943;
b_exp0 = 10'd19; b_exp1 = 10'd414; b_exp2 = 10'd368; b_exp3 = 10'd766;
a_sign0 = 4'd1; a_sign1 = 4'd6; a_sign2 = 4'd6; a_sign3 = 4'd4;
b_sign0 = 4'd5; b_sign1 = 4'd15; b_sign2 = 4'd7; b_sign3 = 4'd0;
@(posedge clk_i);
a_mant0 = 8'd156; a_mant1 = 8'd103; a_mant2 = 8'd27; a_mant3 = 8'd27;
b_mant0 = 8'd250; b_mant1 = 8'd82; b_mant2 = 8'd61; b_mant3 = 8'd147;
a_exp0 = 10'd962; a_exp1 = 10'd45; a_exp2 = 10'd149; a_exp3 = 10'd1021;
b_exp0 = 10'd1001; b_exp1 = 10'd352; b_exp2 = 10'd777; b_exp3 = 10'd416;
a_sign0 = 4'd12; a_sign1 = 4'd5; a_sign2 = 4'd6; a_sign3 = 4'd1;
b_sign0 = 4'd6; b_sign1 = 4'd6; b_sign2 = 4'd4; b_sign3 = 4'd0;
@(posedge clk_i);
shared_exps0 = 8'd99;
shared_exps1 = 8'd119;
a_mant0 = 8'd109; a_mant1 = 8'd221; a_mant2 = 8'd80; a_mant3 = 8'd65;
b_mant0 = 8'd82; b_mant1 = 8'd129; b_mant2 = 8'd168; b_mant3 = 8'd7;
a_exp0 = 10'd611; a_exp1 = 10'd837; a_exp2 = 10'd251; a_exp3 = 10'd755;
b_exp0 = 10'd82; b_exp1 = 10'd126; b_exp2 = 10'd733; b_exp3 = 10'd15;
a_sign0 = 4'd6; a_sign1 = 4'd3; a_sign2 = 4'd2; a_sign3 = 4'd10;
b_sign0 = 4'd5; b_sign1 = 4'd5; b_sign2 = 4'd9; b_sign3 = 4'd5;
@(posedge clk_i);
a_mant0 = 8'd6; a_mant1 = 8'd147; a_mant2 = 8'd72; a_mant3 = 8'd20;
b_mant0 = 8'd38; b_mant1 = 8'd125; b_mant2 = 8'd95; b_mant3 = 8'd169;
a_exp0 = 10'd926; a_exp1 = 10'd187; a_exp2 = 10'd737; a_exp3 = 10'd942;
b_exp0 = 10'd122; b_exp1 = 10'd319; b_exp2 = 10'd765; b_exp3 = 10'd609;
a_sign0 = 4'd7; a_sign1 = 4'd14; a_sign2 = 4'd15; a_sign3 = 4'd8;
b_sign0 = 4'd11; b_sign1 = 4'd4; b_sign2 = 4'd1; b_sign3 = 4'd16;
@(posedge clk_i);
a_mant0 = 8'd54; a_mant1 = 8'd21; a_mant2 = 8'd207; a_mant3 = 8'd14;
b_mant0 = 8'd139; b_mant1 = 8'd56; b_mant2 = 8'd192; b_mant3 = 8'd43;
a_exp0 = 10'd339; a_exp1 = 10'd290; a_exp2 = 10'd424; a_exp3 = 10'd713;
b_exp0 = 10'd730; b_exp1 = 10'd171; b_exp2 = 10'd320; b_exp3 = 10'd117;
a_sign0 = 4'd7; a_sign1 = 4'd6; a_sign2 = 4'd2; a_sign3 = 4'd10;
b_sign0 = 4'd3; b_sign1 = 4'd0; b_sign2 = 4'd6; b_sign3 = 4'd8;
@(posedge clk_i);
a_mant0 = 8'd91; a_mant1 = 8'd172; a_mant2 = 8'd181; a_mant3 = 8'd55;
b_mant0 = 8'd238; b_mant1 = 8'd155; b_mant2 = 8'd111; b_mant3 = 8'd73;
a_exp0 = 10'd684; a_exp1 = 10'd36; a_exp2 = 10'd951; a_exp3 = 10'd444;
b_exp0 = 10'd275; b_exp1 = 10'd886; b_exp2 = 10'd72; b_exp3 = 10'd90;
a_sign0 = 4'd14; a_sign1 = 4'd15; a_sign2 = 4'd12; a_sign3 = 4'd2;
b_sign0 = 4'd15; b_sign1 = 4'd15; b_sign2 = 4'd12; b_sign3 = 4'd9;
@(posedge clk_i);
a_mant0 = 8'd36; a_mant1 = 8'd152; a_mant2 = 8'd170; a_mant3 = 8'd191;
b_mant0 = 8'd86; b_mant1 = 8'd115; b_mant2 = 8'd13; b_mant3 = 8'd14;
a_exp0 = 10'd814; a_exp1 = 10'd583; a_exp2 = 10'd425; a_exp3 = 10'd6;
b_exp0 = 10'd779; b_exp1 = 10'd1000; b_exp2 = 10'd478; b_exp3 = 10'd676;
a_sign0 = 4'd5; a_sign1 = 4'd12; a_sign2 = 4'd5; a_sign3 = 4'd11;
b_sign0 = 4'd4; b_sign1 = 4'd12; b_sign2 = 4'd4; b_sign3 = 4'd10;
@(posedge clk_i);
a_mant0 = 8'd29; a_mant1 = 8'd174; a_mant2 = 8'd133; a_mant3 = 8'd160;
b_mant0 = 8'd65; b_mant1 = 8'd106; b_mant2 = 8'd18; b_mant3 = 8'd224;
a_exp0 = 10'd76; a_exp1 = 10'd96; a_exp2 = 10'd167; a_exp3 = 10'd679;
b_exp0 = 10'd750; b_exp1 = 10'd15; b_exp2 = 10'd274; b_exp3 = 10'd481;
a_sign0 = 4'd3; a_sign1 = 4'd2; a_sign2 = 4'd16; a_sign3 = 4'd9;
b_sign0 = 4'd16; b_sign1 = 4'd4; b_sign2 = 4'd11; b_sign3 = 4'd16;
@(posedge clk_i);
a_mant0 = 8'd228; a_mant1 = 8'd159; a_mant2 = 8'd78; a_mant3 = 8'd253;
b_mant0 = 8'd58; b_mant1 = 8'd237; b_mant2 = 8'd11; b_mant3 = 8'd237;
a_exp0 = 10'd526; a_exp1 = 10'd872; a_exp2 = 10'd47; a_exp3 = 10'd199;
b_exp0 = 10'd12; b_exp1 = 10'd875; b_exp2 = 10'd558; b_exp3 = 10'd282;
a_sign0 = 4'd10; a_sign1 = 4'd2; a_sign2 = 4'd15; a_sign3 = 4'd1;
b_sign0 = 4'd4; b_sign1 = 4'd4; b_sign2 = 4'd8; b_sign3 = 4'd0;
@(posedge clk_i);
a_mant0 = 8'd124; a_mant1 = 8'd157; a_mant2 = 8'd219; a_mant3 = 8'd163;
b_mant0 = 8'd131; b_mant1 = 8'd254; b_mant2 = 8'd131; b_mant3 = 8'd185;
a_exp0 = 10'd13; a_exp1 = 10'd875; a_exp2 = 10'd105; a_exp3 = 10'd421;
b_exp0 = 10'd188; b_exp1 = 10'd218; b_exp2 = 10'd544; b_exp3 = 10'd650;
a_sign0 = 4'd6; a_sign1 = 4'd8; a_sign2 = 4'd11; a_sign3 = 4'd16;
b_sign0 = 4'd13; b_sign1 = 4'd2; b_sign2 = 4'd9; b_sign3 = 4'd7;
@(posedge clk_i);
shared_exps0 = 8'd120;
shared_exps1 = 8'd134;
rstn = 0;
@(posedge clk_i);
rstn = 1;
a_mant0 = 8'd225; a_mant1 = 8'd22; a_mant2 = 8'd41; a_mant3 = 8'd102;
b_mant0 = 8'd32; b_mant1 = 8'd175; b_mant2 = 8'd143; b_mant3 = 8'd236;
a_exp0 = 10'd793; a_exp1 = 10'd620; a_exp2 = 10'd682; a_exp3 = 10'd940;
b_exp0 = 10'd687; b_exp1 = 10'd148; b_exp2 = 10'd537; b_exp3 = 10'd309;
a_sign0 = 4'd16; a_sign1 = 4'd2; a_sign2 = 4'd13; a_sign3 = 4'd16;
b_sign0 = 4'd12; b_sign1 = 4'd7; b_sign2 = 4'd7; b_sign3 = 4'd1;
@(posedge clk_i);
a_mant0 = 8'd100; a_mant1 = 8'd128; a_mant2 = 8'd226; a_mant3 = 8'd142;
b_mant0 = 8'd114; b_mant1 = 8'd193; b_mant2 = 8'd152; b_mant3 = 8'd160;
a_exp0 = 10'd174; a_exp1 = 10'd403; a_exp2 = 10'd456; a_exp3 = 10'd712;
b_exp0 = 10'd147; b_exp1 = 10'd172; b_exp2 = 10'd756; b_exp3 = 10'd983;
a_sign0 = 4'd0; a_sign1 = 4'd7; a_sign2 = 4'd12; a_sign3 = 4'd16;
b_sign0 = 4'd2; b_sign1 = 4'd10; b_sign2 = 4'd4; b_sign3 = 4'd15;
@(posedge clk_i);
a_mant0 = 8'd67; a_mant1 = 8'd125; a_mant2 = 8'd185; a_mant3 = 8'd190;
b_mant0 = 8'd24; b_mant1 = 8'd85; b_mant2 = 8'd110; b_mant3 = 8'd147;
a_exp0 = 10'd504; a_exp1 = 10'd1002; a_exp2 = 10'd52; a_exp3 = 10'd510;
b_exp0 = 10'd838; b_exp1 = 10'd130; b_exp2 = 10'd77; b_exp3 = 10'd900;
a_sign0 = 4'd16; a_sign1 = 4'd4; a_sign2 = 4'd9; a_sign3 = 4'd1;
b_sign0 = 4'd14; b_sign1 = 4'd11; b_sign2 = 4'd0; b_sign3 = 4'd0;
@(posedge clk_i);
a_mant0 = 8'd90; a_mant1 = 8'd237; a_mant2 = 8'd106; a_mant3 = 8'd154;
b_mant0 = 8'd203; b_mant1 = 8'd34; b_mant2 = 8'd151; b_mant3 = 8'd91;
a_exp0 = 10'd474; a_exp1 = 10'd745; a_exp2 = 10'd116; a_exp3 = 10'd310;
b_exp0 = 10'd431; b_exp1 = 10'd736; b_exp2 = 10'd359; b_exp3 = 10'd425;
a_sign0 = 4'd12; a_sign1 = 4'd4; a_sign2 = 4'd15; a_sign3 = 4'd0;
b_sign0 = 4'd3; b_sign1 = 4'd16; b_sign2 = 4'd15; b_sign3 = 4'd8;
@(posedge clk_i);
a_mant0 = 8'd8; a_mant1 = 8'd84; a_mant2 = 8'd42; a_mant3 = 8'd192;
b_mant0 = 8'd218; b_mant1 = 8'd8; b_mant2 = 8'd119; b_mant3 = 8'd164;
a_exp0 = 10'd759; a_exp1 = 10'd151; a_exp2 = 10'd680; a_exp3 = 10'd884;
b_exp0 = 10'd168; b_exp1 = 10'd192; b_exp2 = 10'd619; b_exp3 = 10'd623;
a_sign0 = 4'd12; a_sign1 = 4'd9; a_sign2 = 4'd9; a_sign3 = 4'd8;
b_sign0 = 4'd4; b_sign1 = 4'd16; b_sign2 = 4'd0; b_sign3 = 4'd0;
@(posedge clk_i);
a_mant0 = 8'd183; a_mant1 = 8'd186; a_mant2 = 8'd9; a_mant3 = 8'd69;
b_mant0 = 8'd80; b_mant1 = 8'd74; b_mant2 = 8'd13; b_mant3 = 8'd21;
a_exp0 = 10'd167; a_exp1 = 10'd783; a_exp2 = 10'd152; a_exp3 = 10'd782;
b_exp0 = 10'd892; b_exp1 = 10'd101; b_exp2 = 10'd438; b_exp3 = 10'd391;
a_sign0 = 4'd10; a_sign1 = 4'd1; a_sign2 = 4'd0; a_sign3 = 4'd10;
b_sign0 = 4'd11; b_sign1 = 4'd16; b_sign2 = 4'd4; b_sign3 = 4'd15;
@(posedge clk_i);
a_mant0 = 8'd232; a_mant1 = 8'd68; a_mant2 = 8'd52; a_mant3 = 8'd201;
b_mant0 = 8'd5; b_mant1 = 8'd125; b_mant2 = 8'd18; b_mant3 = 8'd154;
a_exp0 = 10'd360; a_exp1 = 10'd835; a_exp2 = 10'd910; a_exp3 = 10'd366;
b_exp0 = 10'd901; b_exp1 = 10'd735; b_exp2 = 10'd580; b_exp3 = 10'd270;
a_sign0 = 4'd14; a_sign1 = 4'd14; a_sign2 = 4'd8; a_sign3 = 4'd4;
b_sign0 = 4'd1; b_sign1 = 4'd14; b_sign2 = 4'd14; b_sign3 = 4'd2;
@(posedge clk_i);
shared_exps0 = 8'd113;
shared_exps1 = 8'd161;
a_mant0 = 8'd116; a_mant1 = 8'd248; a_mant2 = 8'd12; a_mant3 = 8'd134;
b_mant0 = 8'd26; b_mant1 = 8'd131; b_mant2 = 8'd56; b_mant3 = 8'd96;
a_exp0 = 10'd509; a_exp1 = 10'd339; a_exp2 = 10'd1; a_exp3 = 10'd857;
b_exp0 = 10'd736; b_exp1 = 10'd329; b_exp2 = 10'd680; b_exp3 = 10'd536;
a_sign0 = 4'd9; a_sign1 = 4'd7; a_sign2 = 4'd11; a_sign3 = 4'd3;
b_sign0 = 4'd4; b_sign1 = 4'd5; b_sign2 = 4'd12; b_sign3 = 4'd6;
@(posedge clk_i);
a_mant0 = 8'd50; a_mant1 = 8'd160; a_mant2 = 8'd29; a_mant3 = 8'd93;
b_mant0 = 8'd74; b_mant1 = 8'd103; b_mant2 = 8'd84; b_mant3 = 8'd157;
a_exp0 = 10'd702; a_exp1 = 10'd933; a_exp2 = 10'd568; a_exp3 = 10'd739;
b_exp0 = 10'd1; b_exp1 = 10'd841; b_exp2 = 10'd868; b_exp3 = 10'd338;
a_sign0 = 4'd5; a_sign1 = 4'd16; a_sign2 = 4'd16; a_sign3 = 4'd14;
b_sign0 = 4'd12; b_sign1 = 4'd4; b_sign2 = 4'd16; b_sign3 = 4'd5;
@(posedge clk_i);
a_mant0 = 8'd180; a_mant1 = 8'd70; a_mant2 = 8'd92; a_mant3 = 8'd199;
b_mant0 = 8'd215; b_mant1 = 8'd46; b_mant2 = 8'd43; b_mant3 = 8'd22;
a_exp0 = 10'd633; a_exp1 = 10'd972; a_exp2 = 10'd286; a_exp3 = 10'd406;
b_exp0 = 10'd174; b_exp1 = 10'd500; b_exp2 = 10'd473; b_exp3 = 10'd789;
a_sign0 = 4'd3; a_sign1 = 4'd5; a_sign2 = 4'd2; a_sign3 = 4'd7;
b_sign0 = 4'd16; b_sign1 = 4'd1; b_sign2 = 4'd2; b_sign3 = 4'd0;
@(posedge clk_i);
a_mant0 = 8'd47; a_mant1 = 8'd173; a_mant2 = 8'd67; a_mant3 = 8'd64;
b_mant0 = 8'd224; b_mant1 = 8'd62; b_mant2 = 8'd18; b_mant3 = 8'd254;
a_exp0 = 10'd464; a_exp1 = 10'd848; a_exp2 = 10'd868; a_exp3 = 10'd45;
b_exp0 = 10'd263; b_exp1 = 10'd917; b_exp2 = 10'd832; b_exp3 = 10'd633;
a_sign0 = 4'd10; a_sign1 = 4'd9; a_sign2 = 4'd3; a_sign3 = 4'd6;
b_sign0 = 4'd11; b_sign1 = 4'd5; b_sign2 = 4'd3; b_sign3 = 4'd6;
@(posedge clk_i);
a_mant0 = 8'd9; a_mant1 = 8'd192; a_mant2 = 8'd188; a_mant3 = 8'd197;
b_mant0 = 8'd160; b_mant1 = 8'd221; b_mant2 = 8'd132; b_mant3 = 8'd94;
a_exp0 = 10'd55; a_exp1 = 10'd188; a_exp2 = 10'd954; a_exp3 = 10'd137;
b_exp0 = 10'd439; b_exp1 = 10'd563; b_exp2 = 10'd951; b_exp3 = 10'd661;
a_sign0 = 4'd13; a_sign1 = 4'd15; a_sign2 = 4'd0; a_sign3 = 4'd5;
b_sign0 = 4'd11; b_sign1 = 4'd4; b_sign2 = 4'd5; b_sign3 = 4'd13;
@(posedge clk_i);
a_mant0 = 8'd108; a_mant1 = 8'd83; a_mant2 = 8'd182; a_mant3 = 8'd195;
b_mant0 = 8'd52; b_mant1 = 8'd19; b_mant2 = 8'd100; b_mant3 = 8'd0;
a_exp0 = 10'd722; a_exp1 = 10'd212; a_exp2 = 10'd1005; a_exp3 = 10'd292;
b_exp0 = 10'd855; b_exp1 = 10'd222; b_exp2 = 10'd833; b_exp3 = 10'd0;
a_sign0 = 4'd2; a_sign1 = 4'd16; a_sign2 = 4'd2; a_sign3 = 4'd15;
b_sign0 = 4'd1; b_sign1 = 4'd10; b_sign2 = 4'd2; b_sign3 = 4'd15;
@(posedge clk_i);
a_mant0 = 8'd83; a_mant1 = 8'd67; a_mant2 = 8'd40; a_mant3 = 8'd202;
b_mant0 = 8'd11; b_mant1 = 8'd173; b_mant2 = 8'd18; b_mant3 = 8'd107;
a_exp0 = 10'd747; a_exp1 = 10'd617; a_exp2 = 10'd677; a_exp3 = 10'd240;
b_exp0 = 10'd532; b_exp1 = 10'd454; b_exp2 = 10'd371; b_exp3 = 10'd806;
a_sign0 = 4'd0; a_sign1 = 4'd16; a_sign2 = 4'd4; a_sign3 = 4'd4;
b_sign0 = 4'd3; b_sign1 = 4'd4; b_sign2 = 4'd0; b_sign3 = 4'd4;
@(posedge clk_i);
a_mant0 = 8'd220; a_mant1 = 8'd247; a_mant2 = 8'd47; a_mant3 = 8'd223;
b_mant0 = 8'd151; b_mant1 = 8'd243; b_mant2 = 8'd121; b_mant3 = 8'd247;
a_exp0 = 10'd211; a_exp1 = 10'd952; a_exp2 = 10'd553; a_exp3 = 10'd106;
b_exp0 = 10'd281; b_exp1 = 10'd244; b_exp2 = 10'd1020; b_exp3 = 10'd100;
a_sign0 = 4'd10; a_sign1 = 4'd2; a_sign2 = 4'd5; a_sign3 = 4'd14;
b_sign0 = 4'd4; b_sign1 = 4'd4; b_sign2 = 4'd12; b_sign3 = 4'd8;
@(posedge clk_i);
shared_exps0 = 8'd123;
shared_exps1 = 8'd123;
a_mant0 = 8'd42; a_mant1 = 8'd194; a_mant2 = 8'd187; a_mant3 = 8'd220;
b_mant0 = 8'd195; b_mant1 = 8'd144; b_mant2 = 8'd225; b_mant3 = 8'd240;
a_exp0 = 10'd330; a_exp1 = 10'd60; a_exp2 = 10'd720; a_exp3 = 10'd761;
b_exp0 = 10'd250; b_exp1 = 10'd168; b_exp2 = 10'd524; b_exp3 = 10'd964;
a_sign0 = 4'd0; a_sign1 = 4'd5; a_sign2 = 4'd5; a_sign3 = 4'd12;
b_sign0 = 4'd3; b_sign1 = 4'd2; b_sign2 = 4'd12; b_sign3 = 4'd2;
@(posedge clk_i);
a_mant0 = 8'd166; a_mant1 = 8'd0; a_mant2 = 8'd55; a_mant3 = 8'd206;
b_mant0 = 8'd162; b_mant1 = 8'd206; b_mant2 = 8'd151; b_mant3 = 8'd206;
a_exp0 = 10'd77; a_exp1 = 10'd520; a_exp2 = 10'd359; a_exp3 = 10'd34;
b_exp0 = 10'd134; b_exp1 = 10'd38; b_exp2 = 10'd699; b_exp3 = 10'd976;
a_sign0 = 4'd5; a_sign1 = 4'd10; a_sign2 = 4'd14; a_sign3 = 4'd11;
b_sign0 = 4'd10; b_sign1 = 4'd5; b_sign2 = 4'd4; b_sign3 = 4'd2;
@(posedge clk_i);
a_mant0 = 8'd189; a_mant1 = 8'd194; a_mant2 = 8'd200; a_mant3 = 8'd4;
b_mant0 = 8'd102; b_mant1 = 8'd235; b_mant2 = 8'd29; b_mant3 = 8'd103;
a_exp0 = 10'd14; a_exp1 = 10'd105; a_exp2 = 10'd738; a_exp3 = 10'd37;
b_exp0 = 10'd838; b_exp1 = 10'd139; b_exp2 = 10'd139; b_exp3 = 10'd1011;
a_sign0 = 4'd5; a_sign1 = 4'd9; a_sign2 = 4'd7; a_sign3 = 4'd4;
b_sign0 = 4'd4; b_sign1 = 4'd7; b_sign2 = 4'd14; b_sign3 = 4'd12;
@(posedge clk_i);
a_mant0 = 8'd61; a_mant1 = 8'd200; a_mant2 = 8'd243; a_mant3 = 8'd44;
b_mant0 = 8'd33; b_mant1 = 8'd152; b_mant2 = 8'd111; b_mant3 = 8'd244;
a_exp0 = 10'd209; a_exp1 = 10'd773; a_exp2 = 10'd189; a_exp3 = 10'd515;
b_exp0 = 10'd442; b_exp1 = 10'd919; b_exp2 = 10'd575; b_exp3 = 10'd886;
a_sign0 = 4'd13; a_sign1 = 4'd14; a_sign2 = 4'd5; a_sign3 = 4'd16;
b_sign0 = 4'd4; b_sign1 = 4'd16; b_sign2 = 4'd8; b_sign3 = 4'd10;
@(posedge clk_i);
a_mant0 = 8'd55; a_mant1 = 8'd117; a_mant2 = 8'd66; a_mant3 = 8'd210;
b_mant0 = 8'd47; b_mant1 = 8'd220; b_mant2 = 8'd37; b_mant3 = 8'd97;
a_exp0 = 10'd942; a_exp1 = 10'd552; a_exp2 = 10'd437; a_exp3 = 10'd509;
b_exp0 = 10'd405; b_exp1 = 10'd266; b_exp2 = 10'd948; b_exp3 = 10'd574;
a_sign0 = 4'd14; a_sign1 = 4'd6; a_sign2 = 4'd9; a_sign3 = 4'd7;
b_sign0 = 4'd3; b_sign1 = 4'd8; b_sign2 = 4'd12; b_sign3 = 4'd16;
@(posedge clk_i);
a_mant0 = 8'd47; a_mant1 = 8'd226; a_mant2 = 8'd148; a_mant3 = 8'd207;
b_mant0 = 8'd149; b_mant1 = 8'd243; b_mant2 = 8'd31; b_mant3 = 8'd253;
a_exp0 = 10'd945; a_exp1 = 10'd445; a_exp2 = 10'd715; a_exp3 = 10'd506;
b_exp0 = 10'd775; b_exp1 = 10'd778; b_exp2 = 10'd683; b_exp3 = 10'd5;
a_sign0 = 4'd0; a_sign1 = 4'd16; a_sign2 = 4'd8; a_sign3 = 4'd3;
b_sign0 = 4'd15; b_sign1 = 4'd13; b_sign2 = 4'd3; b_sign3 = 4'd1;
@(posedge clk_i);
a_mant0 = 8'd145; a_mant1 = 8'd15; a_mant2 = 8'd99; a_mant3 = 8'd37;
b_mant0 = 8'd250; b_mant1 = 8'd56; b_mant2 = 8'd163; b_mant3 = 8'd240;
a_exp0 = 10'd200; a_exp1 = 10'd231; a_exp2 = 10'd645; a_exp3 = 10'd22;
b_exp0 = 10'd533; b_exp1 = 10'd928; b_exp2 = 10'd643; b_exp3 = 10'd802;
a_sign0 = 4'd8; a_sign1 = 4'd9; a_sign2 = 4'd9; a_sign3 = 4'd16;
b_sign0 = 4'd0; b_sign1 = 4'd2; b_sign2 = 4'd16; b_sign3 = 4'd12;
@(posedge clk_i);
a_mant0 = 8'd3; a_mant1 = 8'd226; a_mant2 = 8'd183; a_mant3 = 8'd255;
b_mant0 = 8'd220; b_mant1 = 8'd165; b_mant2 = 8'd8; b_mant3 = 8'd58;
a_exp0 = 10'd608; a_exp1 = 10'd752; a_exp2 = 10'd295; a_exp3 = 10'd458;
b_exp0 = 10'd322; b_exp1 = 10'd526; b_exp2 = 10'd788; b_exp3 = 10'd246;
a_sign0 = 4'd1; a_sign1 = 4'd3; a_sign2 = 4'd4; a_sign3 = 4'd3;
b_sign0 = 4'd10; b_sign1 = 4'd1; b_sign2 = 4'd11; b_sign3 = 4'd5;
@(posedge clk_i);
shared_exps0 = 8'd138;
shared_exps1 = 8'd104;
a_mant0 = 8'd59; a_mant1 = 8'd58; a_mant2 = 8'd170; a_mant3 = 8'd55;
b_mant0 = 8'd11; b_mant1 = 8'd40; b_mant2 = 8'd75; b_mant3 = 8'd161;
a_exp0 = 10'd275; a_exp1 = 10'd989; a_exp2 = 10'd68; a_exp3 = 10'd838;
b_exp0 = 10'd59; b_exp1 = 10'd708; b_exp2 = 10'd136; b_exp3 = 10'd739;
a_sign0 = 4'd13; a_sign1 = 4'd11; a_sign2 = 4'd2; a_sign3 = 4'd11;
b_sign0 = 4'd10; b_sign1 = 4'd4; b_sign2 = 4'd9; b_sign3 = 4'd8;
@(posedge clk_i);
a_mant0 = 8'd242; a_mant1 = 8'd19; a_mant2 = 8'd214; a_mant3 = 8'd228;
b_mant0 = 8'd127; b_mant1 = 8'd42; b_mant2 = 8'd38; b_mant3 = 8'd19;
a_exp0 = 10'd1003; a_exp1 = 10'd761; a_exp2 = 10'd248; a_exp3 = 10'd207;
b_exp0 = 10'd990; b_exp1 = 10'd373; b_exp2 = 10'd161; b_exp3 = 10'd764;
a_sign0 = 4'd13; a_sign1 = 4'd12; a_sign2 = 4'd14; a_sign3 = 4'd13;
b_sign0 = 4'd1; b_sign1 = 4'd2; b_sign2 = 4'd6; b_sign3 = 4'd1;
@(posedge clk_i);
a_mant0 = 8'd200; a_mant1 = 8'd201; a_mant2 = 8'd229; a_mant3 = 8'd26;
b_mant0 = 8'd56; b_mant1 = 8'd82; b_mant2 = 8'd225; b_mant3 = 8'd194;
a_exp0 = 10'd322; a_exp1 = 10'd933; a_exp2 = 10'd850; a_exp3 = 10'd869;
b_exp0 = 10'd671; b_exp1 = 10'd187; b_exp2 = 10'd347; b_exp3 = 10'd375;
a_sign0 = 4'd5; a_sign1 = 4'd10; a_sign2 = 4'd6; a_sign3 = 4'd12;
b_sign0 = 4'd10; b_sign1 = 4'd13; b_sign2 = 4'd4; b_sign3 = 4'd13;
@(posedge clk_i);
a_mant0 = 8'd58; a_mant1 = 8'd24; a_mant2 = 8'd194; a_mant3 = 8'd90;
b_mant0 = 8'd50; b_mant1 = 8'd9; b_mant2 = 8'd104; b_mant3 = 8'd96;
a_exp0 = 10'd253; a_exp1 = 10'd552; a_exp2 = 10'd910; a_exp3 = 10'd763;
b_exp0 = 10'd539; b_exp1 = 10'd922; b_exp2 = 10'd202; b_exp3 = 10'd862;
a_sign0 = 4'd15; a_sign1 = 4'd13; a_sign2 = 4'd5; a_sign3 = 4'd15;
b_sign0 = 4'd15; b_sign1 = 4'd9; b_sign2 = 4'd5; b_sign3 = 4'd12;
@(posedge clk_i);
a_mant0 = 8'd178; a_mant1 = 8'd61; a_mant2 = 8'd113; a_mant3 = 8'd176;
b_mant0 = 8'd19; b_mant1 = 8'd46; b_mant2 = 8'd195; b_mant3 = 8'd49;
a_exp0 = 10'd990; a_exp1 = 10'd683; a_exp2 = 10'd395; a_exp3 = 10'd989;
b_exp0 = 10'd11; b_exp1 = 10'd260; b_exp2 = 10'd192; b_exp3 = 10'd374;
a_sign0 = 4'd2; a_sign1 = 4'd1; a_sign2 = 4'd5; a_sign3 = 4'd13;
b_sign0 = 4'd12; b_sign1 = 4'd14; b_sign2 = 4'd7; b_sign3 = 4'd14;
@(posedge clk_i);
a_mant0 = 8'd210; a_mant1 = 8'd68; a_mant2 = 8'd181; a_mant3 = 8'd210;
b_mant0 = 8'd42; b_mant1 = 8'd45; b_mant2 = 8'd52; b_mant3 = 8'd20;
a_exp0 = 10'd77; a_exp1 = 10'd750; a_exp2 = 10'd229; a_exp3 = 10'd0;
b_exp0 = 10'd794; b_exp1 = 10'd380; b_exp2 = 10'd1001; b_exp3 = 10'd183;
a_sign0 = 4'd14; a_sign1 = 4'd1; a_sign2 = 4'd12; a_sign3 = 4'd4;
b_sign0 = 4'd3; b_sign1 = 4'd9; b_sign2 = 4'd12; b_sign3 = 4'd8;
@(posedge clk_i);
a_mant0 = 8'd104; a_mant1 = 8'd114; a_mant2 = 8'd36; a_mant3 = 8'd205;
b_mant0 = 8'd118; b_mant1 = 8'd53; b_mant2 = 8'd75; b_mant3 = 8'd100;
a_exp0 = 10'd370; a_exp1 = 10'd485; a_exp2 = 10'd677; a_exp3 = 10'd647;
b_exp0 = 10'd921; b_exp1 = 10'd789; b_exp2 = 10'd178; b_exp3 = 10'd600;
a_sign0 = 4'd4; a_sign1 = 4'd10; a_sign2 = 4'd2; a_sign3 = 4'd13;
b_sign0 = 4'd7; b_sign1 = 4'd8; b_sign2 = 4'd7; b_sign3 = 4'd3;
@(posedge clk_i);
a_mant0 = 8'd81; a_mant1 = 8'd220; a_mant2 = 8'd32; a_mant3 = 8'd78;
b_mant0 = 8'd158; b_mant1 = 8'd100; b_mant2 = 8'd204; b_mant3 = 8'd167;
a_exp0 = 10'd221; a_exp1 = 10'd414; a_exp2 = 10'd496; a_exp3 = 10'd44;
b_exp0 = 10'd392; b_exp1 = 10'd133; b_exp2 = 10'd192; b_exp3 = 10'd1003;
a_sign0 = 4'd10; a_sign1 = 4'd8; a_sign2 = 4'd15; a_sign3 = 4'd11;
b_sign0 = 4'd5; b_sign1 = 4'd6; b_sign2 = 4'd14; b_sign3 = 4'd7;
@(posedge clk_i);
shared_exps0 = 8'd153;
shared_exps1 = 8'd138;
rstn = 0;
@(posedge clk_i);
rstn = 1;
a_mant0 = 8'd165; a_mant1 = 8'd191; a_mant2 = 8'd145; a_mant3 = 8'd93;
b_mant0 = 8'd114; b_mant1 = 8'd139; b_mant2 = 8'd112; b_mant3 = 8'd174;
a_exp0 = 10'd860; a_exp1 = 10'd798; a_exp2 = 10'd685; a_exp3 = 10'd740;
b_exp0 = 10'd905; b_exp1 = 10'd12; b_exp2 = 10'd215; b_exp3 = 10'd360;
a_sign0 = 4'd1; a_sign1 = 4'd11; a_sign2 = 4'd2; a_sign3 = 4'd2;
b_sign0 = 4'd3; b_sign1 = 4'd11; b_sign2 = 4'd3; b_sign3 = 4'd7;
@(posedge clk_i);
a_mant0 = 8'd181; a_mant1 = 8'd102; a_mant2 = 8'd127; a_mant3 = 8'd34;
b_mant0 = 8'd225; b_mant1 = 8'd86; b_mant2 = 8'd88; b_mant3 = 8'd61;
a_exp0 = 10'd129; a_exp1 = 10'd52; a_exp2 = 10'd229; a_exp3 = 10'd56;
b_exp0 = 10'd138; b_exp1 = 10'd1017; b_exp2 = 10'd721; b_exp3 = 10'd24;
a_sign0 = 4'd3; a_sign1 = 4'd5; a_sign2 = 4'd10; a_sign3 = 4'd11;
b_sign0 = 4'd6; b_sign1 = 4'd1; b_sign2 = 4'd4; b_sign3 = 4'd15;
@(posedge clk_i);
a_mant0 = 8'd13; a_mant1 = 8'd136; a_mant2 = 8'd2; a_mant3 = 8'd151;
b_mant0 = 8'd219; b_mant1 = 8'd98; b_mant2 = 8'd200; b_mant3 = 8'd166;
a_exp0 = 10'd523; a_exp1 = 10'd858; a_exp2 = 10'd62; a_exp3 = 10'd835;
b_exp0 = 10'd153; b_exp1 = 10'd90; b_exp2 = 10'd324; b_exp3 = 10'd110;
a_sign0 = 4'd7; a_sign1 = 4'd8; a_sign2 = 4'd0; a_sign3 = 4'd6;
b_sign0 = 4'd14; b_sign1 = 4'd0; b_sign2 = 4'd10; b_sign3 = 4'd5;
@(posedge clk_i);
a_mant0 = 8'd167; a_mant1 = 8'd11; a_mant2 = 8'd142; a_mant3 = 8'd112;
b_mant0 = 8'd231; b_mant1 = 8'd6; b_mant2 = 8'd231; b_mant3 = 8'd147;
a_exp0 = 10'd593; a_exp1 = 10'd120; a_exp2 = 10'd188; a_exp3 = 10'd71;
b_exp0 = 10'd426; b_exp1 = 10'd806; b_exp2 = 10'd788; b_exp3 = 10'd1012;
a_sign0 = 4'd0; a_sign1 = 4'd8; a_sign2 = 4'd9; a_sign3 = 4'd10;
b_sign0 = 4'd5; b_sign1 = 4'd15; b_sign2 = 4'd9; b_sign3 = 4'd4;
@(posedge clk_i);
a_mant0 = 8'd58; a_mant1 = 8'd107; a_mant2 = 8'd216; a_mant3 = 8'd227;
b_mant0 = 8'd1; b_mant1 = 8'd169; b_mant2 = 8'd89; b_mant3 = 8'd116;
a_exp0 = 10'd652; a_exp1 = 10'd597; a_exp2 = 10'd654; a_exp3 = 10'd104;
b_exp0 = 10'd431; b_exp1 = 10'd295; b_exp2 = 10'd938; b_exp3 = 10'd972;
a_sign0 = 4'd14; a_sign1 = 4'd5; a_sign2 = 4'd12; a_sign3 = 4'd5;
b_sign0 = 4'd2; b_sign1 = 4'd5; b_sign2 = 4'd8; b_sign3 = 4'd16;
@(posedge clk_i);
a_mant0 = 8'd30; a_mant1 = 8'd192; a_mant2 = 8'd3; a_mant3 = 8'd59;
b_mant0 = 8'd245; b_mant1 = 8'd50; b_mant2 = 8'd243; b_mant3 = 8'd107;
a_exp0 = 10'd975; a_exp1 = 10'd216; a_exp2 = 10'd201; a_exp3 = 10'd966;
b_exp0 = 10'd462; b_exp1 = 10'd457; b_exp2 = 10'd314; b_exp3 = 10'd844;
a_sign0 = 4'd7; a_sign1 = 4'd1; a_sign2 = 4'd15; a_sign3 = 4'd10;
b_sign0 = 4'd5; b_sign1 = 4'd0; b_sign2 = 4'd5; b_sign3 = 4'd9;
@(posedge clk_i);
a_mant0 = 8'd11; a_mant1 = 8'd11; a_mant2 = 8'd115; a_mant3 = 8'd178;
b_mant0 = 8'd253; b_mant1 = 8'd189; b_mant2 = 8'd97; b_mant3 = 8'd2;
a_exp0 = 10'd964; a_exp1 = 10'd866; a_exp2 = 10'd180; a_exp3 = 10'd847;
b_exp0 = 10'd412; b_exp1 = 10'd512; b_exp2 = 10'd458; b_exp3 = 10'd796;
a_sign0 = 4'd1; a_sign1 = 4'd15; a_sign2 = 4'd6; a_sign3 = 4'd11;
b_sign0 = 4'd7; b_sign1 = 4'd4; b_sign2 = 4'd13; b_sign3 = 4'd11;
@(posedge clk_i);
shared_exps0 = 8'd112;
shared_exps1 = 8'd109;
a_mant0 = 8'd16; a_mant1 = 8'd180; a_mant2 = 8'd234; a_mant3 = 8'd99;
b_mant0 = 8'd75; b_mant1 = 8'd90; b_mant2 = 8'd28; b_mant3 = 8'd219;
a_exp0 = 10'd1009; a_exp1 = 10'd757; a_exp2 = 10'd190; a_exp3 = 10'd246;
b_exp0 = 10'd741; b_exp1 = 10'd440; b_exp2 = 10'd112; b_exp3 = 10'd457;
a_sign0 = 4'd16; a_sign1 = 4'd15; a_sign2 = 4'd4; a_sign3 = 4'd2;
b_sign0 = 4'd16; b_sign1 = 4'd1; b_sign2 = 4'd10; b_sign3 = 4'd7;
@(posedge clk_i);
a_mant0 = 8'd139; a_mant1 = 8'd180; a_mant2 = 8'd157; a_mant3 = 8'd141;
b_mant0 = 8'd15; b_mant1 = 8'd25; b_mant2 = 8'd147; b_mant3 = 8'd9;
a_exp0 = 10'd786; a_exp1 = 10'd420; a_exp2 = 10'd259; a_exp3 = 10'd337;
b_exp0 = 10'd251; b_exp1 = 10'd506; b_exp2 = 10'd501; b_exp3 = 10'd466;
a_sign0 = 4'd12; a_sign1 = 4'd13; a_sign2 = 4'd0; a_sign3 = 4'd11;
b_sign0 = 4'd4; b_sign1 = 4'd14; b_sign2 = 4'd4; b_sign3 = 4'd13;
@(posedge clk_i);
a_mant0 = 8'd206; a_mant1 = 8'd183; a_mant2 = 8'd175; a_mant3 = 8'd149;
b_mant0 = 8'd179; b_mant1 = 8'd112; b_mant2 = 8'd34; b_mant3 = 8'd233;
a_exp0 = 10'd963; a_exp1 = 10'd868; a_exp2 = 10'd483; a_exp3 = 10'd369;
b_exp0 = 10'd368; b_exp1 = 10'd335; b_exp2 = 10'd676; b_exp3 = 10'd474;
a_sign0 = 4'd16; a_sign1 = 4'd10; a_sign2 = 4'd3; a_sign3 = 4'd0;
b_sign0 = 4'd5; b_sign1 = 4'd9; b_sign2 = 4'd5; b_sign3 = 4'd8;
@(posedge clk_i);
a_mant0 = 8'd47; a_mant1 = 8'd12; a_mant2 = 8'd254; a_mant3 = 8'd245;
b_mant0 = 8'd124; b_mant1 = 8'd24; b_mant2 = 8'd61; b_mant3 = 8'd113;
a_exp0 = 10'd38; a_exp1 = 10'd273; a_exp2 = 10'd546; a_exp3 = 10'd453;
b_exp0 = 10'd324; b_exp1 = 10'd341; b_exp2 = 10'd1011; b_exp3 = 10'd654;
a_sign0 = 4'd12; a_sign1 = 4'd10; a_sign2 = 4'd3; a_sign3 = 4'd11;
b_sign0 = 4'd14; b_sign1 = 4'd16; b_sign2 = 4'd12; b_sign3 = 4'd7;
@(posedge clk_i);
a_mant0 = 8'd183; a_mant1 = 8'd142; a_mant2 = 8'd56; a_mant3 = 8'd59;
b_mant0 = 8'd240; b_mant1 = 8'd172; b_mant2 = 8'd9; b_mant3 = 8'd88;
a_exp0 = 10'd533; a_exp1 = 10'd757; a_exp2 = 10'd588; a_exp3 = 10'd468;
b_exp0 = 10'd831; b_exp1 = 10'd374; b_exp2 = 10'd1019; b_exp3 = 10'd845;
a_sign0 = 4'd4; a_sign1 = 4'd16; a_sign2 = 4'd6; a_sign3 = 4'd1;
b_sign0 = 4'd10; b_sign1 = 4'd10; b_sign2 = 4'd6; b_sign3 = 4'd4;
@(posedge clk_i);
a_mant0 = 8'd82; a_mant1 = 8'd162; a_mant2 = 8'd114; a_mant3 = 8'd226;
b_mant0 = 8'd227; b_mant1 = 8'd202; b_mant2 = 8'd223; b_mant3 = 8'd156;
a_exp0 = 10'd974; a_exp1 = 10'd11; a_exp2 = 10'd43; a_exp3 = 10'd530;
b_exp0 = 10'd690; b_exp1 = 10'd531; b_exp2 = 10'd818; b_exp3 = 10'd786;
a_sign0 = 4'd12; a_sign1 = 4'd14; a_sign2 = 4'd15; a_sign3 = 4'd1;
b_sign0 = 4'd11; b_sign1 = 4'd15; b_sign2 = 4'd14; b_sign3 = 4'd0;
@(posedge clk_i);
a_mant0 = 8'd208; a_mant1 = 8'd178; a_mant2 = 8'd209; a_mant3 = 8'd185;
b_mant0 = 8'd207; b_mant1 = 8'd42; b_mant2 = 8'd242; b_mant3 = 8'd44;
a_exp0 = 10'd317; a_exp1 = 10'd768; a_exp2 = 10'd217; a_exp3 = 10'd828;
b_exp0 = 10'd566; b_exp1 = 10'd781; b_exp2 = 10'd109; b_exp3 = 10'd530;
a_sign0 = 4'd15; a_sign1 = 4'd9; a_sign2 = 4'd1; a_sign3 = 4'd4;
b_sign0 = 4'd1; b_sign1 = 4'd7; b_sign2 = 4'd0; b_sign3 = 4'd12;
@(posedge clk_i);
a_mant0 = 8'd119; a_mant1 = 8'd58; a_mant2 = 8'd215; a_mant3 = 8'd91;
b_mant0 = 8'd182; b_mant1 = 8'd253; b_mant2 = 8'd170; b_mant3 = 8'd178;
a_exp0 = 10'd177; a_exp1 = 10'd559; a_exp2 = 10'd763; a_exp3 = 10'd664;
b_exp0 = 10'd660; b_exp1 = 10'd795; b_exp2 = 10'd276; b_exp3 = 10'd702;
a_sign0 = 4'd4; a_sign1 = 4'd0; a_sign2 = 4'd16; a_sign3 = 4'd10;
b_sign0 = 4'd2; b_sign1 = 4'd1; b_sign2 = 4'd7; b_sign3 = 4'd3;
@(posedge clk_i);
shared_exps0 = 8'd111;
shared_exps1 = 8'd129;
a_mant0 = 8'd122; a_mant1 = 8'd57; a_mant2 = 8'd38; a_mant3 = 8'd18;
b_mant0 = 8'd245; b_mant1 = 8'd53; b_mant2 = 8'd99; b_mant3 = 8'd214;
a_exp0 = 10'd54; a_exp1 = 10'd448; a_exp2 = 10'd359; a_exp3 = 10'd744;
b_exp0 = 10'd184; b_exp1 = 10'd671; b_exp2 = 10'd859; b_exp3 = 10'd560;
a_sign0 = 4'd13; a_sign1 = 4'd16; a_sign2 = 4'd13; a_sign3 = 4'd2;
b_sign0 = 4'd3; b_sign1 = 4'd11; b_sign2 = 4'd2; b_sign3 = 4'd6;
@(posedge clk_i);
a_mant0 = 8'd165; a_mant1 = 8'd127; a_mant2 = 8'd109; a_mant3 = 8'd232;
b_mant0 = 8'd42; b_mant1 = 8'd159; b_mant2 = 8'd172; b_mant3 = 8'd113;
a_exp0 = 10'd180; a_exp1 = 10'd71; a_exp2 = 10'd1006; a_exp3 = 10'd77;
b_exp0 = 10'd706; b_exp1 = 10'd98; b_exp2 = 10'd799; b_exp3 = 10'd961;
a_sign0 = 4'd6; a_sign1 = 4'd11; a_sign2 = 4'd13; a_sign3 = 4'd16;
b_sign0 = 4'd14; b_sign1 = 4'd0; b_sign2 = 4'd2; b_sign3 = 4'd4;
@(posedge clk_i);
a_mant0 = 8'd40; a_mant1 = 8'd45; a_mant2 = 8'd171; a_mant3 = 8'd116;
b_mant0 = 8'd199; b_mant1 = 8'd200; b_mant2 = 8'd153; b_mant3 = 8'd89;
a_exp0 = 10'd781; a_exp1 = 10'd207; a_exp2 = 10'd911; a_exp3 = 10'd118;
b_exp0 = 10'd181; b_exp1 = 10'd251; b_exp2 = 10'd754; b_exp3 = 10'd528;
a_sign0 = 4'd8; a_sign1 = 4'd5; a_sign2 = 4'd8; a_sign3 = 4'd15;
b_sign0 = 4'd16; b_sign1 = 4'd6; b_sign2 = 4'd14; b_sign3 = 4'd13;
@(posedge clk_i);
a_mant0 = 8'd167; a_mant1 = 8'd144; a_mant2 = 8'd90; a_mant3 = 8'd18;
b_mant0 = 8'd26; b_mant1 = 8'd3; b_mant2 = 8'd99; b_mant3 = 8'd23;
a_exp0 = 10'd534; a_exp1 = 10'd296; a_exp2 = 10'd151; a_exp3 = 10'd6;
b_exp0 = 10'd587; b_exp1 = 10'd709; b_exp2 = 10'd778; b_exp3 = 10'd595;
a_sign0 = 4'd13; a_sign1 = 4'd8; a_sign2 = 4'd0; a_sign3 = 4'd1;
b_sign0 = 4'd3; b_sign1 = 4'd9; b_sign2 = 4'd0; b_sign3 = 4'd4;
@(posedge clk_i);
a_mant0 = 8'd54; a_mant1 = 8'd167; a_mant2 = 8'd2; a_mant3 = 8'd188;
b_mant0 = 8'd69; b_mant1 = 8'd175; b_mant2 = 8'd179; b_mant3 = 8'd98;
a_exp0 = 10'd24; a_exp1 = 10'd949; a_exp2 = 10'd620; a_exp3 = 10'd876;
b_exp0 = 10'd793; b_exp1 = 10'd1019; b_exp2 = 10'd188; b_exp3 = 10'd567;
a_sign0 = 4'd7; a_sign1 = 4'd14; a_sign2 = 4'd15; a_sign3 = 4'd0;
b_sign0 = 4'd13; b_sign1 = 4'd13; b_sign2 = 4'd13; b_sign3 = 4'd4;
@(posedge clk_i);
a_mant0 = 8'd97; a_mant1 = 8'd248; a_mant2 = 8'd80; a_mant3 = 8'd107;
b_mant0 = 8'd145; b_mant1 = 8'd187; b_mant2 = 8'd212; b_mant3 = 8'd200;
a_exp0 = 10'd775; a_exp1 = 10'd602; a_exp2 = 10'd664; a_exp3 = 10'd527;
b_exp0 = 10'd722; b_exp1 = 10'd25; b_exp2 = 10'd495; b_exp3 = 10'd921;
a_sign0 = 4'd2; a_sign1 = 4'd10; a_sign2 = 4'd9; a_sign3 = 4'd9;
b_sign0 = 4'd14; b_sign1 = 4'd12; b_sign2 = 4'd6; b_sign3 = 4'd11;
@(posedge clk_i);
a_mant0 = 8'd113; a_mant1 = 8'd219; a_mant2 = 8'd174; a_mant3 = 8'd17;
b_mant0 = 8'd10; b_mant1 = 8'd183; b_mant2 = 8'd134; b_mant3 = 8'd184;
a_exp0 = 10'd143; a_exp1 = 10'd333; a_exp2 = 10'd551; a_exp3 = 10'd214;
b_exp0 = 10'd800; b_exp1 = 10'd833; b_exp2 = 10'd170; b_exp3 = 10'd332;
a_sign0 = 4'd1; a_sign1 = 4'd10; a_sign2 = 4'd10; a_sign3 = 4'd13;
b_sign0 = 4'd2; b_sign1 = 4'd15; b_sign2 = 4'd5; b_sign3 = 4'd11;
@(posedge clk_i);
a_mant0 = 8'd0; a_mant1 = 8'd227; a_mant2 = 8'd209; a_mant3 = 8'd29;
b_mant0 = 8'd163; b_mant1 = 8'd218; b_mant2 = 8'd38; b_mant3 = 8'd238;
a_exp0 = 10'd423; a_exp1 = 10'd63; a_exp2 = 10'd210; a_exp3 = 10'd253;
b_exp0 = 10'd767; b_exp1 = 10'd346; b_exp2 = 10'd336; b_exp3 = 10'd536;
a_sign0 = 4'd16; a_sign1 = 4'd10; a_sign2 = 4'd8; a_sign3 = 4'd12;
b_sign0 = 4'd8; b_sign1 = 4'd9; b_sign2 = 4'd16; b_sign3 = 4'd12;
@(posedge clk_i);
shared_exps0 = 8'd173;
shared_exps1 = 8'd122;
a_mant0 = 8'd135; a_mant1 = 8'd77; a_mant2 = 8'd32; a_mant3 = 8'd200;
b_mant0 = 8'd68; b_mant1 = 8'd180; b_mant2 = 8'd139; b_mant3 = 8'd120;
a_exp0 = 10'd373; a_exp1 = 10'd137; a_exp2 = 10'd85; a_exp3 = 10'd697;
b_exp0 = 10'd358; b_exp1 = 10'd618; b_exp2 = 10'd495; b_exp3 = 10'd348;
a_sign0 = 4'd9; a_sign1 = 4'd7; a_sign2 = 4'd16; a_sign3 = 4'd12;
b_sign0 = 4'd15; b_sign1 = 4'd15; b_sign2 = 4'd0; b_sign3 = 4'd6;
@(posedge clk_i);
a_mant0 = 8'd204; a_mant1 = 8'd10; a_mant2 = 8'd197; a_mant3 = 8'd10;
b_mant0 = 8'd243; b_mant1 = 8'd76; b_mant2 = 8'd37; b_mant3 = 8'd42;
a_exp0 = 10'd199; a_exp1 = 10'd20; a_exp2 = 10'd735; a_exp3 = 10'd673;
b_exp0 = 10'd697; b_exp1 = 10'd551; b_exp2 = 10'd752; b_exp3 = 10'd597;
a_sign0 = 4'd1; a_sign1 = 4'd13; a_sign2 = 4'd6; a_sign3 = 4'd2;
b_sign0 = 4'd6; b_sign1 = 4'd14; b_sign2 = 4'd13; b_sign3 = 4'd7;
@(posedge clk_i);
a_mant0 = 8'd10; a_mant1 = 8'd27; a_mant2 = 8'd241; a_mant3 = 8'd180;
b_mant0 = 8'd61; b_mant1 = 8'd127; b_mant2 = 8'd225; b_mant3 = 8'd93;
a_exp0 = 10'd502; a_exp1 = 10'd102; a_exp2 = 10'd1005; a_exp3 = 10'd729;
b_exp0 = 10'd245; b_exp1 = 10'd502; b_exp2 = 10'd610; b_exp3 = 10'd704;
a_sign0 = 4'd7; a_sign1 = 4'd9; a_sign2 = 4'd14; a_sign3 = 4'd14;
b_sign0 = 4'd7; b_sign1 = 4'd8; b_sign2 = 4'd16; b_sign3 = 4'd13;
@(posedge clk_i);
a_mant0 = 8'd226; a_mant1 = 8'd137; a_mant2 = 8'd119; a_mant3 = 8'd64;
b_mant0 = 8'd159; b_mant1 = 8'd141; b_mant2 = 8'd34; b_mant3 = 8'd250;
a_exp0 = 10'd63; a_exp1 = 10'd689; a_exp2 = 10'd138; a_exp3 = 10'd967;
b_exp0 = 10'd471; b_exp1 = 10'd397; b_exp2 = 10'd976; b_exp3 = 10'd599;
a_sign0 = 4'd2; a_sign1 = 4'd9; a_sign2 = 4'd16; a_sign3 = 4'd16;
b_sign0 = 4'd6; b_sign1 = 4'd12; b_sign2 = 4'd7; b_sign3 = 4'd9;
@(posedge clk_i);
a_mant0 = 8'd163; a_mant1 = 8'd5; a_mant2 = 8'd13; a_mant3 = 8'd50;
b_mant0 = 8'd145; b_mant1 = 8'd192; b_mant2 = 8'd10; b_mant3 = 8'd31;
a_exp0 = 10'd663; a_exp1 = 10'd503; a_exp2 = 10'd845; a_exp3 = 10'd554;
b_exp0 = 10'd703; b_exp1 = 10'd194; b_exp2 = 10'd30; b_exp3 = 10'd443;
a_sign0 = 4'd1; a_sign1 = 4'd0; a_sign2 = 4'd1; a_sign3 = 4'd1;
b_sign0 = 4'd14; b_sign1 = 4'd3; b_sign2 = 4'd1; b_sign3 = 4'd5;
@(posedge clk_i);
a_mant0 = 8'd182; a_mant1 = 8'd237; a_mant2 = 8'd236; a_mant3 = 8'd48;
b_mant0 = 8'd105; b_mant1 = 8'd167; b_mant2 = 8'd229; b_mant3 = 8'd51;
a_exp0 = 10'd837; a_exp1 = 10'd298; a_exp2 = 10'd343; a_exp3 = 10'd600;
b_exp0 = 10'd129; b_exp1 = 10'd958; b_exp2 = 10'd502; b_exp3 = 10'd154;
a_sign0 = 4'd0; a_sign1 = 4'd13; a_sign2 = 4'd13; a_sign3 = 4'd10;
b_sign0 = 4'd4; b_sign1 = 4'd13; b_sign2 = 4'd13; b_sign3 = 4'd11;
@(posedge clk_i);
a_mant0 = 8'd130; a_mant1 = 8'd95; a_mant2 = 8'd12; a_mant3 = 8'd164;
b_mant0 = 8'd64; b_mant1 = 8'd78; b_mant2 = 8'd106; b_mant3 = 8'd182;
a_exp0 = 10'd196; a_exp1 = 10'd262; a_exp2 = 10'd132; a_exp3 = 10'd412;
b_exp0 = 10'd1002; b_exp1 = 10'd527; b_exp2 = 10'd360; b_exp3 = 10'd222;
a_sign0 = 4'd11; a_sign1 = 4'd9; a_sign2 = 4'd5; a_sign3 = 4'd16;
b_sign0 = 4'd2; b_sign1 = 4'd4; b_sign2 = 4'd16; b_sign3 = 4'd4;
@(posedge clk_i);
a_mant0 = 8'd101; a_mant1 = 8'd59; a_mant2 = 8'd245; a_mant3 = 8'd143;
b_mant0 = 8'd246; b_mant1 = 8'd136; b_mant2 = 8'd162; b_mant3 = 8'd115;
a_exp0 = 10'd67; a_exp1 = 10'd967; a_exp2 = 10'd190; a_exp3 = 10'd725;
b_exp0 = 10'd879; b_exp1 = 10'd138; b_exp2 = 10'd619; b_exp3 = 10'd120;
a_sign0 = 4'd6; a_sign1 = 4'd1; a_sign2 = 4'd4; a_sign3 = 4'd0;
b_sign0 = 4'd6; b_sign1 = 4'd12; b_sign2 = 4'd11; b_sign3 = 4'd5;
@(posedge clk_i);
shared_exps0 = 8'd125;
shared_exps1 = 8'd119;
rstn = 0;
@(posedge clk_i);
rstn = 1;
a_mant0 = 8'd75; a_mant1 = 8'd206; a_mant2 = 8'd237; a_mant3 = 8'd193;
b_mant0 = 8'd181; b_mant1 = 8'd28; b_mant2 = 8'd204; b_mant3 = 8'd191;
a_exp0 = 10'd263; a_exp1 = 10'd46; a_exp2 = 10'd780; a_exp3 = 10'd21;
b_exp0 = 10'd771; b_exp1 = 10'd259; b_exp2 = 10'd724; b_exp3 = 10'd991;
a_sign0 = 4'd12; a_sign1 = 4'd16; a_sign2 = 4'd7; a_sign3 = 4'd4;
b_sign0 = 4'd9; b_sign1 = 4'd1; b_sign2 = 4'd6; b_sign3 = 4'd11;
@(posedge clk_i);
a_mant0 = 8'd155; a_mant1 = 8'd22; a_mant2 = 8'd255; a_mant3 = 8'd120;
b_mant0 = 8'd72; b_mant1 = 8'd241; b_mant2 = 8'd233; b_mant3 = 8'd52;
a_exp0 = 10'd399; a_exp1 = 10'd480; a_exp2 = 10'd831; a_exp3 = 10'd297;
b_exp0 = 10'd277; b_exp1 = 10'd103; b_exp2 = 10'd673; b_exp3 = 10'd881;
a_sign0 = 4'd15; a_sign1 = 4'd10; a_sign2 = 4'd14; a_sign3 = 4'd4;
b_sign0 = 4'd11; b_sign1 = 4'd10; b_sign2 = 4'd4; b_sign3 = 4'd14;
@(posedge clk_i);
a_mant0 = 8'd160; a_mant1 = 8'd105; a_mant2 = 8'd175; a_mant3 = 8'd53;
b_mant0 = 8'd211; b_mant1 = 8'd176; b_mant2 = 8'd63; b_mant3 = 8'd89;
a_exp0 = 10'd302; a_exp1 = 10'd225; a_exp2 = 10'd381; a_exp3 = 10'd852;
b_exp0 = 10'd600; b_exp1 = 10'd680; b_exp2 = 10'd865; b_exp3 = 10'd405;
a_sign0 = 4'd14; a_sign1 = 4'd8; a_sign2 = 4'd1; a_sign3 = 4'd15;
b_sign0 = 4'd15; b_sign1 = 4'd7; b_sign2 = 4'd8; b_sign3 = 4'd9;
@(posedge clk_i);
a_mant0 = 8'd213; a_mant1 = 8'd25; a_mant2 = 8'd159; a_mant3 = 8'd219;
b_mant0 = 8'd41; b_mant1 = 8'd162; b_mant2 = 8'd23; b_mant3 = 8'd117;
a_exp0 = 10'd61; a_exp1 = 10'd752; a_exp2 = 10'd462; a_exp3 = 10'd242;
b_exp0 = 10'd137; b_exp1 = 10'd693; b_exp2 = 10'd848; b_exp3 = 10'd509;
a_sign0 = 4'd0; a_sign1 = 4'd14; a_sign2 = 4'd6; a_sign3 = 4'd12;
b_sign0 = 4'd13; b_sign1 = 4'd9; b_sign2 = 4'd6; b_sign3 = 4'd1;
@(posedge clk_i);
a_mant0 = 8'd254; a_mant1 = 8'd3; a_mant2 = 8'd82; a_mant3 = 8'd108;
b_mant0 = 8'd222; b_mant1 = 8'd136; b_mant2 = 8'd142; b_mant3 = 8'd168;
a_exp0 = 10'd236; a_exp1 = 10'd607; a_exp2 = 10'd849; a_exp3 = 10'd36;
b_exp0 = 10'd168; b_exp1 = 10'd319; b_exp2 = 10'd280; b_exp3 = 10'd129;
a_sign0 = 4'd15; a_sign1 = 4'd15; a_sign2 = 4'd4; a_sign3 = 4'd15;
b_sign0 = 4'd15; b_sign1 = 4'd9; b_sign2 = 4'd4; b_sign3 = 4'd9;
@(posedge clk_i);
a_mant0 = 8'd169; a_mant1 = 8'd144; a_mant2 = 8'd224; a_mant3 = 8'd21;
b_mant0 = 8'd15; b_mant1 = 8'd177; b_mant2 = 8'd140; b_mant3 = 8'd244;
a_exp0 = 10'd388; a_exp1 = 10'd555; a_exp2 = 10'd126; a_exp3 = 10'd479;
b_exp0 = 10'd344; b_exp1 = 10'd942; b_exp2 = 10'd486; b_exp3 = 10'd983;
a_sign0 = 4'd5; a_sign1 = 4'd6; a_sign2 = 4'd3; a_sign3 = 4'd11;
b_sign0 = 4'd11; b_sign1 = 4'd13; b_sign2 = 4'd14; b_sign3 = 4'd3;
@(posedge clk_i);
a_mant0 = 8'd164; a_mant1 = 8'd184; a_mant2 = 8'd214; a_mant3 = 8'd120;
b_mant0 = 8'd1; b_mant1 = 8'd126; b_mant2 = 8'd116; b_mant3 = 8'd43;
a_exp0 = 10'd701; a_exp1 = 10'd766; a_exp2 = 10'd633; a_exp3 = 10'd359;
b_exp0 = 10'd305; b_exp1 = 10'd419; b_exp2 = 10'd559; b_exp3 = 10'd1018;
a_sign0 = 4'd12; a_sign1 = 4'd7; a_sign2 = 4'd6; a_sign3 = 4'd0;
b_sign0 = 4'd14; b_sign1 = 4'd4; b_sign2 = 4'd5; b_sign3 = 4'd13;
@(posedge clk_i);
shared_exps0 = 8'd127;
shared_exps1 = 8'd133;
a_mant0 = 8'd62; a_mant1 = 8'd51; a_mant2 = 8'd8; a_mant3 = 8'd30;
b_mant0 = 8'd177; b_mant1 = 8'd219; b_mant2 = 8'd112; b_mant3 = 8'd163;
a_exp0 = 10'd773; a_exp1 = 10'd579; a_exp2 = 10'd53; a_exp3 = 10'd658;
b_exp0 = 10'd301; b_exp1 = 10'd221; b_exp2 = 10'd363; b_exp3 = 10'd302;
a_sign0 = 4'd11; a_sign1 = 4'd10; a_sign2 = 4'd3; a_sign3 = 4'd15;
b_sign0 = 4'd10; b_sign1 = 4'd12; b_sign2 = 4'd8; b_sign3 = 4'd6;
@(posedge clk_i);
a_mant0 = 8'd18; a_mant1 = 8'd137; a_mant2 = 8'd122; a_mant3 = 8'd212;
b_mant0 = 8'd200; b_mant1 = 8'd163; b_mant2 = 8'd20; b_mant3 = 8'd199;
a_exp0 = 10'd155; a_exp1 = 10'd690; a_exp2 = 10'd284; a_exp3 = 10'd95;
b_exp0 = 10'd977; b_exp1 = 10'd532; b_exp2 = 10'd976; b_exp3 = 10'd928;
a_sign0 = 4'd2; a_sign1 = 4'd14; a_sign2 = 4'd0; a_sign3 = 4'd3;
b_sign0 = 4'd9; b_sign1 = 4'd13; b_sign2 = 4'd13; b_sign3 = 4'd0;
@(posedge clk_i);
a_mant0 = 8'd39; a_mant1 = 8'd37; a_mant2 = 8'd159; a_mant3 = 8'd63;
b_mant0 = 8'd138; b_mant1 = 8'd216; b_mant2 = 8'd220; b_mant3 = 8'd254;
a_exp0 = 10'd592; a_exp1 = 10'd33; a_exp2 = 10'd152; a_exp3 = 10'd1003;
b_exp0 = 10'd78; b_exp1 = 10'd206; b_exp2 = 10'd165; b_exp3 = 10'd892;
a_sign0 = 4'd1; a_sign1 = 4'd4; a_sign2 = 4'd10; a_sign3 = 4'd12;
b_sign0 = 4'd10; b_sign1 = 4'd0; b_sign2 = 4'd2; b_sign3 = 4'd9;
@(posedge clk_i);
a_mant0 = 8'd30; a_mant1 = 8'd171; a_mant2 = 8'd243; a_mant3 = 8'd218;
b_mant0 = 8'd118; b_mant1 = 8'd234; b_mant2 = 8'd155; b_mant3 = 8'd9;
a_exp0 = 10'd108; a_exp1 = 10'd217; a_exp2 = 10'd404; a_exp3 = 10'd22;
b_exp0 = 10'd358; b_exp1 = 10'd512; b_exp2 = 10'd116; b_exp3 = 10'd89;
a_sign0 = 4'd11; a_sign1 = 4'd14; a_sign2 = 4'd6; a_sign3 = 4'd9;
b_sign0 = 4'd13; b_sign1 = 4'd8; b_sign2 = 4'd14; b_sign3 = 4'd9;
@(posedge clk_i);
a_mant0 = 8'd113; a_mant1 = 8'd164; a_mant2 = 8'd21; a_mant3 = 8'd243;
b_mant0 = 8'd244; b_mant1 = 8'd77; b_mant2 = 8'd46; b_mant3 = 8'd39;
a_exp0 = 10'd845; a_exp1 = 10'd506; a_exp2 = 10'd543; a_exp3 = 10'd510;
b_exp0 = 10'd496; b_exp1 = 10'd466; b_exp2 = 10'd268; b_exp3 = 10'd988;
a_sign0 = 4'd8; a_sign1 = 4'd10; a_sign2 = 4'd16; a_sign3 = 4'd14;
b_sign0 = 4'd16; b_sign1 = 4'd0; b_sign2 = 4'd9; b_sign3 = 4'd8;
@(posedge clk_i);
a_mant0 = 8'd127; a_mant1 = 8'd76; a_mant2 = 8'd148; a_mant3 = 8'd244;
b_mant0 = 8'd2; b_mant1 = 8'd202; b_mant2 = 8'd155; b_mant3 = 8'd38;
a_exp0 = 10'd17; a_exp1 = 10'd765; a_exp2 = 10'd940; a_exp3 = 10'd895;
b_exp0 = 10'd790; b_exp1 = 10'd906; b_exp2 = 10'd890; b_exp3 = 10'd43;
a_sign0 = 4'd8; a_sign1 = 4'd1; a_sign2 = 4'd6; a_sign3 = 4'd15;
b_sign0 = 4'd9; b_sign1 = 4'd4; b_sign2 = 4'd4; b_sign3 = 4'd16;
@(posedge clk_i);
a_mant0 = 8'd15; a_mant1 = 8'd253; a_mant2 = 8'd246; a_mant3 = 8'd40;
b_mant0 = 8'd139; b_mant1 = 8'd191; b_mant2 = 8'd209; b_mant3 = 8'd235;
a_exp0 = 10'd408; a_exp1 = 10'd548; a_exp2 = 10'd379; a_exp3 = 10'd266;
b_exp0 = 10'd275; b_exp1 = 10'd129; b_exp2 = 10'd987; b_exp3 = 10'd597;
a_sign0 = 4'd4; a_sign1 = 4'd9; a_sign2 = 4'd11; a_sign3 = 4'd0;
b_sign0 = 4'd3; b_sign1 = 4'd5; b_sign2 = 4'd4; b_sign3 = 4'd14;
@(posedge clk_i);
a_mant0 = 8'd202; a_mant1 = 8'd184; a_mant2 = 8'd130; a_mant3 = 8'd216;
b_mant0 = 8'd3; b_mant1 = 8'd173; b_mant2 = 8'd253; b_mant3 = 8'd198;
a_exp0 = 10'd871; a_exp1 = 10'd217; a_exp2 = 10'd223; a_exp3 = 10'd327;
b_exp0 = 10'd40; b_exp1 = 10'd731; b_exp2 = 10'd595; b_exp3 = 10'd320;
a_sign0 = 4'd3; a_sign1 = 4'd14; a_sign2 = 4'd0; a_sign3 = 4'd1;
b_sign0 = 4'd9; b_sign1 = 4'd1; b_sign2 = 4'd10; b_sign3 = 4'd11;
@(posedge clk_i);
shared_exps0 = 8'd127;
shared_exps1 = 8'd122;
a_mant0 = 8'd219; a_mant1 = 8'd10; a_mant2 = 8'd200; a_mant3 = 8'd21;
b_mant0 = 8'd117; b_mant1 = 8'd169; b_mant2 = 8'd183; b_mant3 = 8'd83;
a_exp0 = 10'd437; a_exp1 = 10'd785; a_exp2 = 10'd217; a_exp3 = 10'd490;
b_exp0 = 10'd197; b_exp1 = 10'd840; b_exp2 = 10'd917; b_exp3 = 10'd297;
a_sign0 = 4'd16; a_sign1 = 4'd11; a_sign2 = 4'd12; a_sign3 = 4'd1;
b_sign0 = 4'd0; b_sign1 = 4'd16; b_sign2 = 4'd2; b_sign3 = 4'd0;
@(posedge clk_i);
a_mant0 = 8'd43; a_mant1 = 8'd126; a_mant2 = 8'd215; a_mant3 = 8'd4;
b_mant0 = 8'd174; b_mant1 = 8'd129; b_mant2 = 8'd162; b_mant3 = 8'd36;
a_exp0 = 10'd487; a_exp1 = 10'd690; a_exp2 = 10'd342; a_exp3 = 10'd172;
b_exp0 = 10'd788; b_exp1 = 10'd801; b_exp2 = 10'd433; b_exp3 = 10'd42;
a_sign0 = 4'd4; a_sign1 = 4'd3; a_sign2 = 4'd6; a_sign3 = 4'd10;
b_sign0 = 4'd10; b_sign1 = 4'd0; b_sign2 = 4'd7; b_sign3 = 4'd0;
@(posedge clk_i);
a_mant0 = 8'd219; a_mant1 = 8'd6; a_mant2 = 8'd236; a_mant3 = 8'd154;
b_mant0 = 8'd76; b_mant1 = 8'd93; b_mant2 = 8'd238; b_mant3 = 8'd230;
a_exp0 = 10'd226; a_exp1 = 10'd1002; a_exp2 = 10'd173; a_exp3 = 10'd966;
b_exp0 = 10'd567; b_exp1 = 10'd917; b_exp2 = 10'd680; b_exp3 = 10'd546;
a_sign0 = 4'd4; a_sign1 = 4'd5; a_sign2 = 4'd10; a_sign3 = 4'd3;
b_sign0 = 4'd13; b_sign1 = 4'd10; b_sign2 = 4'd10; b_sign3 = 4'd10;
@(posedge clk_i);
a_mant0 = 8'd223; a_mant1 = 8'd217; a_mant2 = 8'd1; a_mant3 = 8'd106;
b_mant0 = 8'd197; b_mant1 = 8'd254; b_mant2 = 8'd230; b_mant3 = 8'd112;
a_exp0 = 10'd912; a_exp1 = 10'd338; a_exp2 = 10'd654; a_exp3 = 10'd289;
b_exp0 = 10'd445; b_exp1 = 10'd750; b_exp2 = 10'd258; b_exp3 = 10'd553;
a_sign0 = 4'd15; a_sign1 = 4'd13; a_sign2 = 4'd8; a_sign3 = 4'd3;
b_sign0 = 4'd4; b_sign1 = 4'd16; b_sign2 = 4'd12; b_sign3 = 4'd10;
@(posedge clk_i);
a_mant0 = 8'd25; a_mant1 = 8'd2; a_mant2 = 8'd223; a_mant3 = 8'd153;
b_mant0 = 8'd105; b_mant1 = 8'd45; b_mant2 = 8'd163; b_mant3 = 8'd11;
a_exp0 = 10'd320; a_exp1 = 10'd905; a_exp2 = 10'd490; a_exp3 = 10'd833;
b_exp0 = 10'd642; b_exp1 = 10'd334; b_exp2 = 10'd878; b_exp3 = 10'd79;
a_sign0 = 4'd5; a_sign1 = 4'd3; a_sign2 = 4'd10; a_sign3 = 4'd1;
b_sign0 = 4'd3; b_sign1 = 4'd14; b_sign2 = 4'd0; b_sign3 = 4'd5;
@(posedge clk_i);
a_mant0 = 8'd60; a_mant1 = 8'd54; a_mant2 = 8'd101; a_mant3 = 8'd198;
b_mant0 = 8'd99; b_mant1 = 8'd101; b_mant2 = 8'd169; b_mant3 = 8'd22;
a_exp0 = 10'd665; a_exp1 = 10'd40; a_exp2 = 10'd590; a_exp3 = 10'd807;
b_exp0 = 10'd263; b_exp1 = 10'd668; b_exp2 = 10'd40; b_exp3 = 10'd956;
a_sign0 = 4'd10; a_sign1 = 4'd7; a_sign2 = 4'd10; a_sign3 = 4'd15;
b_sign0 = 4'd11; b_sign1 = 4'd1; b_sign2 = 4'd2; b_sign3 = 4'd3;
@(posedge clk_i);
a_mant0 = 8'd160; a_mant1 = 8'd159; a_mant2 = 8'd129; a_mant3 = 8'd244;
b_mant0 = 8'd158; b_mant1 = 8'd151; b_mant2 = 8'd247; b_mant3 = 8'd103;
a_exp0 = 10'd59; a_exp1 = 10'd157; a_exp2 = 10'd218; a_exp3 = 10'd767;
b_exp0 = 10'd538; b_exp1 = 10'd379; b_exp2 = 10'd625; b_exp3 = 10'd441;
a_sign0 = 4'd2; a_sign1 = 4'd7; a_sign2 = 4'd1; a_sign3 = 4'd7;
b_sign0 = 4'd0; b_sign1 = 4'd14; b_sign2 = 4'd2; b_sign3 = 4'd14;
@(posedge clk_i);
a_mant0 = 8'd72; a_mant1 = 8'd71; a_mant2 = 8'd173; a_mant3 = 8'd176;
b_mant0 = 8'd96; b_mant1 = 8'd6; b_mant2 = 8'd70; b_mant3 = 8'd183;
a_exp0 = 10'd327; a_exp1 = 10'd621; a_exp2 = 10'd614; a_exp3 = 10'd867;
b_exp0 = 10'd747; b_exp1 = 10'd533; b_exp2 = 10'd611; b_exp3 = 10'd272;
a_sign0 = 4'd13; a_sign1 = 4'd1; a_sign2 = 4'd13; a_sign3 = 4'd16;
b_sign0 = 4'd7; b_sign1 = 4'd1; b_sign2 = 4'd8; b_sign3 = 4'd6;
@(posedge clk_i);
shared_exps0 = 8'd161;
shared_exps1 = 8'd134;
a_mant0 = 8'd232; a_mant1 = 8'd68; a_mant2 = 8'd103; a_mant3 = 8'd78;
b_mant0 = 8'd252; b_mant1 = 8'd86; b_mant2 = 8'd13; b_mant3 = 8'd27;
a_exp0 = 10'd354; a_exp1 = 10'd810; a_exp2 = 10'd560; a_exp3 = 10'd922;
b_exp0 = 10'd655; b_exp1 = 10'd655; b_exp2 = 10'd716; b_exp3 = 10'd190;
a_sign0 = 4'd3; a_sign1 = 4'd16; a_sign2 = 4'd14; a_sign3 = 4'd12;
b_sign0 = 4'd7; b_sign1 = 4'd7; b_sign2 = 4'd6; b_sign3 = 4'd14;
@(posedge clk_i);
a_mant0 = 8'd187; a_mant1 = 8'd53; a_mant2 = 8'd56; a_mant3 = 8'd66;
b_mant0 = 8'd198; b_mant1 = 8'd253; b_mant2 = 8'd209; b_mant3 = 8'd35;
a_exp0 = 10'd371; a_exp1 = 10'd702; a_exp2 = 10'd327; a_exp3 = 10'd150;
b_exp0 = 10'd953; b_exp1 = 10'd53; b_exp2 = 10'd22; b_exp3 = 10'd288;
a_sign0 = 4'd0; a_sign1 = 4'd8; a_sign2 = 4'd3; a_sign3 = 4'd1;
b_sign0 = 4'd3; b_sign1 = 4'd10; b_sign2 = 4'd7; b_sign3 = 4'd11;
@(posedge clk_i);
a_mant0 = 8'd202; a_mant1 = 8'd94; a_mant2 = 8'd29; a_mant3 = 8'd178;
b_mant0 = 8'd239; b_mant1 = 8'd150; b_mant2 = 8'd200; b_mant3 = 8'd236;
a_exp0 = 10'd348; a_exp1 = 10'd956; a_exp2 = 10'd624; a_exp3 = 10'd935;
b_exp0 = 10'd18; b_exp1 = 10'd812; b_exp2 = 10'd964; b_exp3 = 10'd1005;
a_sign0 = 4'd5; a_sign1 = 4'd3; a_sign2 = 4'd9; a_sign3 = 4'd8;
b_sign0 = 4'd6; b_sign1 = 4'd5; b_sign2 = 4'd12; b_sign3 = 4'd10;
@(posedge clk_i);
a_mant0 = 8'd163; a_mant1 = 8'd54; a_mant2 = 8'd179; a_mant3 = 8'd158;
b_mant0 = 8'd40; b_mant1 = 8'd92; b_mant2 = 8'd234; b_mant3 = 8'd141;
a_exp0 = 10'd903; a_exp1 = 10'd193; a_exp2 = 10'd247; a_exp3 = 10'd984;
b_exp0 = 10'd937; b_exp1 = 10'd193; b_exp2 = 10'd692; b_exp3 = 10'd586;
a_sign0 = 4'd16; a_sign1 = 4'd11; a_sign2 = 4'd6; a_sign3 = 4'd2;
b_sign0 = 4'd1; b_sign1 = 4'd0; b_sign2 = 4'd6; b_sign3 = 4'd5;
@(posedge clk_i);
a_mant0 = 8'd73; a_mant1 = 8'd94; a_mant2 = 8'd126; a_mant3 = 8'd53;
b_mant0 = 8'd203; b_mant1 = 8'd206; b_mant2 = 8'd103; b_mant3 = 8'd249;
a_exp0 = 10'd404; a_exp1 = 10'd8; a_exp2 = 10'd255; a_exp3 = 10'd169;
b_exp0 = 10'd963; b_exp1 = 10'd776; b_exp2 = 10'd874; b_exp3 = 10'd343;
a_sign0 = 4'd9; a_sign1 = 4'd2; a_sign2 = 4'd13; a_sign3 = 4'd14;
b_sign0 = 4'd15; b_sign1 = 4'd4; b_sign2 = 4'd13; b_sign3 = 4'd0;
@(posedge clk_i);
a_mant0 = 8'd12; a_mant1 = 8'd177; a_mant2 = 8'd154; a_mant3 = 8'd16;
b_mant0 = 8'd153; b_mant1 = 8'd73; b_mant2 = 8'd207; b_mant3 = 8'd43;
a_exp0 = 10'd484; a_exp1 = 10'd841; a_exp2 = 10'd994; a_exp3 = 10'd385;
b_exp0 = 10'd857; b_exp1 = 10'd713; b_exp2 = 10'd933; b_exp3 = 10'd274;
a_sign0 = 4'd10; a_sign1 = 4'd15; a_sign2 = 4'd3; a_sign3 = 4'd7;
b_sign0 = 4'd12; b_sign1 = 4'd13; b_sign2 = 4'd6; b_sign3 = 4'd16;
@(posedge clk_i);
a_mant0 = 8'd178; a_mant1 = 8'd167; a_mant2 = 8'd198; a_mant3 = 8'd143;
b_mant0 = 8'd67; b_mant1 = 8'd46; b_mant2 = 8'd118; b_mant3 = 8'd36;
a_exp0 = 10'd851; a_exp1 = 10'd425; a_exp2 = 10'd737; a_exp3 = 10'd409;
b_exp0 = 10'd944; b_exp1 = 10'd130; b_exp2 = 10'd86; b_exp3 = 10'd750;
a_sign0 = 4'd10; a_sign1 = 4'd14; a_sign2 = 4'd15; a_sign3 = 4'd4;
b_sign0 = 4'd9; b_sign1 = 4'd14; b_sign2 = 4'd14; b_sign3 = 4'd8;
@(posedge clk_i);
a_mant0 = 8'd170; a_mant1 = 8'd41; a_mant2 = 8'd68; a_mant3 = 8'd9;
b_mant0 = 8'd221; b_mant1 = 8'd140; b_mant2 = 8'd36; b_mant3 = 8'd86;
a_exp0 = 10'd957; a_exp1 = 10'd228; a_exp2 = 10'd717; a_exp3 = 10'd255;
b_exp0 = 10'd48; b_exp1 = 10'd721; b_exp2 = 10'd962; b_exp3 = 10'd97;
a_sign0 = 4'd12; a_sign1 = 4'd10; a_sign2 = 4'd12; a_sign3 = 4'd7;
b_sign0 = 4'd10; b_sign1 = 4'd9; b_sign2 = 4'd7; b_sign3 = 4'd8;
@(posedge clk_i);
shared_exps0 = 8'd136;
shared_exps1 = 8'd118;
rstn = 0;
@(posedge clk_i);
rstn = 1;
a_mant0 = 8'd180; a_mant1 = 8'd218; a_mant2 = 8'd4; a_mant3 = 8'd95;
b_mant0 = 8'd37; b_mant1 = 8'd143; b_mant2 = 8'd4; b_mant3 = 8'd195;
a_exp0 = 10'd235; a_exp1 = 10'd304; a_exp2 = 10'd655; a_exp3 = 10'd754;
b_exp0 = 10'd925; b_exp1 = 10'd693; b_exp2 = 10'd806; b_exp3 = 10'd43;
a_sign0 = 4'd2; a_sign1 = 4'd2; a_sign2 = 4'd12; a_sign3 = 4'd0;
b_sign0 = 4'd4; b_sign1 = 4'd7; b_sign2 = 4'd13; b_sign3 = 4'd9;
@(posedge clk_i);
a_mant0 = 8'd114; a_mant1 = 8'd92; a_mant2 = 8'd107; a_mant3 = 8'd160;
b_mant0 = 8'd189; b_mant1 = 8'd6; b_mant2 = 8'd4; b_mant3 = 8'd99;
a_exp0 = 10'd220; a_exp1 = 10'd598; a_exp2 = 10'd518; a_exp3 = 10'd682;
b_exp0 = 10'd379; b_exp1 = 10'd264; b_exp2 = 10'd187; b_exp3 = 10'd185;
a_sign0 = 4'd5; a_sign1 = 4'd13; a_sign2 = 4'd9; a_sign3 = 4'd5;
b_sign0 = 4'd8; b_sign1 = 4'd7; b_sign2 = 4'd5; b_sign3 = 4'd0;
@(posedge clk_i);
a_mant0 = 8'd146; a_mant1 = 8'd28; a_mant2 = 8'd14; a_mant3 = 8'd63;
b_mant0 = 8'd36; b_mant1 = 8'd194; b_mant2 = 8'd199; b_mant3 = 8'd229;
a_exp0 = 10'd649; a_exp1 = 10'd240; a_exp2 = 10'd228; a_exp3 = 10'd889;
b_exp0 = 10'd436; b_exp1 = 10'd327; b_exp2 = 10'd672; b_exp3 = 10'd645;
a_sign0 = 4'd5; a_sign1 = 4'd1; a_sign2 = 4'd12; a_sign3 = 4'd3;
b_sign0 = 4'd0; b_sign1 = 4'd2; b_sign2 = 4'd6; b_sign3 = 4'd4;
@(posedge clk_i);
a_mant0 = 8'd73; a_mant1 = 8'd115; a_mant2 = 8'd106; a_mant3 = 8'd238;
b_mant0 = 8'd239; b_mant1 = 8'd16; b_mant2 = 8'd113; b_mant3 = 8'd193;
a_exp0 = 10'd967; a_exp1 = 10'd95; a_exp2 = 10'd505; a_exp3 = 10'd814;
b_exp0 = 10'd592; b_exp1 = 10'd423; b_exp2 = 10'd96; b_exp3 = 10'd818;
a_sign0 = 4'd15; a_sign1 = 4'd8; a_sign2 = 4'd14; a_sign3 = 4'd5;
b_sign0 = 4'd0; b_sign1 = 4'd10; b_sign2 = 4'd2; b_sign3 = 4'd14;
@(posedge clk_i);
a_mant0 = 8'd153; a_mant1 = 8'd200; a_mant2 = 8'd84; a_mant3 = 8'd113;
b_mant0 = 8'd177; b_mant1 = 8'd172; b_mant2 = 8'd142; b_mant3 = 8'd79;
a_exp0 = 10'd70; a_exp1 = 10'd853; a_exp2 = 10'd1014; a_exp3 = 10'd835;
b_exp0 = 10'd820; b_exp1 = 10'd917; b_exp2 = 10'd331; b_exp3 = 10'd949;
a_sign0 = 4'd11; a_sign1 = 4'd16; a_sign2 = 4'd9; a_sign3 = 4'd3;
b_sign0 = 4'd15; b_sign1 = 4'd2; b_sign2 = 4'd16; b_sign3 = 4'd5;
@(posedge clk_i);
a_mant0 = 8'd174; a_mant1 = 8'd209; a_mant2 = 8'd157; a_mant3 = 8'd163;
b_mant0 = 8'd31; b_mant1 = 8'd200; b_mant2 = 8'd35; b_mant3 = 8'd33;
a_exp0 = 10'd996; a_exp1 = 10'd609; a_exp2 = 10'd446; a_exp3 = 10'd24;
b_exp0 = 10'd142; b_exp1 = 10'd667; b_exp2 = 10'd398; b_exp3 = 10'd685;
a_sign0 = 4'd11; a_sign1 = 4'd12; a_sign2 = 4'd2; a_sign3 = 4'd14;
b_sign0 = 4'd10; b_sign1 = 4'd1; b_sign2 = 4'd15; b_sign3 = 4'd15;
@(posedge clk_i);
a_mant0 = 8'd91; a_mant1 = 8'd211; a_mant2 = 8'd9; a_mant3 = 8'd227;
b_mant0 = 8'd221; b_mant1 = 8'd53; b_mant2 = 8'd184; b_mant3 = 8'd180;
a_exp0 = 10'd407; a_exp1 = 10'd882; a_exp2 = 10'd73; a_exp3 = 10'd659;
b_exp0 = 10'd332; b_exp1 = 10'd678; b_exp2 = 10'd456; b_exp3 = 10'd162;
a_sign0 = 4'd15; a_sign1 = 4'd1; a_sign2 = 4'd6; a_sign3 = 4'd12;
b_sign0 = 4'd12; b_sign1 = 4'd6; b_sign2 = 4'd10; b_sign3 = 4'd13;
@(posedge clk_i);
shared_exps0 = 8'd129;
shared_exps1 = 8'd113;
a_mant0 = 8'd28; a_mant1 = 8'd200; a_mant2 = 8'd164; a_mant3 = 8'd251;
b_mant0 = 8'd230; b_mant1 = 8'd41; b_mant2 = 8'd66; b_mant3 = 8'd15;
a_exp0 = 10'd32; a_exp1 = 10'd220; a_exp2 = 10'd429; a_exp3 = 10'd991;
b_exp0 = 10'd295; b_exp1 = 10'd724; b_exp2 = 10'd178; b_exp3 = 10'd828;
a_sign0 = 4'd4; a_sign1 = 4'd8; a_sign2 = 4'd14; a_sign3 = 4'd16;
b_sign0 = 4'd9; b_sign1 = 4'd7; b_sign2 = 4'd7; b_sign3 = 4'd5;
@(posedge clk_i);
a_mant0 = 8'd1; a_mant1 = 8'd193; a_mant2 = 8'd157; a_mant3 = 8'd188;
b_mant0 = 8'd48; b_mant1 = 8'd41; b_mant2 = 8'd45; b_mant3 = 8'd14;
a_exp0 = 10'd687; a_exp1 = 10'd755; a_exp2 = 10'd363; a_exp3 = 10'd889;
b_exp0 = 10'd732; b_exp1 = 10'd945; b_exp2 = 10'd484; b_exp3 = 10'd121;
a_sign0 = 4'd4; a_sign1 = 4'd10; a_sign2 = 4'd4; a_sign3 = 4'd1;
b_sign0 = 4'd13; b_sign1 = 4'd16; b_sign2 = 4'd0; b_sign3 = 4'd11;
@(posedge clk_i);
a_mant0 = 8'd204; a_mant1 = 8'd180; a_mant2 = 8'd251; a_mant3 = 8'd62;
b_mant0 = 8'd227; b_mant1 = 8'd210; b_mant2 = 8'd77; b_mant3 = 8'd70;
a_exp0 = 10'd976; a_exp1 = 10'd514; a_exp2 = 10'd104; a_exp3 = 10'd292;
b_exp0 = 10'd197; b_exp1 = 10'd730; b_exp2 = 10'd957; b_exp3 = 10'd201;
a_sign0 = 4'd13; a_sign1 = 4'd4; a_sign2 = 4'd9; a_sign3 = 4'd7;
b_sign0 = 4'd9; b_sign1 = 4'd14; b_sign2 = 4'd16; b_sign3 = 4'd6;
@(posedge clk_i);
a_mant0 = 8'd213; a_mant1 = 8'd123; a_mant2 = 8'd83; a_mant3 = 8'd239;
b_mant0 = 8'd116; b_mant1 = 8'd109; b_mant2 = 8'd60; b_mant3 = 8'd102;
a_exp0 = 10'd709; a_exp1 = 10'd332; a_exp2 = 10'd761; a_exp3 = 10'd250;
b_exp0 = 10'd951; b_exp1 = 10'd216; b_exp2 = 10'd796; b_exp3 = 10'd488;
a_sign0 = 4'd5; a_sign1 = 4'd0; a_sign2 = 4'd13; a_sign3 = 4'd6;
b_sign0 = 4'd8; b_sign1 = 4'd7; b_sign2 = 4'd7; b_sign3 = 4'd3;
@(posedge clk_i);
a_mant0 = 8'd154; a_mant1 = 8'd0; a_mant2 = 8'd188; a_mant3 = 8'd73;
b_mant0 = 8'd159; b_mant1 = 8'd252; b_mant2 = 8'd115; b_mant3 = 8'd122;
a_exp0 = 10'd940; a_exp1 = 10'd225; a_exp2 = 10'd244; a_exp3 = 10'd6;
b_exp0 = 10'd557; b_exp1 = 10'd434; b_exp2 = 10'd600; b_exp3 = 10'd138;
a_sign0 = 4'd12; a_sign1 = 4'd8; a_sign2 = 4'd13; a_sign3 = 4'd8;
b_sign0 = 4'd11; b_sign1 = 4'd5; b_sign2 = 4'd1; b_sign3 = 4'd13;
@(posedge clk_i);
a_mant0 = 8'd50; a_mant1 = 8'd246; a_mant2 = 8'd63; a_mant3 = 8'd159;
b_mant0 = 8'd3; b_mant1 = 8'd176; b_mant2 = 8'd226; b_mant3 = 8'd246;
a_exp0 = 10'd707; a_exp1 = 10'd507; a_exp2 = 10'd64; a_exp3 = 10'd21;
b_exp0 = 10'd495; b_exp1 = 10'd225; b_exp2 = 10'd47; b_exp3 = 10'd903;
a_sign0 = 4'd9; a_sign1 = 4'd11; a_sign2 = 4'd11; a_sign3 = 4'd10;
b_sign0 = 4'd9; b_sign1 = 4'd10; b_sign2 = 4'd7; b_sign3 = 4'd14;
@(posedge clk_i);
a_mant0 = 8'd188; a_mant1 = 8'd234; a_mant2 = 8'd48; a_mant3 = 8'd178;
b_mant0 = 8'd124; b_mant1 = 8'd248; b_mant2 = 8'd35; b_mant3 = 8'd158;
a_exp0 = 10'd882; a_exp1 = 10'd899; a_exp2 = 10'd393; a_exp3 = 10'd873;
b_exp0 = 10'd458; b_exp1 = 10'd330; b_exp2 = 10'd690; b_exp3 = 10'd258;
a_sign0 = 4'd12; a_sign1 = 4'd10; a_sign2 = 4'd1; a_sign3 = 4'd13;
b_sign0 = 4'd14; b_sign1 = 4'd4; b_sign2 = 4'd9; b_sign3 = 4'd9;
@(posedge clk_i);
a_mant0 = 8'd228; a_mant1 = 8'd14; a_mant2 = 8'd250; a_mant3 = 8'd104;
b_mant0 = 8'd209; b_mant1 = 8'd2; b_mant2 = 8'd75; b_mant3 = 8'd170;
a_exp0 = 10'd107; a_exp1 = 10'd585; a_exp2 = 10'd993; a_exp3 = 10'd213;
b_exp0 = 10'd233; b_exp1 = 10'd861; b_exp2 = 10'd732; b_exp3 = 10'd196;
a_sign0 = 4'd3; a_sign1 = 4'd2; a_sign2 = 4'd5; a_sign3 = 4'd8;
b_sign0 = 4'd6; b_sign1 = 4'd10; b_sign2 = 4'd16; b_sign3 = 4'd7;
@(posedge clk_i);
shared_exps0 = 8'd123;
shared_exps1 = 8'd125;
a_mant0 = 8'd99; a_mant1 = 8'd1; a_mant2 = 8'd229; a_mant3 = 8'd135;
b_mant0 = 8'd108; b_mant1 = 8'd80; b_mant2 = 8'd60; b_mant3 = 8'd3;
a_exp0 = 10'd962; a_exp1 = 10'd327; a_exp2 = 10'd38; a_exp3 = 10'd768;
b_exp0 = 10'd689; b_exp1 = 10'd154; b_exp2 = 10'd995; b_exp3 = 10'd505;
a_sign0 = 4'd16; a_sign1 = 4'd6; a_sign2 = 4'd0; a_sign3 = 4'd14;
b_sign0 = 4'd9; b_sign1 = 4'd8; b_sign2 = 4'd0; b_sign3 = 4'd4;
@(posedge clk_i);
a_mant0 = 8'd56; a_mant1 = 8'd118; a_mant2 = 8'd208; a_mant3 = 8'd99;
b_mant0 = 8'd243; b_mant1 = 8'd33; b_mant2 = 8'd146; b_mant3 = 8'd18;
a_exp0 = 10'd487; a_exp1 = 10'd979; a_exp2 = 10'd793; a_exp3 = 10'd325;
b_exp0 = 10'd927; b_exp1 = 10'd209; b_exp2 = 10'd52; b_exp3 = 10'd179;
a_sign0 = 4'd5; a_sign1 = 4'd10; a_sign2 = 4'd14; a_sign3 = 4'd9;
b_sign0 = 4'd6; b_sign1 = 4'd10; b_sign2 = 4'd15; b_sign3 = 4'd5;
@(posedge clk_i);
a_mant0 = 8'd32; a_mant1 = 8'd149; a_mant2 = 8'd52; a_mant3 = 8'd96;
b_mant0 = 8'd71; b_mant1 = 8'd53; b_mant2 = 8'd25; b_mant3 = 8'd133;
a_exp0 = 10'd269; a_exp1 = 10'd304; a_exp2 = 10'd364; a_exp3 = 10'd830;
b_exp0 = 10'd991; b_exp1 = 10'd725; b_exp2 = 10'd687; b_exp3 = 10'd410;
a_sign0 = 4'd8; a_sign1 = 4'd11; a_sign2 = 4'd1; a_sign3 = 4'd6;
b_sign0 = 4'd4; b_sign1 = 4'd9; b_sign2 = 4'd13; b_sign3 = 4'd12;
@(posedge clk_i);
a_mant0 = 8'd202; a_mant1 = 8'd248; a_mant2 = 8'd23; a_mant3 = 8'd73;
b_mant0 = 8'd146; b_mant1 = 8'd137; b_mant2 = 8'd184; b_mant3 = 8'd137;
a_exp0 = 10'd950; a_exp1 = 10'd819; a_exp2 = 10'd452; a_exp3 = 10'd805;
b_exp0 = 10'd286; b_exp1 = 10'd890; b_exp2 = 10'd15; b_exp3 = 10'd98;
a_sign0 = 4'd1; a_sign1 = 4'd2; a_sign2 = 4'd3; a_sign3 = 4'd8;
b_sign0 = 4'd10; b_sign1 = 4'd8; b_sign2 = 4'd14; b_sign3 = 4'd7;
@(posedge clk_i);
a_mant0 = 8'd44; a_mant1 = 8'd69; a_mant2 = 8'd155; a_mant3 = 8'd226;
b_mant0 = 8'd214; b_mant1 = 8'd21; b_mant2 = 8'd101; b_mant3 = 8'd227;
a_exp0 = 10'd400; a_exp1 = 10'd972; a_exp2 = 10'd314; a_exp3 = 10'd597;
b_exp0 = 10'd452; b_exp1 = 10'd324; b_exp2 = 10'd584; b_exp3 = 10'd102;
a_sign0 = 4'd6; a_sign1 = 4'd3; a_sign2 = 4'd15; a_sign3 = 4'd9;
b_sign0 = 4'd16; b_sign1 = 4'd15; b_sign2 = 4'd10; b_sign3 = 4'd14;
@(posedge clk_i);
a_mant0 = 8'd110; a_mant1 = 8'd40; a_mant2 = 8'd143; a_mant3 = 8'd65;
b_mant0 = 8'd40; b_mant1 = 8'd197; b_mant2 = 8'd41; b_mant3 = 8'd3;
a_exp0 = 10'd123; a_exp1 = 10'd196; a_exp2 = 10'd259; a_exp3 = 10'd178;
b_exp0 = 10'd97; b_exp1 = 10'd395; b_exp2 = 10'd453; b_exp3 = 10'd6;
a_sign0 = 4'd9; a_sign1 = 4'd15; a_sign2 = 4'd12; a_sign3 = 4'd15;
b_sign0 = 4'd12; b_sign1 = 4'd11; b_sign2 = 4'd6; b_sign3 = 4'd11;
@(posedge clk_i);
a_mant0 = 8'd57; a_mant1 = 8'd94; a_mant2 = 8'd90; a_mant3 = 8'd175;
b_mant0 = 8'd77; b_mant1 = 8'd186; b_mant2 = 8'd15; b_mant3 = 8'd187;
a_exp0 = 10'd600; a_exp1 = 10'd888; a_exp2 = 10'd92; a_exp3 = 10'd313;
b_exp0 = 10'd360; b_exp1 = 10'd173; b_exp2 = 10'd865; b_exp3 = 10'd428;
a_sign0 = 4'd1; a_sign1 = 4'd14; a_sign2 = 4'd6; a_sign3 = 4'd16;
b_sign0 = 4'd16; b_sign1 = 4'd15; b_sign2 = 4'd13; b_sign3 = 4'd14;
@(posedge clk_i);
a_mant0 = 8'd216; a_mant1 = 8'd214; a_mant2 = 8'd250; a_mant3 = 8'd196;
b_mant0 = 8'd71; b_mant1 = 8'd249; b_mant2 = 8'd204; b_mant3 = 8'd163;
a_exp0 = 10'd994; a_exp1 = 10'd815; a_exp2 = 10'd145; a_exp3 = 10'd202;
b_exp0 = 10'd880; b_exp1 = 10'd802; b_exp2 = 10'd661; b_exp3 = 10'd524;
a_sign0 = 4'd14; a_sign1 = 4'd0; a_sign2 = 4'd1; a_sign3 = 4'd12;
b_sign0 = 4'd1; b_sign1 = 4'd8; b_sign2 = 4'd6; b_sign3 = 4'd5;
@(posedge clk_i);
shared_exps0 = 8'd117;
shared_exps1 = 8'd147;
a_mant0 = 8'd228; a_mant1 = 8'd119; a_mant2 = 8'd10; a_mant3 = 8'd87;
b_mant0 = 8'd215; b_mant1 = 8'd137; b_mant2 = 8'd186; b_mant3 = 8'd87;
a_exp0 = 10'd726; a_exp1 = 10'd831; a_exp2 = 10'd177; a_exp3 = 10'd324;
b_exp0 = 10'd872; b_exp1 = 10'd645; b_exp2 = 10'd79; b_exp3 = 10'd910;
a_sign0 = 4'd11; a_sign1 = 4'd10; a_sign2 = 4'd14; a_sign3 = 4'd7;
b_sign0 = 4'd12; b_sign1 = 4'd5; b_sign2 = 4'd13; b_sign3 = 4'd8;
@(posedge clk_i);
a_mant0 = 8'd9; a_mant1 = 8'd238; a_mant2 = 8'd92; a_mant3 = 8'd6;
b_mant0 = 8'd24; b_mant1 = 8'd108; b_mant2 = 8'd183; b_mant3 = 8'd240;
a_exp0 = 10'd412; a_exp1 = 10'd438; a_exp2 = 10'd441; a_exp3 = 10'd729;
b_exp0 = 10'd196; b_exp1 = 10'd1002; b_exp2 = 10'd101; b_exp3 = 10'd807;
a_sign0 = 4'd10; a_sign1 = 4'd16; a_sign2 = 4'd2; a_sign3 = 4'd11;
b_sign0 = 4'd10; b_sign1 = 4'd11; b_sign2 = 4'd0; b_sign3 = 4'd9;
@(posedge clk_i);
a_mant0 = 8'd59; a_mant1 = 8'd193; a_mant2 = 8'd97; a_mant3 = 8'd152;
b_mant0 = 8'd137; b_mant1 = 8'd21; b_mant2 = 8'd74; b_mant3 = 8'd209;
a_exp0 = 10'd92; a_exp1 = 10'd582; a_exp2 = 10'd829; a_exp3 = 10'd547;
b_exp0 = 10'd786; b_exp1 = 10'd236; b_exp2 = 10'd326; b_exp3 = 10'd540;
a_sign0 = 4'd16; a_sign1 = 4'd6; a_sign2 = 4'd6; a_sign3 = 4'd2;
b_sign0 = 4'd5; b_sign1 = 4'd2; b_sign2 = 4'd10; b_sign3 = 4'd7;
@(posedge clk_i);
a_mant0 = 8'd183; a_mant1 = 8'd10; a_mant2 = 8'd21; a_mant3 = 8'd158;
b_mant0 = 8'd34; b_mant1 = 8'd3; b_mant2 = 8'd233; b_mant3 = 8'd124;
a_exp0 = 10'd760; a_exp1 = 10'd272; a_exp2 = 10'd496; a_exp3 = 10'd734;
b_exp0 = 10'd260; b_exp1 = 10'd349; b_exp2 = 10'd575; b_exp3 = 10'd343;
a_sign0 = 4'd15; a_sign1 = 4'd15; a_sign2 = 4'd0; a_sign3 = 4'd1;
b_sign0 = 4'd5; b_sign1 = 4'd15; b_sign2 = 4'd1; b_sign3 = 4'd12;
@(posedge clk_i);
a_mant0 = 8'd247; a_mant1 = 8'd57; a_mant2 = 8'd12; a_mant3 = 8'd178;
b_mant0 = 8'd238; b_mant1 = 8'd102; b_mant2 = 8'd142; b_mant3 = 8'd45;
a_exp0 = 10'd280; a_exp1 = 10'd981; a_exp2 = 10'd583; a_exp3 = 10'd371;
b_exp0 = 10'd114; b_exp1 = 10'd714; b_exp2 = 10'd574; b_exp3 = 10'd189;
a_sign0 = 4'd8; a_sign1 = 4'd13; a_sign2 = 4'd7; a_sign3 = 4'd6;
b_sign0 = 4'd16; b_sign1 = 4'd2; b_sign2 = 4'd8; b_sign3 = 4'd15;
@(posedge clk_i);
a_mant0 = 8'd214; a_mant1 = 8'd177; a_mant2 = 8'd63; a_mant3 = 8'd111;
b_mant0 = 8'd67; b_mant1 = 8'd56; b_mant2 = 8'd68; b_mant3 = 8'd86;
a_exp0 = 10'd367; a_exp1 = 10'd714; a_exp2 = 10'd840; a_exp3 = 10'd210;
b_exp0 = 10'd494; b_exp1 = 10'd720; b_exp2 = 10'd930; b_exp3 = 10'd138;
a_sign0 = 4'd13; a_sign1 = 4'd16; a_sign2 = 4'd9; a_sign3 = 4'd5;
b_sign0 = 4'd10; b_sign1 = 4'd4; b_sign2 = 4'd7; b_sign3 = 4'd6;
@(posedge clk_i);
a_mant0 = 8'd252; a_mant1 = 8'd35; a_mant2 = 8'd245; a_mant3 = 8'd67;
b_mant0 = 8'd245; b_mant1 = 8'd50; b_mant2 = 8'd197; b_mant3 = 8'd134;
a_exp0 = 10'd943; a_exp1 = 10'd238; a_exp2 = 10'd689; a_exp3 = 10'd395;
b_exp0 = 10'd84; b_exp1 = 10'd48; b_exp2 = 10'd112; b_exp3 = 10'd305;
a_sign0 = 4'd1; a_sign1 = 4'd11; a_sign2 = 4'd15; a_sign3 = 4'd15;
b_sign0 = 4'd1; b_sign1 = 4'd13; b_sign2 = 4'd7; b_sign3 = 4'd11;
@(posedge clk_i);
a_mant0 = 8'd73; a_mant1 = 8'd177; a_mant2 = 8'd39; a_mant3 = 8'd242;
b_mant0 = 8'd155; b_mant1 = 8'd179; b_mant2 = 8'd162; b_mant3 = 8'd18;
a_exp0 = 10'd81; a_exp1 = 10'd290; a_exp2 = 10'd356; a_exp3 = 10'd359;
b_exp0 = 10'd197; b_exp1 = 10'd635; b_exp2 = 10'd962; b_exp3 = 10'd310;
a_sign0 = 4'd13; a_sign1 = 4'd9; a_sign2 = 4'd4; a_sign3 = 4'd8;
b_sign0 = 4'd5; b_sign1 = 4'd6; b_sign2 = 4'd15; b_sign3 = 4'd12;
@(posedge clk_i);
shared_exps0 = 8'd129;
shared_exps1 = 8'd143;
rstn = 0;
@(posedge clk_i);
rstn = 1;
a_mant0 = 8'd126; a_mant1 = 8'd172; a_mant2 = 8'd178; a_mant3 = 8'd17;
b_mant0 = 8'd98; b_mant1 = 8'd12; b_mant2 = 8'd66; b_mant3 = 8'd174;
a_exp0 = 10'd374; a_exp1 = 10'd220; a_exp2 = 10'd691; a_exp3 = 10'd71;
b_exp0 = 10'd98; b_exp1 = 10'd1008; b_exp2 = 10'd178; b_exp3 = 10'd13;
a_sign0 = 4'd7; a_sign1 = 4'd6; a_sign2 = 4'd15; a_sign3 = 4'd15;
b_sign0 = 4'd10; b_sign1 = 4'd8; b_sign2 = 4'd14; b_sign3 = 4'd0;
@(posedge clk_i);
a_mant0 = 8'd169; a_mant1 = 8'd123; a_mant2 = 8'd64; a_mant3 = 8'd51;
b_mant0 = 8'd224; b_mant1 = 8'd213; b_mant2 = 8'd189; b_mant3 = 8'd28;
a_exp0 = 10'd194; a_exp1 = 10'd966; a_exp2 = 10'd864; a_exp3 = 10'd1008;
b_exp0 = 10'd525; b_exp1 = 10'd405; b_exp2 = 10'd526; b_exp3 = 10'd426;
a_sign0 = 4'd0; a_sign1 = 4'd0; a_sign2 = 4'd0; a_sign3 = 4'd6;
b_sign0 = 4'd16; b_sign1 = 4'd8; b_sign2 = 4'd3; b_sign3 = 4'd14;
@(posedge clk_i);
a_mant0 = 8'd153; a_mant1 = 8'd53; a_mant2 = 8'd100; a_mant3 = 8'd209;
b_mant0 = 8'd56; b_mant1 = 8'd237; b_mant2 = 8'd17; b_mant3 = 8'd135;
a_exp0 = 10'd391; a_exp1 = 10'd996; a_exp2 = 10'd419; a_exp3 = 10'd93;
b_exp0 = 10'd933; b_exp1 = 10'd69; b_exp2 = 10'd50; b_exp3 = 10'd376;
a_sign0 = 4'd12; a_sign1 = 4'd4; a_sign2 = 4'd1; a_sign3 = 4'd8;
b_sign0 = 4'd8; b_sign1 = 4'd9; b_sign2 = 4'd12; b_sign3 = 4'd13;
@(posedge clk_i);
a_mant0 = 8'd91; a_mant1 = 8'd229; a_mant2 = 8'd18; a_mant3 = 8'd141;
b_mant0 = 8'd4; b_mant1 = 8'd141; b_mant2 = 8'd210; b_mant3 = 8'd136;
a_exp0 = 10'd322; a_exp1 = 10'd125; a_exp2 = 10'd821; a_exp3 = 10'd552;
b_exp0 = 10'd741; b_exp1 = 10'd851; b_exp2 = 10'd31; b_exp3 = 10'd346;
a_sign0 = 4'd15; a_sign1 = 4'd0; a_sign2 = 4'd2; a_sign3 = 4'd9;
b_sign0 = 4'd10; b_sign1 = 4'd11; b_sign2 = 4'd1; b_sign3 = 4'd3;
@(posedge clk_i);
a_mant0 = 8'd146; a_mant1 = 8'd241; a_mant2 = 8'd25; a_mant3 = 8'd211;
b_mant0 = 8'd55; b_mant1 = 8'd95; b_mant2 = 8'd74; b_mant3 = 8'd80;
a_exp0 = 10'd18; a_exp1 = 10'd490; a_exp2 = 10'd202; a_exp3 = 10'd833;
b_exp0 = 10'd801; b_exp1 = 10'd495; b_exp2 = 10'd956; b_exp3 = 10'd518;
a_sign0 = 4'd3; a_sign1 = 4'd4; a_sign2 = 4'd14; a_sign3 = 4'd11;
b_sign0 = 4'd16; b_sign1 = 4'd15; b_sign2 = 4'd7; b_sign3 = 4'd13;
@(posedge clk_i);
a_mant0 = 8'd72; a_mant1 = 8'd127; a_mant2 = 8'd16; a_mant3 = 8'd68;
b_mant0 = 8'd90; b_mant1 = 8'd135; b_mant2 = 8'd9; b_mant3 = 8'd220;
a_exp0 = 10'd170; a_exp1 = 10'd37; a_exp2 = 10'd181; a_exp3 = 10'd615;
b_exp0 = 10'd587; b_exp1 = 10'd831; b_exp2 = 10'd282; b_exp3 = 10'd534;
a_sign0 = 4'd2; a_sign1 = 4'd14; a_sign2 = 4'd11; a_sign3 = 4'd4;
b_sign0 = 4'd15; b_sign1 = 4'd6; b_sign2 = 4'd16; b_sign3 = 4'd1;
@(posedge clk_i);
a_mant0 = 8'd169; a_mant1 = 8'd106; a_mant2 = 8'd143; a_mant3 = 8'd240;
b_mant0 = 8'd13; b_mant1 = 8'd92; b_mant2 = 8'd48; b_mant3 = 8'd68;
a_exp0 = 10'd467; a_exp1 = 10'd87; a_exp2 = 10'd799; a_exp3 = 10'd707;
b_exp0 = 10'd701; b_exp1 = 10'd719; b_exp2 = 10'd572; b_exp3 = 10'd818;
a_sign0 = 4'd9; a_sign1 = 4'd3; a_sign2 = 4'd14; a_sign3 = 4'd9;
b_sign0 = 4'd2; b_sign1 = 4'd9; b_sign2 = 4'd16; b_sign3 = 4'd9;
@(posedge clk_i);
shared_exps0 = 8'd120;
shared_exps1 = 8'd133;
a_mant0 = 8'd91; a_mant1 = 8'd160; a_mant2 = 8'd250; a_mant3 = 8'd110;
b_mant0 = 8'd109; b_mant1 = 8'd123; b_mant2 = 8'd232; b_mant3 = 8'd14;
a_exp0 = 10'd1022; a_exp1 = 10'd114; a_exp2 = 10'd519; a_exp3 = 10'd844;
b_exp0 = 10'd820; b_exp1 = 10'd6; b_exp2 = 10'd545; b_exp3 = 10'd509;
a_sign0 = 4'd16; a_sign1 = 4'd6; a_sign2 = 4'd6; a_sign3 = 4'd0;
b_sign0 = 4'd5; b_sign1 = 4'd1; b_sign2 = 4'd2; b_sign3 = 4'd16;
@(posedge clk_i);
a_mant0 = 8'd193; a_mant1 = 8'd7; a_mant2 = 8'd149; a_mant3 = 8'd251;
b_mant0 = 8'd77; b_mant1 = 8'd184; b_mant2 = 8'd103; b_mant3 = 8'd63;
a_exp0 = 10'd639; a_exp1 = 10'd406; a_exp2 = 10'd59; a_exp3 = 10'd611;
b_exp0 = 10'd693; b_exp1 = 10'd1021; b_exp2 = 10'd1019; b_exp3 = 10'd961;
a_sign0 = 4'd15; a_sign1 = 4'd10; a_sign2 = 4'd0; a_sign3 = 4'd11;
b_sign0 = 4'd4; b_sign1 = 4'd11; b_sign2 = 4'd7; b_sign3 = 4'd0;
@(posedge clk_i);
a_mant0 = 8'd189; a_mant1 = 8'd120; a_mant2 = 8'd78; a_mant3 = 8'd217;
b_mant0 = 8'd132; b_mant1 = 8'd211; b_mant2 = 8'd71; b_mant3 = 8'd119;
a_exp0 = 10'd613; a_exp1 = 10'd335; a_exp2 = 10'd556; a_exp3 = 10'd108;
b_exp0 = 10'd934; b_exp1 = 10'd183; b_exp2 = 10'd37; b_exp3 = 10'd990;
a_sign0 = 4'd0; a_sign1 = 4'd3; a_sign2 = 4'd4; a_sign3 = 4'd9;
b_sign0 = 4'd14; b_sign1 = 4'd6; b_sign2 = 4'd10; b_sign3 = 4'd4;
@(posedge clk_i);
a_mant0 = 8'd118; a_mant1 = 8'd175; a_mant2 = 8'd223; a_mant3 = 8'd16;
b_mant0 = 8'd68; b_mant1 = 8'd26; b_mant2 = 8'd211; b_mant3 = 8'd187;
a_exp0 = 10'd969; a_exp1 = 10'd760; a_exp2 = 10'd112; a_exp3 = 10'd497;
b_exp0 = 10'd343; b_exp1 = 10'd385; b_exp2 = 10'd216; b_exp3 = 10'd813;
a_sign0 = 4'd2; a_sign1 = 4'd10; a_sign2 = 4'd0; a_sign3 = 4'd1;
b_sign0 = 4'd15; b_sign1 = 4'd11; b_sign2 = 4'd13; b_sign3 = 4'd3;
@(posedge clk_i);
a_mant0 = 8'd103; a_mant1 = 8'd121; a_mant2 = 8'd168; a_mant3 = 8'd32;
b_mant0 = 8'd189; b_mant1 = 8'd148; b_mant2 = 8'd168; b_mant3 = 8'd210;
a_exp0 = 10'd707; a_exp1 = 10'd285; a_exp2 = 10'd76; a_exp3 = 10'd989;
b_exp0 = 10'd948; b_exp1 = 10'd962; b_exp2 = 10'd339; b_exp3 = 10'd829;
a_sign0 = 4'd5; a_sign1 = 4'd14; a_sign2 = 4'd8; a_sign3 = 4'd16;
b_sign0 = 4'd13; b_sign1 = 4'd7; b_sign2 = 4'd15; b_sign3 = 4'd14;
@(posedge clk_i);
a_mant0 = 8'd231; a_mant1 = 8'd103; a_mant2 = 8'd181; a_mant3 = 8'd131;
b_mant0 = 8'd87; b_mant1 = 8'd110; b_mant2 = 8'd213; b_mant3 = 8'd60;
a_exp0 = 10'd336; a_exp1 = 10'd821; a_exp2 = 10'd647; a_exp3 = 10'd306;
b_exp0 = 10'd826; b_exp1 = 10'd800; b_exp2 = 10'd220; b_exp3 = 10'd742;
a_sign0 = 4'd11; a_sign1 = 4'd14; a_sign2 = 4'd6; a_sign3 = 4'd6;
b_sign0 = 4'd10; b_sign1 = 4'd11; b_sign2 = 4'd1; b_sign3 = 4'd7;
@(posedge clk_i);
a_mant0 = 8'd130; a_mant1 = 8'd30; a_mant2 = 8'd14; a_mant3 = 8'd35;
b_mant0 = 8'd6; b_mant1 = 8'd43; b_mant2 = 8'd162; b_mant3 = 8'd195;
a_exp0 = 10'd851; a_exp1 = 10'd1003; a_exp2 = 10'd491; a_exp3 = 10'd497;
b_exp0 = 10'd561; b_exp1 = 10'd300; b_exp2 = 10'd367; b_exp3 = 10'd954;
a_sign0 = 4'd4; a_sign1 = 4'd7; a_sign2 = 4'd10; a_sign3 = 4'd6;
b_sign0 = 4'd11; b_sign1 = 4'd16; b_sign2 = 4'd7; b_sign3 = 4'd6;
@(posedge clk_i);
a_mant0 = 8'd99; a_mant1 = 8'd9; a_mant2 = 8'd188; a_mant3 = 8'd48;
b_mant0 = 8'd248; b_mant1 = 8'd100; b_mant2 = 8'd99; b_mant3 = 8'd185;
a_exp0 = 10'd282; a_exp1 = 10'd87; a_exp2 = 10'd940; a_exp3 = 10'd490;
b_exp0 = 10'd910; b_exp1 = 10'd80; b_exp2 = 10'd334; b_exp3 = 10'd109;
a_sign0 = 4'd12; a_sign1 = 4'd3; a_sign2 = 4'd8; a_sign3 = 4'd3;
b_sign0 = 4'd8; b_sign1 = 4'd10; b_sign2 = 4'd11; b_sign3 = 4'd8;
@(posedge clk_i);
shared_exps0 = 8'd112;
shared_exps1 = 8'd102;
a_mant0 = 8'd31; a_mant1 = 8'd126; a_mant2 = 8'd53; a_mant3 = 8'd15;
b_mant0 = 8'd104; b_mant1 = 8'd13; b_mant2 = 8'd228; b_mant3 = 8'd92;
a_exp0 = 10'd751; a_exp1 = 10'd447; a_exp2 = 10'd331; a_exp3 = 10'd488;
b_exp0 = 10'd154; b_exp1 = 10'd941; b_exp2 = 10'd387; b_exp3 = 10'd664;
a_sign0 = 4'd3; a_sign1 = 4'd10; a_sign2 = 4'd16; a_sign3 = 4'd8;
b_sign0 = 4'd4; b_sign1 = 4'd12; b_sign2 = 4'd1; b_sign3 = 4'd3;
@(posedge clk_i);
a_mant0 = 8'd30; a_mant1 = 8'd33; a_mant2 = 8'd159; a_mant3 = 8'd83;
b_mant0 = 8'd146; b_mant1 = 8'd185; b_mant2 = 8'd72; b_mant3 = 8'd179;
a_exp0 = 10'd117; a_exp1 = 10'd384; a_exp2 = 10'd919; a_exp3 = 10'd1019;
b_exp0 = 10'd454; b_exp1 = 10'd743; b_exp2 = 10'd608; b_exp3 = 10'd876;
a_sign0 = 4'd12; a_sign1 = 4'd7; a_sign2 = 4'd7; a_sign3 = 4'd11;
b_sign0 = 4'd12; b_sign1 = 4'd3; b_sign2 = 4'd0; b_sign3 = 4'd5;
@(posedge clk_i);
a_mant0 = 8'd162; a_mant1 = 8'd94; a_mant2 = 8'd186; a_mant3 = 8'd14;
b_mant0 = 8'd129; b_mant1 = 8'd198; b_mant2 = 8'd24; b_mant3 = 8'd67;
a_exp0 = 10'd382; a_exp1 = 10'd364; a_exp2 = 10'd607; a_exp3 = 10'd902;
b_exp0 = 10'd753; b_exp1 = 10'd851; b_exp2 = 10'd82; b_exp3 = 10'd298;
a_sign0 = 4'd0; a_sign1 = 4'd9; a_sign2 = 4'd4; a_sign3 = 4'd1;
b_sign0 = 4'd13; b_sign1 = 4'd5; b_sign2 = 4'd11; b_sign3 = 4'd9;
@(posedge clk_i);
a_mant0 = 8'd208; a_mant1 = 8'd109; a_mant2 = 8'd228; a_mant3 = 8'd207;
b_mant0 = 8'd65; b_mant1 = 8'd205; b_mant2 = 8'd43; b_mant3 = 8'd189;
a_exp0 = 10'd154; a_exp1 = 10'd636; a_exp2 = 10'd588; a_exp3 = 10'd99;
b_exp0 = 10'd123; b_exp1 = 10'd275; b_exp2 = 10'd271; b_exp3 = 10'd961;
a_sign0 = 4'd2; a_sign1 = 4'd6; a_sign2 = 4'd9; a_sign3 = 4'd2;
b_sign0 = 4'd1; b_sign1 = 4'd3; b_sign2 = 4'd1; b_sign3 = 4'd8;
@(posedge clk_i);
a_mant0 = 8'd166; a_mant1 = 8'd73; a_mant2 = 8'd109; a_mant3 = 8'd84;
b_mant0 = 8'd34; b_mant1 = 8'd109; b_mant2 = 8'd134; b_mant3 = 8'd205;
a_exp0 = 10'd633; a_exp1 = 10'd938; a_exp2 = 10'd503; a_exp3 = 10'd240;
b_exp0 = 10'd108; b_exp1 = 10'd401; b_exp2 = 10'd470; b_exp3 = 10'd231;
a_sign0 = 4'd15; a_sign1 = 4'd11; a_sign2 = 4'd15; a_sign3 = 4'd6;
b_sign0 = 4'd14; b_sign1 = 4'd3; b_sign2 = 4'd14; b_sign3 = 4'd14;
@(posedge clk_i);
a_mant0 = 8'd59; a_mant1 = 8'd238; a_mant2 = 8'd244; a_mant3 = 8'd137;
b_mant0 = 8'd188; b_mant1 = 8'd103; b_mant2 = 8'd223; b_mant3 = 8'd216;
a_exp0 = 10'd7; a_exp1 = 10'd407; a_exp2 = 10'd1000; a_exp3 = 10'd639;
b_exp0 = 10'd397; b_exp1 = 10'd136; b_exp2 = 10'd815; b_exp3 = 10'd955;
a_sign0 = 4'd8; a_sign1 = 4'd6; a_sign2 = 4'd6; a_sign3 = 4'd3;
b_sign0 = 4'd10; b_sign1 = 4'd13; b_sign2 = 4'd1; b_sign3 = 4'd1;
@(posedge clk_i);
a_mant0 = 8'd216; a_mant1 = 8'd96; a_mant2 = 8'd115; a_mant3 = 8'd48;
b_mant0 = 8'd152; b_mant1 = 8'd216; b_mant2 = 8'd241; b_mant3 = 8'd223;
a_exp0 = 10'd753; a_exp1 = 10'd803; a_exp2 = 10'd506; a_exp3 = 10'd135;
b_exp0 = 10'd696; b_exp1 = 10'd191; b_exp2 = 10'd454; b_exp3 = 10'd1017;
a_sign0 = 4'd2; a_sign1 = 4'd11; a_sign2 = 4'd12; a_sign3 = 4'd13;
b_sign0 = 4'd10; b_sign1 = 4'd12; b_sign2 = 4'd6; b_sign3 = 4'd9;
@(posedge clk_i);
a_mant0 = 8'd182; a_mant1 = 8'd96; a_mant2 = 8'd213; a_mant3 = 8'd199;
b_mant0 = 8'd105; b_mant1 = 8'd18; b_mant2 = 8'd127; b_mant3 = 8'd19;
a_exp0 = 10'd295; a_exp1 = 10'd807; a_exp2 = 10'd810; a_exp3 = 10'd791;
b_exp0 = 10'd2; b_exp1 = 10'd201; b_exp2 = 10'd687; b_exp3 = 10'd637;
a_sign0 = 4'd4; a_sign1 = 4'd14; a_sign2 = 4'd13; a_sign3 = 4'd13;
b_sign0 = 4'd10; b_sign1 = 4'd9; b_sign2 = 4'd4; b_sign3 = 4'd14;
@(posedge clk_i);
shared_exps0 = 8'd149;
shared_exps1 = 8'd114;
a_mant0 = 8'd14; a_mant1 = 8'd199; a_mant2 = 8'd187; a_mant3 = 8'd21;
b_mant0 = 8'd112; b_mant1 = 8'd225; b_mant2 = 8'd14; b_mant3 = 8'd234;
a_exp0 = 10'd146; a_exp1 = 10'd555; a_exp2 = 10'd694; a_exp3 = 10'd413;
b_exp0 = 10'd114; b_exp1 = 10'd149; b_exp2 = 10'd46; b_exp3 = 10'd911;
a_sign0 = 4'd8; a_sign1 = 4'd2; a_sign2 = 4'd11; a_sign3 = 4'd0;
b_sign0 = 4'd8; b_sign1 = 4'd8; b_sign2 = 4'd11; b_sign3 = 4'd1;
@(posedge clk_i);
a_mant0 = 8'd152; a_mant1 = 8'd244; a_mant2 = 8'd63; a_mant3 = 8'd131;
b_mant0 = 8'd166; b_mant1 = 8'd212; b_mant2 = 8'd157; b_mant3 = 8'd28;
a_exp0 = 10'd422; a_exp1 = 10'd484; a_exp2 = 10'd152; a_exp3 = 10'd302;
b_exp0 = 10'd570; b_exp1 = 10'd389; b_exp2 = 10'd1002; b_exp3 = 10'd473;
a_sign0 = 4'd9; a_sign1 = 4'd8; a_sign2 = 4'd1; a_sign3 = 4'd16;
b_sign0 = 4'd1; b_sign1 = 4'd16; b_sign2 = 4'd1; b_sign3 = 4'd14;
@(posedge clk_i);
a_mant0 = 8'd66; a_mant1 = 8'd104; a_mant2 = 8'd99; a_mant3 = 8'd172;
b_mant0 = 8'd78; b_mant1 = 8'd110; b_mant2 = 8'd215; b_mant3 = 8'd191;
a_exp0 = 10'd703; a_exp1 = 10'd676; a_exp2 = 10'd732; a_exp3 = 10'd382;
b_exp0 = 10'd588; b_exp1 = 10'd109; b_exp2 = 10'd1002; b_exp3 = 10'd473;
a_sign0 = 4'd3; a_sign1 = 4'd14; a_sign2 = 4'd15; a_sign3 = 4'd3;
b_sign0 = 4'd10; b_sign1 = 4'd2; b_sign2 = 4'd3; b_sign3 = 4'd5;
@(posedge clk_i);
a_mant0 = 8'd228; a_mant1 = 8'd127; a_mant2 = 8'd144; a_mant3 = 8'd195;
b_mant0 = 8'd211; b_mant1 = 8'd173; b_mant2 = 8'd8; b_mant3 = 8'd187;
a_exp0 = 10'd344; a_exp1 = 10'd858; a_exp2 = 10'd658; a_exp3 = 10'd781;
b_exp0 = 10'd299; b_exp1 = 10'd921; b_exp2 = 10'd355; b_exp3 = 10'd553;
a_sign0 = 4'd4; a_sign1 = 4'd8; a_sign2 = 4'd0; a_sign3 = 4'd1;
b_sign0 = 4'd7; b_sign1 = 4'd1; b_sign2 = 4'd11; b_sign3 = 4'd3;
@(posedge clk_i);
a_mant0 = 8'd125; a_mant1 = 8'd214; a_mant2 = 8'd124; a_mant3 = 8'd131;
b_mant0 = 8'd35; b_mant1 = 8'd77; b_mant2 = 8'd214; b_mant3 = 8'd16;
a_exp0 = 10'd171; a_exp1 = 10'd339; a_exp2 = 10'd489; a_exp3 = 10'd997;
b_exp0 = 10'd882; b_exp1 = 10'd137; b_exp2 = 10'd675; b_exp3 = 10'd872;
a_sign0 = 4'd16; a_sign1 = 4'd11; a_sign2 = 4'd5; a_sign3 = 4'd4;
b_sign0 = 4'd3; b_sign1 = 4'd12; b_sign2 = 4'd12; b_sign3 = 4'd10;
@(posedge clk_i);
a_mant0 = 8'd148; a_mant1 = 8'd208; a_mant2 = 8'd13; a_mant3 = 8'd184;
b_mant0 = 8'd170; b_mant1 = 8'd2; b_mant2 = 8'd104; b_mant3 = 8'd75;
a_exp0 = 10'd593; a_exp1 = 10'd662; a_exp2 = 10'd867; a_exp3 = 10'd135;
b_exp0 = 10'd93; b_exp1 = 10'd831; b_exp2 = 10'd438; b_exp3 = 10'd430;
a_sign0 = 4'd1; a_sign1 = 4'd0; a_sign2 = 4'd6; a_sign3 = 4'd6;
b_sign0 = 4'd6; b_sign1 = 4'd0; b_sign2 = 4'd12; b_sign3 = 4'd11;
@(posedge clk_i);
a_mant0 = 8'd58; a_mant1 = 8'd102; a_mant2 = 8'd222; a_mant3 = 8'd10;
b_mant0 = 8'd2; b_mant1 = 8'd154; b_mant2 = 8'd216; b_mant3 = 8'd140;
a_exp0 = 10'd330; a_exp1 = 10'd686; a_exp2 = 10'd558; a_exp3 = 10'd116;
b_exp0 = 10'd485; b_exp1 = 10'd952; b_exp2 = 10'd597; b_exp3 = 10'd602;
a_sign0 = 4'd13; a_sign1 = 4'd5; a_sign2 = 4'd14; a_sign3 = 4'd5;
b_sign0 = 4'd15; b_sign1 = 4'd10; b_sign2 = 4'd0; b_sign3 = 4'd9;
@(posedge clk_i);
a_mant0 = 8'd212; a_mant1 = 8'd206; a_mant2 = 8'd217; a_mant3 = 8'd224;
b_mant0 = 8'd181; b_mant1 = 8'd57; b_mant2 = 8'd103; b_mant3 = 8'd242;
a_exp0 = 10'd937; a_exp1 = 10'd339; a_exp2 = 10'd323; a_exp3 = 10'd431;
b_exp0 = 10'd479; b_exp1 = 10'd359; b_exp2 = 10'd712; b_exp3 = 10'd985;
a_sign0 = 4'd5; a_sign1 = 4'd12; a_sign2 = 4'd16; a_sign3 = 4'd9;
b_sign0 = 4'd5; b_sign1 = 4'd3; b_sign2 = 4'd9; b_sign3 = 4'd1;
@(posedge clk_i);
shared_exps0 = 8'd142;
shared_exps1 = 8'd129;
rstn = 0;
@(posedge clk_i);
rstn = 1;
a_mant0 = 8'd107; a_mant1 = 8'd119; a_mant2 = 8'd252; a_mant3 = 8'd63;
b_mant0 = 8'd115; b_mant1 = 8'd84; b_mant2 = 8'd172; b_mant3 = 8'd204;
a_exp0 = 10'd957; a_exp1 = 10'd48; a_exp2 = 10'd72; a_exp3 = 10'd42;
b_exp0 = 10'd485; b_exp1 = 10'd321; b_exp2 = 10'd869; b_exp3 = 10'd683;
a_sign0 = 4'd16; a_sign1 = 4'd13; a_sign2 = 4'd0; a_sign3 = 4'd11;
b_sign0 = 4'd3; b_sign1 = 4'd2; b_sign2 = 4'd4; b_sign3 = 4'd8;
@(posedge clk_i);
a_mant0 = 8'd33; a_mant1 = 8'd175; a_mant2 = 8'd190; a_mant3 = 8'd47;
b_mant0 = 8'd155; b_mant1 = 8'd230; b_mant2 = 8'd6; b_mant3 = 8'd194;
a_exp0 = 10'd9; a_exp1 = 10'd446; a_exp2 = 10'd903; a_exp3 = 10'd31;
b_exp0 = 10'd626; b_exp1 = 10'd65; b_exp2 = 10'd444; b_exp3 = 10'd132;
a_sign0 = 4'd7; a_sign1 = 4'd10; a_sign2 = 4'd10; a_sign3 = 4'd1;
b_sign0 = 4'd7; b_sign1 = 4'd14; b_sign2 = 4'd11; b_sign3 = 4'd2;
@(posedge clk_i);
a_mant0 = 8'd79; a_mant1 = 8'd124; a_mant2 = 8'd101; a_mant3 = 8'd36;
b_mant0 = 8'd210; b_mant1 = 8'd171; b_mant2 = 8'd46; b_mant3 = 8'd65;
a_exp0 = 10'd822; a_exp1 = 10'd859; a_exp2 = 10'd762; a_exp3 = 10'd926;
b_exp0 = 10'd353; b_exp1 = 10'd476; b_exp2 = 10'd790; b_exp3 = 10'd572;
a_sign0 = 4'd5; a_sign1 = 4'd11; a_sign2 = 4'd6; a_sign3 = 4'd1;
b_sign0 = 4'd12; b_sign1 = 4'd5; b_sign2 = 4'd12; b_sign3 = 4'd8;
@(posedge clk_i);
a_mant0 = 8'd85; a_mant1 = 8'd92; a_mant2 = 8'd162; a_mant3 = 8'd214;
b_mant0 = 8'd30; b_mant1 = 8'd63; b_mant2 = 8'd228; b_mant3 = 8'd146;
a_exp0 = 10'd68; a_exp1 = 10'd592; a_exp2 = 10'd716; a_exp3 = 10'd656;
b_exp0 = 10'd722; b_exp1 = 10'd712; b_exp2 = 10'd414; b_exp3 = 10'd845;
a_sign0 = 4'd6; a_sign1 = 4'd12; a_sign2 = 4'd15; a_sign3 = 4'd12;
b_sign0 = 4'd8; b_sign1 = 4'd1; b_sign2 = 4'd12; b_sign3 = 4'd11;
@(posedge clk_i);
a_mant0 = 8'd2; a_mant1 = 8'd43; a_mant2 = 8'd209; a_mant3 = 8'd147;
b_mant0 = 8'd132; b_mant1 = 8'd139; b_mant2 = 8'd187; b_mant3 = 8'd205;
a_exp0 = 10'd674; a_exp1 = 10'd998; a_exp2 = 10'd460; a_exp3 = 10'd302;
b_exp0 = 10'd341; b_exp1 = 10'd360; b_exp2 = 10'd1023; b_exp3 = 10'd391;
a_sign0 = 4'd6; a_sign1 = 4'd0; a_sign2 = 4'd8; a_sign3 = 4'd7;
b_sign0 = 4'd8; b_sign1 = 4'd2; b_sign2 = 4'd16; b_sign3 = 4'd4;
@(posedge clk_i);
a_mant0 = 8'd10; a_mant1 = 8'd105; a_mant2 = 8'd96; a_mant3 = 8'd105;
b_mant0 = 8'd8; b_mant1 = 8'd225; b_mant2 = 8'd195; b_mant3 = 8'd13;
a_exp0 = 10'd974; a_exp1 = 10'd414; a_exp2 = 10'd405; a_exp3 = 10'd182;
b_exp0 = 10'd559; b_exp1 = 10'd962; b_exp2 = 10'd775; b_exp3 = 10'd995;
a_sign0 = 4'd9; a_sign1 = 4'd4; a_sign2 = 4'd9; a_sign3 = 4'd10;
b_sign0 = 4'd10; b_sign1 = 4'd3; b_sign2 = 4'd13; b_sign3 = 4'd8;
@(posedge clk_i);
a_mant0 = 8'd162; a_mant1 = 8'd208; a_mant2 = 8'd141; a_mant3 = 8'd54;
b_mant0 = 8'd144; b_mant1 = 8'd48; b_mant2 = 8'd33; b_mant3 = 8'd60;
a_exp0 = 10'd986; a_exp1 = 10'd272; a_exp2 = 10'd410; a_exp3 = 10'd140;
b_exp0 = 10'd351; b_exp1 = 10'd503; b_exp2 = 10'd922; b_exp3 = 10'd516;
a_sign0 = 4'd12; a_sign1 = 4'd5; a_sign2 = 4'd11; a_sign3 = 4'd14;
b_sign0 = 4'd11; b_sign1 = 4'd9; b_sign2 = 4'd3; b_sign3 = 4'd6;
@(posedge clk_i);
shared_exps0 = 8'd127;
shared_exps1 = 8'd149;
a_mant0 = 8'd243; a_mant1 = 8'd17; a_mant2 = 8'd213; a_mant3 = 8'd63;
b_mant0 = 8'd26; b_mant1 = 8'd5; b_mant2 = 8'd182; b_mant3 = 8'd141;
a_exp0 = 10'd103; a_exp1 = 10'd48; a_exp2 = 10'd457; a_exp3 = 10'd656;
b_exp0 = 10'd732; b_exp1 = 10'd284; b_exp2 = 10'd645; b_exp3 = 10'd388;
a_sign0 = 4'd1; a_sign1 = 4'd15; a_sign2 = 4'd4; a_sign3 = 4'd9;
b_sign0 = 4'd11; b_sign1 = 4'd5; b_sign2 = 4'd0; b_sign3 = 4'd8;
@(posedge clk_i);
a_mant0 = 8'd56; a_mant1 = 8'd174; a_mant2 = 8'd236; a_mant3 = 8'd170;
b_mant0 = 8'd233; b_mant1 = 8'd27; b_mant2 = 8'd102; b_mant3 = 8'd143;
a_exp0 = 10'd311; a_exp1 = 10'd829; a_exp2 = 10'd441; a_exp3 = 10'd381;
b_exp0 = 10'd676; b_exp1 = 10'd61; b_exp2 = 10'd635; b_exp3 = 10'd863;
a_sign0 = 4'd9; a_sign1 = 4'd13; a_sign2 = 4'd0; a_sign3 = 4'd6;
b_sign0 = 4'd10; b_sign1 = 4'd14; b_sign2 = 4'd2; b_sign3 = 4'd2;
@(posedge clk_i);
a_mant0 = 8'd65; a_mant1 = 8'd15; a_mant2 = 8'd209; a_mant3 = 8'd132;
b_mant0 = 8'd130; b_mant1 = 8'd190; b_mant2 = 8'd199; b_mant3 = 8'd99;
a_exp0 = 10'd778; a_exp1 = 10'd236; a_exp2 = 10'd493; a_exp3 = 10'd526;
b_exp0 = 10'd726; b_exp1 = 10'd716; b_exp2 = 10'd912; b_exp3 = 10'd519;
a_sign0 = 4'd1; a_sign1 = 4'd12; a_sign2 = 4'd0; a_sign3 = 4'd4;
b_sign0 = 4'd4; b_sign1 = 4'd0; b_sign2 = 4'd6; b_sign3 = 4'd4;
@(posedge clk_i);
a_mant0 = 8'd179; a_mant1 = 8'd253; a_mant2 = 8'd113; a_mant3 = 8'd23;
b_mant0 = 8'd245; b_mant1 = 8'd149; b_mant2 = 8'd187; b_mant3 = 8'd113;
a_exp0 = 10'd465; a_exp1 = 10'd374; a_exp2 = 10'd637; a_exp3 = 10'd420;
b_exp0 = 10'd118; b_exp1 = 10'd688; b_exp2 = 10'd595; b_exp3 = 10'd737;
a_sign0 = 4'd5; a_sign1 = 4'd14; a_sign2 = 4'd15; a_sign3 = 4'd0;
b_sign0 = 4'd14; b_sign1 = 4'd1; b_sign2 = 4'd10; b_sign3 = 4'd5;
@(posedge clk_i);
a_mant0 = 8'd183; a_mant1 = 8'd122; a_mant2 = 8'd250; a_mant3 = 8'd185;
b_mant0 = 8'd35; b_mant1 = 8'd41; b_mant2 = 8'd202; b_mant3 = 8'd160;
a_exp0 = 10'd776; a_exp1 = 10'd751; a_exp2 = 10'd515; a_exp3 = 10'd680;
b_exp0 = 10'd857; b_exp1 = 10'd259; b_exp2 = 10'd760; b_exp3 = 10'd803;
a_sign0 = 4'd2; a_sign1 = 4'd9; a_sign2 = 4'd16; a_sign3 = 4'd6;
b_sign0 = 4'd12; b_sign1 = 4'd16; b_sign2 = 4'd8; b_sign3 = 4'd5;
@(posedge clk_i);
a_mant0 = 8'd115; a_mant1 = 8'd199; a_mant2 = 8'd239; a_mant3 = 8'd17;
b_mant0 = 8'd97; b_mant1 = 8'd48; b_mant2 = 8'd132; b_mant3 = 8'd255;
a_exp0 = 10'd1018; a_exp1 = 10'd572; a_exp2 = 10'd666; a_exp3 = 10'd458;
b_exp0 = 10'd921; b_exp1 = 10'd204; b_exp2 = 10'd892; b_exp3 = 10'd419;
a_sign0 = 4'd13; a_sign1 = 4'd0; a_sign2 = 4'd0; a_sign3 = 4'd8;
b_sign0 = 4'd3; b_sign1 = 4'd9; b_sign2 = 4'd10; b_sign3 = 4'd13;
@(posedge clk_i);
a_mant0 = 8'd215; a_mant1 = 8'd204; a_mant2 = 8'd142; a_mant3 = 8'd124;
b_mant0 = 8'd133; b_mant1 = 8'd167; b_mant2 = 8'd10; b_mant3 = 8'd95;
a_exp0 = 10'd158; a_exp1 = 10'd791; a_exp2 = 10'd1012; a_exp3 = 10'd325;
b_exp0 = 10'd791; b_exp1 = 10'd681; b_exp2 = 10'd932; b_exp3 = 10'd954;
a_sign0 = 4'd15; a_sign1 = 4'd8; a_sign2 = 4'd10; a_sign3 = 4'd4;
b_sign0 = 4'd2; b_sign1 = 4'd8; b_sign2 = 4'd16; b_sign3 = 4'd13;
@(posedge clk_i);
a_mant0 = 8'd83; a_mant1 = 8'd67; a_mant2 = 8'd135; a_mant3 = 8'd56;
b_mant0 = 8'd35; b_mant1 = 8'd112; b_mant2 = 8'd24; b_mant3 = 8'd70;
a_exp0 = 10'd691; a_exp1 = 10'd578; a_exp2 = 10'd276; a_exp3 = 10'd656;
b_exp0 = 10'd858; b_exp1 = 10'd993; b_exp2 = 10'd681; b_exp3 = 10'd33;
a_sign0 = 4'd5; a_sign1 = 4'd13; a_sign2 = 4'd13; a_sign3 = 4'd12;
b_sign0 = 4'd16; b_sign1 = 4'd15; b_sign2 = 4'd2; b_sign3 = 4'd12;
@(posedge clk_i);
shared_exps0 = 8'd142;
shared_exps1 = 8'd140;
a_mant0 = 8'd177; a_mant1 = 8'd156; a_mant2 = 8'd213; a_mant3 = 8'd249;
b_mant0 = 8'd101; b_mant1 = 8'd148; b_mant2 = 8'd144; b_mant3 = 8'd114;
a_exp0 = 10'd231; a_exp1 = 10'd967; a_exp2 = 10'd694; a_exp3 = 10'd148;
b_exp0 = 10'd1007; b_exp1 = 10'd326; b_exp2 = 10'd810; b_exp3 = 10'd109;
a_sign0 = 4'd12; a_sign1 = 4'd6; a_sign2 = 4'd10; a_sign3 = 4'd9;
b_sign0 = 4'd16; b_sign1 = 4'd12; b_sign2 = 4'd0; b_sign3 = 4'd2;
@(posedge clk_i);
a_mant0 = 8'd52; a_mant1 = 8'd36; a_mant2 = 8'd5; a_mant3 = 8'd111;
b_mant0 = 8'd147; b_mant1 = 8'd136; b_mant2 = 8'd180; b_mant3 = 8'd229;
a_exp0 = 10'd289; a_exp1 = 10'd842; a_exp2 = 10'd461; a_exp3 = 10'd249;
b_exp0 = 10'd271; b_exp1 = 10'd779; b_exp2 = 10'd316; b_exp3 = 10'd395;
a_sign0 = 4'd6; a_sign1 = 4'd16; a_sign2 = 4'd0; a_sign3 = 4'd16;
b_sign0 = 4'd15; b_sign1 = 4'd8; b_sign2 = 4'd5; b_sign3 = 4'd14;
@(posedge clk_i);
a_mant0 = 8'd29; a_mant1 = 8'd150; a_mant2 = 8'd91; a_mant3 = 8'd228;
b_mant0 = 8'd163; b_mant1 = 8'd102; b_mant2 = 8'd217; b_mant3 = 8'd88;
a_exp0 = 10'd258; a_exp1 = 10'd111; a_exp2 = 10'd296; a_exp3 = 10'd803;
b_exp0 = 10'd595; b_exp1 = 10'd361; b_exp2 = 10'd276; b_exp3 = 10'd997;
a_sign0 = 4'd12; a_sign1 = 4'd10; a_sign2 = 4'd6; a_sign3 = 4'd2;
b_sign0 = 4'd8; b_sign1 = 4'd14; b_sign2 = 4'd10; b_sign3 = 4'd5;
@(posedge clk_i);
a_mant0 = 8'd246; a_mant1 = 8'd115; a_mant2 = 8'd93; a_mant3 = 8'd153;
b_mant0 = 8'd183; b_mant1 = 8'd127; b_mant2 = 8'd213; b_mant3 = 8'd115;
a_exp0 = 10'd620; a_exp1 = 10'd739; a_exp2 = 10'd626; a_exp3 = 10'd48;
b_exp0 = 10'd556; b_exp1 = 10'd110; b_exp2 = 10'd836; b_exp3 = 10'd873;
a_sign0 = 4'd7; a_sign1 = 4'd6; a_sign2 = 4'd1; a_sign3 = 4'd2;
b_sign0 = 4'd13; b_sign1 = 4'd4; b_sign2 = 4'd9; b_sign3 = 4'd9;
@(posedge clk_i);
a_mant0 = 8'd175; a_mant1 = 8'd159; a_mant2 = 8'd228; a_mant3 = 8'd114;
b_mant0 = 8'd94; b_mant1 = 8'd169; b_mant2 = 8'd2; b_mant3 = 8'd231;
a_exp0 = 10'd562; a_exp1 = 10'd398; a_exp2 = 10'd174; a_exp3 = 10'd122;
b_exp0 = 10'd323; b_exp1 = 10'd231; b_exp2 = 10'd643; b_exp3 = 10'd331;
a_sign0 = 4'd10; a_sign1 = 4'd8; a_sign2 = 4'd14; a_sign3 = 4'd6;
b_sign0 = 4'd4; b_sign1 = 4'd6; b_sign2 = 4'd13; b_sign3 = 4'd6;
@(posedge clk_i);
a_mant0 = 8'd232; a_mant1 = 8'd187; a_mant2 = 8'd166; a_mant3 = 8'd187;
b_mant0 = 8'd42; b_mant1 = 8'd136; b_mant2 = 8'd254; b_mant3 = 8'd20;
a_exp0 = 10'd104; a_exp1 = 10'd32; a_exp2 = 10'd49; a_exp3 = 10'd35;
b_exp0 = 10'd231; b_exp1 = 10'd364; b_exp2 = 10'd135; b_exp3 = 10'd616;
a_sign0 = 4'd0; a_sign1 = 4'd0; a_sign2 = 4'd2; a_sign3 = 4'd3;
b_sign0 = 4'd12; b_sign1 = 4'd13; b_sign2 = 4'd3; b_sign3 = 4'd10;
@(posedge clk_i);
a_mant0 = 8'd80; a_mant1 = 8'd104; a_mant2 = 8'd54; a_mant3 = 8'd30;
b_mant0 = 8'd23; b_mant1 = 8'd11; b_mant2 = 8'd177; b_mant3 = 8'd244;
a_exp0 = 10'd535; a_exp1 = 10'd56; a_exp2 = 10'd110; a_exp3 = 10'd23;
b_exp0 = 10'd925; b_exp1 = 10'd960; b_exp2 = 10'd791; b_exp3 = 10'd212;
a_sign0 = 4'd3; a_sign1 = 4'd14; a_sign2 = 4'd5; a_sign3 = 4'd4;
b_sign0 = 4'd10; b_sign1 = 4'd0; b_sign2 = 4'd3; b_sign3 = 4'd11;
@(posedge clk_i);
a_mant0 = 8'd63; a_mant1 = 8'd126; a_mant2 = 8'd152; a_mant3 = 8'd175;
b_mant0 = 8'd81; b_mant1 = 8'd68; b_mant2 = 8'd56; b_mant3 = 8'd6;
a_exp0 = 10'd945; a_exp1 = 10'd871; a_exp2 = 10'd264; a_exp3 = 10'd1008;
b_exp0 = 10'd653; b_exp1 = 10'd379; b_exp2 = 10'd615; b_exp3 = 10'd116;
a_sign0 = 4'd13; a_sign1 = 4'd11; a_sign2 = 4'd8; a_sign3 = 4'd3;
b_sign0 = 4'd10; b_sign1 = 4'd14; b_sign2 = 4'd3; b_sign3 = 4'd10;
@(posedge clk_i);
shared_exps0 = 8'd152;
shared_exps1 = 8'd113;
a_mant0 = 8'd175; a_mant1 = 8'd42; a_mant2 = 8'd128; a_mant3 = 8'd216;
b_mant0 = 8'd44; b_mant1 = 8'd204; b_mant2 = 8'd158; b_mant3 = 8'd116;
a_exp0 = 10'd478; a_exp1 = 10'd471; a_exp2 = 10'd331; a_exp3 = 10'd561;
b_exp0 = 10'd950; b_exp1 = 10'd600; b_exp2 = 10'd736; b_exp3 = 10'd873;
a_sign0 = 4'd2; a_sign1 = 4'd7; a_sign2 = 4'd11; a_sign3 = 4'd13;
b_sign0 = 4'd10; b_sign1 = 4'd1; b_sign2 = 4'd15; b_sign3 = 4'd13;
@(posedge clk_i);
a_mant0 = 8'd49; a_mant1 = 8'd245; a_mant2 = 8'd78; a_mant3 = 8'd10;
b_mant0 = 8'd140; b_mant1 = 8'd85; b_mant2 = 8'd158; b_mant3 = 8'd86;
a_exp0 = 10'd394; a_exp1 = 10'd882; a_exp2 = 10'd248; a_exp3 = 10'd1008;
b_exp0 = 10'd739; b_exp1 = 10'd172; b_exp2 = 10'd911; b_exp3 = 10'd763;
a_sign0 = 4'd3; a_sign1 = 4'd1; a_sign2 = 4'd11; a_sign3 = 4'd13;
b_sign0 = 4'd14; b_sign1 = 4'd7; b_sign2 = 4'd14; b_sign3 = 4'd10;
@(posedge clk_i);
a_mant0 = 8'd26; a_mant1 = 8'd66; a_mant2 = 8'd81; a_mant3 = 8'd34;
b_mant0 = 8'd168; b_mant1 = 8'd129; b_mant2 = 8'd59; b_mant3 = 8'd12;
a_exp0 = 10'd261; a_exp1 = 10'd271; a_exp2 = 10'd337; a_exp3 = 10'd945;
b_exp0 = 10'd249; b_exp1 = 10'd603; b_exp2 = 10'd263; b_exp3 = 10'd896;
a_sign0 = 4'd0; a_sign1 = 4'd0; a_sign2 = 4'd1; a_sign3 = 4'd6;
b_sign0 = 4'd16; b_sign1 = 4'd1; b_sign2 = 4'd3; b_sign3 = 4'd11;
@(posedge clk_i);
a_mant0 = 8'd226; a_mant1 = 8'd121; a_mant2 = 8'd138; a_mant3 = 8'd186;
b_mant0 = 8'd171; b_mant1 = 8'd201; b_mant2 = 8'd145; b_mant3 = 8'd176;
a_exp0 = 10'd318; a_exp1 = 10'd362; a_exp2 = 10'd336; a_exp3 = 10'd147;
b_exp0 = 10'd264; b_exp1 = 10'd801; b_exp2 = 10'd82; b_exp3 = 10'd605;
a_sign0 = 4'd0; a_sign1 = 4'd1; a_sign2 = 4'd4; a_sign3 = 4'd7;
b_sign0 = 4'd16; b_sign1 = 4'd7; b_sign2 = 4'd5; b_sign3 = 4'd11;
@(posedge clk_i);
a_mant0 = 8'd143; a_mant1 = 8'd175; a_mant2 = 8'd81; a_mant3 = 8'd149;
b_mant0 = 8'd24; b_mant1 = 8'd238; b_mant2 = 8'd143; b_mant3 = 8'd79;
a_exp0 = 10'd394; a_exp1 = 10'd289; a_exp2 = 10'd244; a_exp3 = 10'd188;
b_exp0 = 10'd690; b_exp1 = 10'd521; b_exp2 = 10'd254; b_exp3 = 10'd791;
a_sign0 = 4'd9; a_sign1 = 4'd5; a_sign2 = 4'd0; a_sign3 = 4'd2;
b_sign0 = 4'd2; b_sign1 = 4'd12; b_sign2 = 4'd6; b_sign3 = 4'd1;
@(posedge clk_i);
a_mant0 = 8'd117; a_mant1 = 8'd207; a_mant2 = 8'd240; a_mant3 = 8'd85;
b_mant0 = 8'd20; b_mant1 = 8'd36; b_mant2 = 8'd149; b_mant3 = 8'd230;
a_exp0 = 10'd283; a_exp1 = 10'd678; a_exp2 = 10'd133; a_exp3 = 10'd8;
b_exp0 = 10'd276; b_exp1 = 10'd34; b_exp2 = 10'd588; b_exp3 = 10'd893;
a_sign0 = 4'd15; a_sign1 = 4'd4; a_sign2 = 4'd13; a_sign3 = 4'd10;
b_sign0 = 4'd7; b_sign1 = 4'd0; b_sign2 = 4'd9; b_sign3 = 4'd7;
@(posedge clk_i);
a_mant0 = 8'd107; a_mant1 = 8'd147; a_mant2 = 8'd82; a_mant3 = 8'd32;
b_mant0 = 8'd35; b_mant1 = 8'd34; b_mant2 = 8'd182; b_mant3 = 8'd214;
a_exp0 = 10'd1003; a_exp1 = 10'd822; a_exp2 = 10'd662; a_exp3 = 10'd421;
b_exp0 = 10'd94; b_exp1 = 10'd594; b_exp2 = 10'd857; b_exp3 = 10'd135;
a_sign0 = 4'd5; a_sign1 = 4'd8; a_sign2 = 4'd0; a_sign3 = 4'd9;
b_sign0 = 4'd7; b_sign1 = 4'd15; b_sign2 = 4'd1; b_sign3 = 4'd7;
@(posedge clk_i);
a_mant0 = 8'd244; a_mant1 = 8'd162; a_mant2 = 8'd129; a_mant3 = 8'd61;
b_mant0 = 8'd232; b_mant1 = 8'd206; b_mant2 = 8'd193; b_mant3 = 8'd225;
a_exp0 = 10'd581; a_exp1 = 10'd655; a_exp2 = 10'd446; a_exp3 = 10'd575;
b_exp0 = 10'd29; b_exp1 = 10'd113; b_exp2 = 10'd46; b_exp3 = 10'd628;
a_sign0 = 4'd2; a_sign1 = 4'd14; a_sign2 = 4'd13; a_sign3 = 4'd15;
b_sign0 = 4'd5; b_sign1 = 4'd10; b_sign2 = 4'd16; b_sign3 = 4'd15;
@(posedge clk_i);
shared_exps0 = 8'd170;
shared_exps1 = 8'd140;
rstn = 0;
@(posedge clk_i);
rstn = 1;
a_mant0 = 8'd45; a_mant1 = 8'd35; a_mant2 = 8'd144; a_mant3 = 8'd157;
b_mant0 = 8'd189; b_mant1 = 8'd214; b_mant2 = 8'd143; b_mant3 = 8'd143;
a_exp0 = 10'd553; a_exp1 = 10'd409; a_exp2 = 10'd529; a_exp3 = 10'd655;
b_exp0 = 10'd1016; b_exp1 = 10'd122; b_exp2 = 10'd379; b_exp3 = 10'd522;
a_sign0 = 4'd0; a_sign1 = 4'd9; a_sign2 = 4'd11; a_sign3 = 4'd8;
b_sign0 = 4'd16; b_sign1 = 4'd7; b_sign2 = 4'd14; b_sign3 = 4'd3;
@(posedge clk_i);
a_mant0 = 8'd222; a_mant1 = 8'd173; a_mant2 = 8'd95; a_mant3 = 8'd155;
b_mant0 = 8'd150; b_mant1 = 8'd86; b_mant2 = 8'd12; b_mant3 = 8'd89;
a_exp0 = 10'd96; a_exp1 = 10'd586; a_exp2 = 10'd858; a_exp3 = 10'd9;
b_exp0 = 10'd824; b_exp1 = 10'd279; b_exp2 = 10'd831; b_exp3 = 10'd345;
a_sign0 = 4'd6; a_sign1 = 4'd7; a_sign2 = 4'd8; a_sign3 = 4'd3;
b_sign0 = 4'd16; b_sign1 = 4'd14; b_sign2 = 4'd5; b_sign3 = 4'd4;
@(posedge clk_i);
a_mant0 = 8'd191; a_mant1 = 8'd12; a_mant2 = 8'd222; a_mant3 = 8'd51;
b_mant0 = 8'd152; b_mant1 = 8'd28; b_mant2 = 8'd184; b_mant3 = 8'd135;
a_exp0 = 10'd366; a_exp1 = 10'd965; a_exp2 = 10'd303; a_exp3 = 10'd370;
b_exp0 = 10'd888; b_exp1 = 10'd9; b_exp2 = 10'd760; b_exp3 = 10'd216;
a_sign0 = 4'd12; a_sign1 = 4'd1; a_sign2 = 4'd9; a_sign3 = 4'd15;
b_sign0 = 4'd14; b_sign1 = 4'd12; b_sign2 = 4'd0; b_sign3 = 4'd0;
@(posedge clk_i);
a_mant0 = 8'd85; a_mant1 = 8'd169; a_mant2 = 8'd201; a_mant3 = 8'd199;
b_mant0 = 8'd107; b_mant1 = 8'd109; b_mant2 = 8'd184; b_mant3 = 8'd68;
a_exp0 = 10'd803; a_exp1 = 10'd301; a_exp2 = 10'd456; a_exp3 = 10'd552;
b_exp0 = 10'd256; b_exp1 = 10'd299; b_exp2 = 10'd633; b_exp3 = 10'd432;
a_sign0 = 4'd12; a_sign1 = 4'd16; a_sign2 = 4'd13; a_sign3 = 4'd3;
b_sign0 = 4'd14; b_sign1 = 4'd3; b_sign2 = 4'd10; b_sign3 = 4'd11;
@(posedge clk_i);
a_mant0 = 8'd216; a_mant1 = 8'd80; a_mant2 = 8'd69; a_mant3 = 8'd100;
b_mant0 = 8'd198; b_mant1 = 8'd64; b_mant2 = 8'd85; b_mant3 = 8'd66;
a_exp0 = 10'd475; a_exp1 = 10'd648; a_exp2 = 10'd440; a_exp3 = 10'd72;
b_exp0 = 10'd686; b_exp1 = 10'd867; b_exp2 = 10'd882; b_exp3 = 10'd931;
a_sign0 = 4'd4; a_sign1 = 4'd3; a_sign2 = 4'd2; a_sign3 = 4'd10;
b_sign0 = 4'd1; b_sign1 = 4'd9; b_sign2 = 4'd6; b_sign3 = 4'd9;
@(posedge clk_i);
a_mant0 = 8'd121; a_mant1 = 8'd75; a_mant2 = 8'd68; a_mant3 = 8'd43;
b_mant0 = 8'd216; b_mant1 = 8'd23; b_mant2 = 8'd0; b_mant3 = 8'd202;
a_exp0 = 10'd608; a_exp1 = 10'd878; a_exp2 = 10'd854; a_exp3 = 10'd820;
b_exp0 = 10'd56; b_exp1 = 10'd857; b_exp2 = 10'd120; b_exp3 = 10'd659;
a_sign0 = 4'd4; a_sign1 = 4'd0; a_sign2 = 4'd4; a_sign3 = 4'd12;
b_sign0 = 4'd3; b_sign1 = 4'd14; b_sign2 = 4'd10; b_sign3 = 4'd7;
@(posedge clk_i);
a_mant0 = 8'd37; a_mant1 = 8'd171; a_mant2 = 8'd245; a_mant3 = 8'd104;
b_mant0 = 8'd225; b_mant1 = 8'd30; b_mant2 = 8'd72; b_mant3 = 8'd1;
a_exp0 = 10'd580; a_exp1 = 10'd217; a_exp2 = 10'd854; a_exp3 = 10'd919;
b_exp0 = 10'd841; b_exp1 = 10'd862; b_exp2 = 10'd739; b_exp3 = 10'd785;
a_sign0 = 4'd3; a_sign1 = 4'd9; a_sign2 = 4'd15; a_sign3 = 4'd8;
b_sign0 = 4'd11; b_sign1 = 4'd2; b_sign2 = 4'd4; b_sign3 = 4'd14;
@(posedge clk_i);
shared_exps0 = 8'd115;
shared_exps1 = 8'd82;
a_mant0 = 8'd243; a_mant1 = 8'd21; a_mant2 = 8'd136; a_mant3 = 8'd92;
b_mant0 = 8'd158; b_mant1 = 8'd12; b_mant2 = 8'd217; b_mant3 = 8'd78;
a_exp0 = 10'd370; a_exp1 = 10'd735; a_exp2 = 10'd742; a_exp3 = 10'd769;
b_exp0 = 10'd18; b_exp1 = 10'd940; b_exp2 = 10'd699; b_exp3 = 10'd450;
a_sign0 = 4'd5; a_sign1 = 4'd13; a_sign2 = 4'd5; a_sign3 = 4'd10;
b_sign0 = 4'd9; b_sign1 = 4'd12; b_sign2 = 4'd2; b_sign3 = 4'd10;
@(posedge clk_i);
a_mant0 = 8'd43; a_mant1 = 8'd148; a_mant2 = 8'd50; a_mant3 = 8'd156;
b_mant0 = 8'd214; b_mant1 = 8'd59; b_mant2 = 8'd130; b_mant3 = 8'd152;
a_exp0 = 10'd186; a_exp1 = 10'd381; a_exp2 = 10'd115; a_exp3 = 10'd898;
b_exp0 = 10'd940; b_exp1 = 10'd428; b_exp2 = 10'd944; b_exp3 = 10'd539;
a_sign0 = 4'd2; a_sign1 = 4'd4; a_sign2 = 4'd5; a_sign3 = 4'd5;
b_sign0 = 4'd5; b_sign1 = 4'd7; b_sign2 = 4'd6; b_sign3 = 4'd4;
@(posedge clk_i);
a_mant0 = 8'd196; a_mant1 = 8'd18; a_mant2 = 8'd141; a_mant3 = 8'd25;
b_mant0 = 8'd94; b_mant1 = 8'd229; b_mant2 = 8'd88; b_mant3 = 8'd48;
a_exp0 = 10'd33; a_exp1 = 10'd613; a_exp2 = 10'd573; a_exp3 = 10'd590;
b_exp0 = 10'd482; b_exp1 = 10'd662; b_exp2 = 10'd292; b_exp3 = 10'd94;
a_sign0 = 4'd4; a_sign1 = 4'd12; a_sign2 = 4'd10; a_sign3 = 4'd8;
b_sign0 = 4'd0; b_sign1 = 4'd13; b_sign2 = 4'd6; b_sign3 = 4'd0;
@(posedge clk_i);
a_mant0 = 8'd63; a_mant1 = 8'd75; a_mant2 = 8'd127; a_mant3 = 8'd3;
b_mant0 = 8'd56; b_mant1 = 8'd252; b_mant2 = 8'd203; b_mant3 = 8'd209;
a_exp0 = 10'd437; a_exp1 = 10'd155; a_exp2 = 10'd91; a_exp3 = 10'd399;
b_exp0 = 10'd303; b_exp1 = 10'd865; b_exp2 = 10'd79; b_exp3 = 10'd342;
a_sign0 = 4'd0; a_sign1 = 4'd15; a_sign2 = 4'd2; a_sign3 = 4'd4;
b_sign0 = 4'd12; b_sign1 = 4'd5; b_sign2 = 4'd2; b_sign3 = 4'd3;
@(posedge clk_i);
a_mant0 = 8'd179; a_mant1 = 8'd66; a_mant2 = 8'd137; a_mant3 = 8'd232;
b_mant0 = 8'd117; b_mant1 = 8'd214; b_mant2 = 8'd162; b_mant3 = 8'd146;
a_exp0 = 10'd304; a_exp1 = 10'd899; a_exp2 = 10'd999; a_exp3 = 10'd791;
b_exp0 = 10'd24; b_exp1 = 10'd987; b_exp2 = 10'd714; b_exp3 = 10'd306;
a_sign0 = 4'd7; a_sign1 = 4'd12; a_sign2 = 4'd1; a_sign3 = 4'd9;
b_sign0 = 4'd16; b_sign1 = 4'd2; b_sign2 = 4'd11; b_sign3 = 4'd1;
@(posedge clk_i);
a_mant0 = 8'd129; a_mant1 = 8'd46; a_mant2 = 8'd50; a_mant3 = 8'd132;
b_mant0 = 8'd156; b_mant1 = 8'd204; b_mant2 = 8'd6; b_mant3 = 8'd89;
a_exp0 = 10'd420; a_exp1 = 10'd43; a_exp2 = 10'd199; a_exp3 = 10'd5;
b_exp0 = 10'd1002; b_exp1 = 10'd340; b_exp2 = 10'd121; b_exp3 = 10'd425;
a_sign0 = 4'd8; a_sign1 = 4'd6; a_sign2 = 4'd2; a_sign3 = 4'd2;
b_sign0 = 4'd8; b_sign1 = 4'd9; b_sign2 = 4'd13; b_sign3 = 4'd16;
@(posedge clk_i);
a_mant0 = 8'd253; a_mant1 = 8'd38; a_mant2 = 8'd74; a_mant3 = 8'd12;
b_mant0 = 8'd210; b_mant1 = 8'd104; b_mant2 = 8'd54; b_mant3 = 8'd248;
a_exp0 = 10'd167; a_exp1 = 10'd634; a_exp2 = 10'd412; a_exp3 = 10'd444;
b_exp0 = 10'd928; b_exp1 = 10'd541; b_exp2 = 10'd996; b_exp3 = 10'd283;
a_sign0 = 4'd13; a_sign1 = 4'd13; a_sign2 = 4'd1; a_sign3 = 4'd10;
b_sign0 = 4'd15; b_sign1 = 4'd14; b_sign2 = 4'd15; b_sign3 = 4'd13;
@(posedge clk_i);
a_mant0 = 8'd204; a_mant1 = 8'd185; a_mant2 = 8'd21; a_mant3 = 8'd171;
b_mant0 = 8'd172; b_mant1 = 8'd41; b_mant2 = 8'd248; b_mant3 = 8'd28;
a_exp0 = 10'd114; a_exp1 = 10'd123; a_exp2 = 10'd550; a_exp3 = 10'd447;
b_exp0 = 10'd791; b_exp1 = 10'd706; b_exp2 = 10'd795; b_exp3 = 10'd333;
a_sign0 = 4'd1; a_sign1 = 4'd2; a_sign2 = 4'd15; a_sign3 = 4'd10;
b_sign0 = 4'd5; b_sign1 = 4'd11; b_sign2 = 4'd2; b_sign3 = 4'd14;
@(posedge clk_i);
shared_exps0 = 8'd110;
shared_exps1 = 8'd140;
a_mant0 = 8'd144; a_mant1 = 8'd116; a_mant2 = 8'd103; a_mant3 = 8'd167;
b_mant0 = 8'd8; b_mant1 = 8'd163; b_mant2 = 8'd58; b_mant3 = 8'd200;
a_exp0 = 10'd904; a_exp1 = 10'd111; a_exp2 = 10'd739; a_exp3 = 10'd31;
b_exp0 = 10'd39; b_exp1 = 10'd490; b_exp2 = 10'd421; b_exp3 = 10'd85;
a_sign0 = 4'd4; a_sign1 = 4'd3; a_sign2 = 4'd16; a_sign3 = 4'd12;
b_sign0 = 4'd5; b_sign1 = 4'd15; b_sign2 = 4'd9; b_sign3 = 4'd3;
@(posedge clk_i);
a_mant0 = 8'd28; a_mant1 = 8'd119; a_mant2 = 8'd246; a_mant3 = 8'd205;
b_mant0 = 8'd213; b_mant1 = 8'd28; b_mant2 = 8'd50; b_mant3 = 8'd63;
a_exp0 = 10'd321; a_exp1 = 10'd873; a_exp2 = 10'd516; a_exp3 = 10'd149;
b_exp0 = 10'd73; b_exp1 = 10'd492; b_exp2 = 10'd476; b_exp3 = 10'd458;
a_sign0 = 4'd16; a_sign1 = 4'd5; a_sign2 = 4'd16; a_sign3 = 4'd9;
b_sign0 = 4'd13; b_sign1 = 4'd8; b_sign2 = 4'd13; b_sign3 = 4'd16;
@(posedge clk_i);
a_mant0 = 8'd59; a_mant1 = 8'd63; a_mant2 = 8'd129; a_mant3 = 8'd206;
b_mant0 = 8'd189; b_mant1 = 8'd150; b_mant2 = 8'd145; b_mant3 = 8'd196;
a_exp0 = 10'd94; a_exp1 = 10'd788; a_exp2 = 10'd893; a_exp3 = 10'd1012;
b_exp0 = 10'd295; b_exp1 = 10'd544; b_exp2 = 10'd567; b_exp3 = 10'd629;
a_sign0 = 4'd3; a_sign1 = 4'd1; a_sign2 = 4'd6; a_sign3 = 4'd15;
b_sign0 = 4'd10; b_sign1 = 4'd15; b_sign2 = 4'd10; b_sign3 = 4'd4;
@(posedge clk_i);
a_mant0 = 8'd6; a_mant1 = 8'd80; a_mant2 = 8'd66; a_mant3 = 8'd27;
b_mant0 = 8'd168; b_mant1 = 8'd136; b_mant2 = 8'd158; b_mant3 = 8'd162;
a_exp0 = 10'd680; a_exp1 = 10'd784; a_exp2 = 10'd188; a_exp3 = 10'd575;
b_exp0 = 10'd376; b_exp1 = 10'd80; b_exp2 = 10'd980; b_exp3 = 10'd155;
a_sign0 = 4'd7; a_sign1 = 4'd13; a_sign2 = 4'd12; a_sign3 = 4'd2;
b_sign0 = 4'd8; b_sign1 = 4'd6; b_sign2 = 4'd9; b_sign3 = 4'd9;
@(posedge clk_i);
a_mant0 = 8'd87; a_mant1 = 8'd214; a_mant2 = 8'd131; a_mant3 = 8'd83;
b_mant0 = 8'd194; b_mant1 = 8'd34; b_mant2 = 8'd20; b_mant3 = 8'd117;
a_exp0 = 10'd706; a_exp1 = 10'd302; a_exp2 = 10'd246; a_exp3 = 10'd639;
b_exp0 = 10'd195; b_exp1 = 10'd500; b_exp2 = 10'd520; b_exp3 = 10'd214;
a_sign0 = 4'd0; a_sign1 = 4'd7; a_sign2 = 4'd12; a_sign3 = 4'd13;
b_sign0 = 4'd1; b_sign1 = 4'd16; b_sign2 = 4'd9; b_sign3 = 4'd10;
@(posedge clk_i);
a_mant0 = 8'd245; a_mant1 = 8'd180; a_mant2 = 8'd35; a_mant3 = 8'd80;
b_mant0 = 8'd167; b_mant1 = 8'd32; b_mant2 = 8'd96; b_mant3 = 8'd201;
a_exp0 = 10'd951; a_exp1 = 10'd807; a_exp2 = 10'd259; a_exp3 = 10'd167;
b_exp0 = 10'd456; b_exp1 = 10'd346; b_exp2 = 10'd603; b_exp3 = 10'd124;
a_sign0 = 4'd1; a_sign1 = 4'd9; a_sign2 = 4'd0; a_sign3 = 4'd16;
b_sign0 = 4'd2; b_sign1 = 4'd15; b_sign2 = 4'd4; b_sign3 = 4'd10;
@(posedge clk_i);
a_mant0 = 8'd169; a_mant1 = 8'd100; a_mant2 = 8'd93; a_mant3 = 8'd206;
b_mant0 = 8'd33; b_mant1 = 8'd128; b_mant2 = 8'd124; b_mant3 = 8'd119;
a_exp0 = 10'd420; a_exp1 = 10'd578; a_exp2 = 10'd85; a_exp3 = 10'd135;
b_exp0 = 10'd123; b_exp1 = 10'd641; b_exp2 = 10'd1000; b_exp3 = 10'd295;
a_sign0 = 4'd9; a_sign1 = 4'd1; a_sign2 = 4'd3; a_sign3 = 4'd9;
b_sign0 = 4'd10; b_sign1 = 4'd4; b_sign2 = 4'd10; b_sign3 = 4'd11;
@(posedge clk_i);
a_mant0 = 8'd79; a_mant1 = 8'd19; a_mant2 = 8'd177; a_mant3 = 8'd120;
b_mant0 = 8'd240; b_mant1 = 8'd231; b_mant2 = 8'd135; b_mant3 = 8'd215;
a_exp0 = 10'd424; a_exp1 = 10'd303; a_exp2 = 10'd912; a_exp3 = 10'd941;
b_exp0 = 10'd795; b_exp1 = 10'd205; b_exp2 = 10'd479; b_exp3 = 10'd922;
a_sign0 = 4'd1; a_sign1 = 4'd8; a_sign2 = 4'd9; a_sign3 = 4'd9;
b_sign0 = 4'd6; b_sign1 = 4'd6; b_sign2 = 4'd0; b_sign3 = 4'd7;
@(posedge clk_i);
shared_exps0 = 8'd142;
shared_exps1 = 8'd96;
a_mant0 = 8'd250; a_mant1 = 8'd231; a_mant2 = 8'd113; a_mant3 = 8'd59;
b_mant0 = 8'd191; b_mant1 = 8'd221; b_mant2 = 8'd34; b_mant3 = 8'd90;
a_exp0 = 10'd163; a_exp1 = 10'd758; a_exp2 = 10'd442; a_exp3 = 10'd888;
b_exp0 = 10'd420; b_exp1 = 10'd679; b_exp2 = 10'd584; b_exp3 = 10'd196;
a_sign0 = 4'd6; a_sign1 = 4'd0; a_sign2 = 4'd0; a_sign3 = 4'd1;
b_sign0 = 4'd1; b_sign1 = 4'd13; b_sign2 = 4'd16; b_sign3 = 4'd9;
@(posedge clk_i);
a_mant0 = 8'd2; a_mant1 = 8'd7; a_mant2 = 8'd95; a_mant3 = 8'd252;
b_mant0 = 8'd169; b_mant1 = 8'd187; b_mant2 = 8'd162; b_mant3 = 8'd186;
a_exp0 = 10'd284; a_exp1 = 10'd783; a_exp2 = 10'd968; a_exp3 = 10'd335;
b_exp0 = 10'd688; b_exp1 = 10'd755; b_exp2 = 10'd956; b_exp3 = 10'd878;
a_sign0 = 4'd0; a_sign1 = 4'd15; a_sign2 = 4'd4; a_sign3 = 4'd4;
b_sign0 = 4'd10; b_sign1 = 4'd0; b_sign2 = 4'd12; b_sign3 = 4'd14;
@(posedge clk_i);
a_mant0 = 8'd172; a_mant1 = 8'd181; a_mant2 = 8'd52; a_mant3 = 8'd118;
b_mant0 = 8'd132; b_mant1 = 8'd179; b_mant2 = 8'd199; b_mant3 = 8'd111;
a_exp0 = 10'd941; a_exp1 = 10'd386; a_exp2 = 10'd842; a_exp3 = 10'd452;
b_exp0 = 10'd754; b_exp1 = 10'd341; b_exp2 = 10'd915; b_exp3 = 10'd763;
a_sign0 = 4'd8; a_sign1 = 4'd12; a_sign2 = 4'd13; a_sign3 = 4'd7;
b_sign0 = 4'd7; b_sign1 = 4'd10; b_sign2 = 4'd11; b_sign3 = 4'd6;
@(posedge clk_i);
a_mant0 = 8'd125; a_mant1 = 8'd217; a_mant2 = 8'd0; a_mant3 = 8'd74;
b_mant0 = 8'd96; b_mant1 = 8'd236; b_mant2 = 8'd14; b_mant3 = 8'd244;
a_exp0 = 10'd264; a_exp1 = 10'd913; a_exp2 = 10'd303; a_exp3 = 10'd758;
b_exp0 = 10'd362; b_exp1 = 10'd357; b_exp2 = 10'd41; b_exp3 = 10'd392;
a_sign0 = 4'd10; a_sign1 = 4'd10; a_sign2 = 4'd12; a_sign3 = 4'd4;
b_sign0 = 4'd6; b_sign1 = 4'd9; b_sign2 = 4'd12; b_sign3 = 4'd16;
@(posedge clk_i);
a_mant0 = 8'd32; a_mant1 = 8'd199; a_mant2 = 8'd104; a_mant3 = 8'd231;
b_mant0 = 8'd216; b_mant1 = 8'd74; b_mant2 = 8'd159; b_mant3 = 8'd238;
a_exp0 = 10'd390; a_exp1 = 10'd741; a_exp2 = 10'd695; a_exp3 = 10'd785;
b_exp0 = 10'd677; b_exp1 = 10'd34; b_exp2 = 10'd261; b_exp3 = 10'd440;
a_sign0 = 4'd6; a_sign1 = 4'd1; a_sign2 = 4'd7; a_sign3 = 4'd7;
b_sign0 = 4'd4; b_sign1 = 4'd0; b_sign2 = 4'd7; b_sign3 = 4'd10;
@(posedge clk_i);
a_mant0 = 8'd108; a_mant1 = 8'd227; a_mant2 = 8'd233; a_mant3 = 8'd99;
b_mant0 = 8'd5; b_mant1 = 8'd92; b_mant2 = 8'd126; b_mant3 = 8'd207;
a_exp0 = 10'd928; a_exp1 = 10'd960; a_exp2 = 10'd271; a_exp3 = 10'd664;
b_exp0 = 10'd184; b_exp1 = 10'd25; b_exp2 = 10'd52; b_exp3 = 10'd962;
a_sign0 = 4'd1; a_sign1 = 4'd10; a_sign2 = 4'd10; a_sign3 = 4'd9;
b_sign0 = 4'd8; b_sign1 = 4'd14; b_sign2 = 4'd11; b_sign3 = 4'd2;
@(posedge clk_i);
a_mant0 = 8'd44; a_mant1 = 8'd224; a_mant2 = 8'd211; a_mant3 = 8'd99;
b_mant0 = 8'd117; b_mant1 = 8'd205; b_mant2 = 8'd65; b_mant3 = 8'd211;
a_exp0 = 10'd363; a_exp1 = 10'd487; a_exp2 = 10'd252; a_exp3 = 10'd791;
b_exp0 = 10'd205; b_exp1 = 10'd233; b_exp2 = 10'd918; b_exp3 = 10'd306;
a_sign0 = 4'd10; a_sign1 = 4'd11; a_sign2 = 4'd9; a_sign3 = 4'd16;
b_sign0 = 4'd14; b_sign1 = 4'd6; b_sign2 = 4'd6; b_sign3 = 4'd7;
@(posedge clk_i);
a_mant0 = 8'd235; a_mant1 = 8'd150; a_mant2 = 8'd223; a_mant3 = 8'd188;
b_mant0 = 8'd170; b_mant1 = 8'd21; b_mant2 = 8'd12; b_mant3 = 8'd45;
a_exp0 = 10'd884; a_exp1 = 10'd273; a_exp2 = 10'd51; a_exp3 = 10'd955;
b_exp0 = 10'd718; b_exp1 = 10'd657; b_exp2 = 10'd339; b_exp3 = 10'd637;
a_sign0 = 4'd15; a_sign1 = 4'd10; a_sign2 = 4'd6; a_sign3 = 4'd9;
b_sign0 = 4'd10; b_sign1 = 4'd9; b_sign2 = 4'd14; b_sign3 = 4'd13;
@(posedge clk_i);
shared_exps0 = 8'd137;
shared_exps1 = 8'd115;
rstn = 0;
@(posedge clk_i);
rstn = 1;
a_mant0 = 8'd178; a_mant1 = 8'd224; a_mant2 = 8'd223; a_mant3 = 8'd21;
b_mant0 = 8'd193; b_mant1 = 8'd26; b_mant2 = 8'd160; b_mant3 = 8'd208;
a_exp0 = 10'd784; a_exp1 = 10'd703; a_exp2 = 10'd80; a_exp3 = 10'd994;
b_exp0 = 10'd21; b_exp1 = 10'd473; b_exp2 = 10'd403; b_exp3 = 10'd298;
a_sign0 = 4'd4; a_sign1 = 4'd0; a_sign2 = 4'd6; a_sign3 = 4'd1;
b_sign0 = 4'd10; b_sign1 = 4'd3; b_sign2 = 4'd14; b_sign3 = 4'd16;
@(posedge clk_i);
a_mant0 = 8'd60; a_mant1 = 8'd233; a_mant2 = 8'd6; a_mant3 = 8'd127;
b_mant0 = 8'd96; b_mant1 = 8'd48; b_mant2 = 8'd68; b_mant3 = 8'd102;
a_exp0 = 10'd301; a_exp1 = 10'd128; a_exp2 = 10'd618; a_exp3 = 10'd408;
b_exp0 = 10'd274; b_exp1 = 10'd342; b_exp2 = 10'd549; b_exp3 = 10'd946;
a_sign0 = 4'd9; a_sign1 = 4'd12; a_sign2 = 4'd3; a_sign3 = 4'd10;
b_sign0 = 4'd11; b_sign1 = 4'd1; b_sign2 = 4'd3; b_sign3 = 4'd14;
@(posedge clk_i);
a_mant0 = 8'd147; a_mant1 = 8'd173; a_mant2 = 8'd5; a_mant3 = 8'd143;
b_mant0 = 8'd191; b_mant1 = 8'd0; b_mant2 = 8'd92; b_mant3 = 8'd10;
a_exp0 = 10'd704; a_exp1 = 10'd694; a_exp2 = 10'd81; a_exp3 = 10'd292;
b_exp0 = 10'd730; b_exp1 = 10'd158; b_exp2 = 10'd245; b_exp3 = 10'd16;
a_sign0 = 4'd12; a_sign1 = 4'd6; a_sign2 = 4'd16; a_sign3 = 4'd1;
b_sign0 = 4'd16; b_sign1 = 4'd14; b_sign2 = 4'd2; b_sign3 = 4'd10;
@(posedge clk_i);
a_mant0 = 8'd160; a_mant1 = 8'd201; a_mant2 = 8'd220; a_mant3 = 8'd145;
b_mant0 = 8'd114; b_mant1 = 8'd99; b_mant2 = 8'd29; b_mant3 = 8'd168;
a_exp0 = 10'd611; a_exp1 = 10'd601; a_exp2 = 10'd516; a_exp3 = 10'd675;
b_exp0 = 10'd942; b_exp1 = 10'd376; b_exp2 = 10'd314; b_exp3 = 10'd325;
a_sign0 = 4'd4; a_sign1 = 4'd4; a_sign2 = 4'd4; a_sign3 = 4'd10;
b_sign0 = 4'd16; b_sign1 = 4'd16; b_sign2 = 4'd1; b_sign3 = 4'd4;
@(posedge clk_i);
a_mant0 = 8'd154; a_mant1 = 8'd214; a_mant2 = 8'd237; a_mant3 = 8'd6;
b_mant0 = 8'd199; b_mant1 = 8'd116; b_mant2 = 8'd14; b_mant3 = 8'd147;
a_exp0 = 10'd280; a_exp1 = 10'd132; a_exp2 = 10'd296; a_exp3 = 10'd788;
b_exp0 = 10'd327; b_exp1 = 10'd866; b_exp2 = 10'd11; b_exp3 = 10'd800;
a_sign0 = 4'd16; a_sign1 = 4'd2; a_sign2 = 4'd4; a_sign3 = 4'd11;
b_sign0 = 4'd6; b_sign1 = 4'd12; b_sign2 = 4'd5; b_sign3 = 4'd12;
@(posedge clk_i);
a_mant0 = 8'd37; a_mant1 = 8'd162; a_mant2 = 8'd181; a_mant3 = 8'd101;
b_mant0 = 8'd4; b_mant1 = 8'd230; b_mant2 = 8'd171; b_mant3 = 8'd225;
a_exp0 = 10'd659; a_exp1 = 10'd323; a_exp2 = 10'd162; a_exp3 = 10'd512;
b_exp0 = 10'd636; b_exp1 = 10'd196; b_exp2 = 10'd866; b_exp3 = 10'd618;
a_sign0 = 4'd6; a_sign1 = 4'd7; a_sign2 = 4'd6; a_sign3 = 4'd0;
b_sign0 = 4'd8; b_sign1 = 4'd9; b_sign2 = 4'd13; b_sign3 = 4'd13;
@(posedge clk_i);
a_mant0 = 8'd9; a_mant1 = 8'd144; a_mant2 = 8'd41; a_mant3 = 8'd137;
b_mant0 = 8'd17; b_mant1 = 8'd24; b_mant2 = 8'd2; b_mant3 = 8'd174;
a_exp0 = 10'd802; a_exp1 = 10'd200; a_exp2 = 10'd59; a_exp3 = 10'd993;
b_exp0 = 10'd822; b_exp1 = 10'd101; b_exp2 = 10'd926; b_exp3 = 10'd420;
a_sign0 = 4'd4; a_sign1 = 4'd11; a_sign2 = 4'd16; a_sign3 = 4'd6;
b_sign0 = 4'd5; b_sign1 = 4'd3; b_sign2 = 4'd8; b_sign3 = 4'd1;
@(posedge clk_i);
shared_exps0 = 8'd146;
shared_exps1 = 8'd127;
a_mant0 = 8'd53; a_mant1 = 8'd81; a_mant2 = 8'd88; a_mant3 = 8'd217;
b_mant0 = 8'd34; b_mant1 = 8'd55; b_mant2 = 8'd131; b_mant3 = 8'd106;
a_exp0 = 10'd131; a_exp1 = 10'd783; a_exp2 = 10'd209; a_exp3 = 10'd575;
b_exp0 = 10'd549; b_exp1 = 10'd592; b_exp2 = 10'd655; b_exp3 = 10'd250;
a_sign0 = 4'd10; a_sign1 = 4'd15; a_sign2 = 4'd10; a_sign3 = 4'd8;
b_sign0 = 4'd10; b_sign1 = 4'd1; b_sign2 = 4'd13; b_sign3 = 4'd11;
@(posedge clk_i);
a_mant0 = 8'd6; a_mant1 = 8'd72; a_mant2 = 8'd42; a_mant3 = 8'd73;
b_mant0 = 8'd236; b_mant1 = 8'd189; b_mant2 = 8'd191; b_mant3 = 8'd253;
a_exp0 = 10'd934; a_exp1 = 10'd466; a_exp2 = 10'd64; a_exp3 = 10'd188;
b_exp0 = 10'd873; b_exp1 = 10'd881; b_exp2 = 10'd252; b_exp3 = 10'd829;
a_sign0 = 4'd5; a_sign1 = 4'd14; a_sign2 = 4'd15; a_sign3 = 4'd2;
b_sign0 = 4'd4; b_sign1 = 4'd10; b_sign2 = 4'd2; b_sign3 = 4'd12;
@(posedge clk_i);
a_mant0 = 8'd193; a_mant1 = 8'd54; a_mant2 = 8'd249; a_mant3 = 8'd56;
b_mant0 = 8'd169; b_mant1 = 8'd93; b_mant2 = 8'd15; b_mant3 = 8'd8;
a_exp0 = 10'd571; a_exp1 = 10'd590; a_exp2 = 10'd834; a_exp3 = 10'd909;
b_exp0 = 10'd919; b_exp1 = 10'd208; b_exp2 = 10'd400; b_exp3 = 10'd610;
a_sign0 = 4'd10; a_sign1 = 4'd15; a_sign2 = 4'd13; a_sign3 = 4'd10;
b_sign0 = 4'd13; b_sign1 = 4'd8; b_sign2 = 4'd2; b_sign3 = 4'd14;
@(posedge clk_i);
a_mant0 = 8'd193; a_mant1 = 8'd130; a_mant2 = 8'd210; a_mant3 = 8'd214;
b_mant0 = 8'd38; b_mant1 = 8'd90; b_mant2 = 8'd75; b_mant3 = 8'd112;
a_exp0 = 10'd46; a_exp1 = 10'd163; a_exp2 = 10'd970; a_exp3 = 10'd669;
b_exp0 = 10'd13; b_exp1 = 10'd87; b_exp2 = 10'd27; b_exp3 = 10'd805;
a_sign0 = 4'd11; a_sign1 = 4'd15; a_sign2 = 4'd10; a_sign3 = 4'd4;
b_sign0 = 4'd4; b_sign1 = 4'd2; b_sign2 = 4'd2; b_sign3 = 4'd5;
@(posedge clk_i);
a_mant0 = 8'd161; a_mant1 = 8'd87; a_mant2 = 8'd193; a_mant3 = 8'd62;
b_mant0 = 8'd63; b_mant1 = 8'd211; b_mant2 = 8'd81; b_mant3 = 8'd89;
a_exp0 = 10'd11; a_exp1 = 10'd569; a_exp2 = 10'd103; a_exp3 = 10'd417;
b_exp0 = 10'd824; b_exp1 = 10'd94; b_exp2 = 10'd599; b_exp3 = 10'd345;
a_sign0 = 4'd14; a_sign1 = 4'd1; a_sign2 = 4'd4; a_sign3 = 4'd11;
b_sign0 = 4'd4; b_sign1 = 4'd4; b_sign2 = 4'd7; b_sign3 = 4'd15;
@(posedge clk_i);
a_mant0 = 8'd191; a_mant1 = 8'd228; a_mant2 = 8'd62; a_mant3 = 8'd174;
b_mant0 = 8'd51; b_mant1 = 8'd246; b_mant2 = 8'd139; b_mant3 = 8'd87;
a_exp0 = 10'd671; a_exp1 = 10'd431; a_exp2 = 10'd148; a_exp3 = 10'd938;
b_exp0 = 10'd832; b_exp1 = 10'd31; b_exp2 = 10'd654; b_exp3 = 10'd305;
a_sign0 = 4'd10; a_sign1 = 4'd7; a_sign2 = 4'd4; a_sign3 = 4'd16;
b_sign0 = 4'd16; b_sign1 = 4'd10; b_sign2 = 4'd13; b_sign3 = 4'd12;
@(posedge clk_i);
a_mant0 = 8'd158; a_mant1 = 8'd85; a_mant2 = 8'd152; a_mant3 = 8'd124;
b_mant0 = 8'd53; b_mant1 = 8'd111; b_mant2 = 8'd179; b_mant3 = 8'd36;
a_exp0 = 10'd879; a_exp1 = 10'd948; a_exp2 = 10'd685; a_exp3 = 10'd793;
b_exp0 = 10'd518; b_exp1 = 10'd48; b_exp2 = 10'd641; b_exp3 = 10'd561;
a_sign0 = 4'd1; a_sign1 = 4'd14; a_sign2 = 4'd13; a_sign3 = 4'd1;
b_sign0 = 4'd0; b_sign1 = 4'd4; b_sign2 = 4'd2; b_sign3 = 4'd12;
@(posedge clk_i);
a_mant0 = 8'd236; a_mant1 = 8'd213; a_mant2 = 8'd71; a_mant3 = 8'd12;
b_mant0 = 8'd138; b_mant1 = 8'd129; b_mant2 = 8'd1; b_mant3 = 8'd130;
a_exp0 = 10'd561; a_exp1 = 10'd472; a_exp2 = 10'd840; a_exp3 = 10'd476;
b_exp0 = 10'd1006; b_exp1 = 10'd60; b_exp2 = 10'd663; b_exp3 = 10'd221;
a_sign0 = 4'd0; a_sign1 = 4'd13; a_sign2 = 4'd6; a_sign3 = 4'd14;
b_sign0 = 4'd3; b_sign1 = 4'd13; b_sign2 = 4'd4; b_sign3 = 4'd4;
@(posedge clk_i);
shared_exps0 = 8'd118;
shared_exps1 = 8'd123;
a_mant0 = 8'd245; a_mant1 = 8'd41; a_mant2 = 8'd234; a_mant3 = 8'd69;
b_mant0 = 8'd104; b_mant1 = 8'd101; b_mant2 = 8'd63; b_mant3 = 8'd48;
a_exp0 = 10'd687; a_exp1 = 10'd403; a_exp2 = 10'd979; a_exp3 = 10'd769;
b_exp0 = 10'd410; b_exp1 = 10'd514; b_exp2 = 10'd491; b_exp3 = 10'd705;
a_sign0 = 4'd9; a_sign1 = 4'd1; a_sign2 = 4'd12; a_sign3 = 4'd13;
b_sign0 = 4'd7; b_sign1 = 4'd6; b_sign2 = 4'd5; b_sign3 = 4'd0;
@(posedge clk_i);
a_mant0 = 8'd61; a_mant1 = 8'd179; a_mant2 = 8'd16; a_mant3 = 8'd65;
b_mant0 = 8'd154; b_mant1 = 8'd101; b_mant2 = 8'd41; b_mant3 = 8'd115;
a_exp0 = 10'd156; a_exp1 = 10'd674; a_exp2 = 10'd34; a_exp3 = 10'd453;
b_exp0 = 10'd923; b_exp1 = 10'd993; b_exp2 = 10'd155; b_exp3 = 10'd937;
a_sign0 = 4'd15; a_sign1 = 4'd1; a_sign2 = 4'd2; a_sign3 = 4'd5;
b_sign0 = 4'd11; b_sign1 = 4'd7; b_sign2 = 4'd5; b_sign3 = 4'd9;
@(posedge clk_i);
a_mant0 = 8'd181; a_mant1 = 8'd205; a_mant2 = 8'd180; a_mant3 = 8'd47;
b_mant0 = 8'd47; b_mant1 = 8'd26; b_mant2 = 8'd53; b_mant3 = 8'd126;
a_exp0 = 10'd413; a_exp1 = 10'd598; a_exp2 = 10'd597; a_exp3 = 10'd219;
b_exp0 = 10'd145; b_exp1 = 10'd921; b_exp2 = 10'd19; b_exp3 = 10'd983;
a_sign0 = 4'd7; a_sign1 = 4'd11; a_sign2 = 4'd11; a_sign3 = 4'd6;
b_sign0 = 4'd11; b_sign1 = 4'd2; b_sign2 = 4'd1; b_sign3 = 4'd9;
@(posedge clk_i);
a_mant0 = 8'd55; a_mant1 = 8'd243; a_mant2 = 8'd222; a_mant3 = 8'd122;
b_mant0 = 8'd201; b_mant1 = 8'd168; b_mant2 = 8'd216; b_mant3 = 8'd96;
a_exp0 = 10'd727; a_exp1 = 10'd697; a_exp2 = 10'd835; a_exp3 = 10'd588;
b_exp0 = 10'd428; b_exp1 = 10'd127; b_exp2 = 10'd773; b_exp3 = 10'd227;
a_sign0 = 4'd16; a_sign1 = 4'd1; a_sign2 = 4'd11; a_sign3 = 4'd3;
b_sign0 = 4'd8; b_sign1 = 4'd10; b_sign2 = 4'd14; b_sign3 = 4'd8;
@(posedge clk_i);
a_mant0 = 8'd117; a_mant1 = 8'd65; a_mant2 = 8'd116; a_mant3 = 8'd5;
b_mant0 = 8'd47; b_mant1 = 8'd236; b_mant2 = 8'd126; b_mant3 = 8'd13;
a_exp0 = 10'd296; a_exp1 = 10'd518; a_exp2 = 10'd183; a_exp3 = 10'd944;
b_exp0 = 10'd326; b_exp1 = 10'd602; b_exp2 = 10'd709; b_exp3 = 10'd836;
a_sign0 = 4'd3; a_sign1 = 4'd2; a_sign2 = 4'd6; a_sign3 = 4'd5;
b_sign0 = 4'd9; b_sign1 = 4'd8; b_sign2 = 4'd16; b_sign3 = 4'd0;
@(posedge clk_i);
a_mant0 = 8'd114; a_mant1 = 8'd167; a_mant2 = 8'd213; a_mant3 = 8'd96;
b_mant0 = 8'd229; b_mant1 = 8'd186; b_mant2 = 8'd136; b_mant3 = 8'd177;
a_exp0 = 10'd683; a_exp1 = 10'd446; a_exp2 = 10'd339; a_exp3 = 10'd630;
b_exp0 = 10'd285; b_exp1 = 10'd990; b_exp2 = 10'd303; b_exp3 = 10'd204;
a_sign0 = 4'd6; a_sign1 = 4'd15; a_sign2 = 4'd3; a_sign3 = 4'd14;
b_sign0 = 4'd16; b_sign1 = 4'd1; b_sign2 = 4'd3; b_sign3 = 4'd2;
@(posedge clk_i);
a_mant0 = 8'd109; a_mant1 = 8'd53; a_mant2 = 8'd132; a_mant3 = 8'd198;
b_mant0 = 8'd174; b_mant1 = 8'd154; b_mant2 = 8'd173; b_mant3 = 8'd54;
a_exp0 = 10'd61; a_exp1 = 10'd774; a_exp2 = 10'd664; a_exp3 = 10'd41;
b_exp0 = 10'd777; b_exp1 = 10'd154; b_exp2 = 10'd739; b_exp3 = 10'd486;
a_sign0 = 4'd8; a_sign1 = 4'd15; a_sign2 = 4'd8; a_sign3 = 4'd15;
b_sign0 = 4'd12; b_sign1 = 4'd7; b_sign2 = 4'd2; b_sign3 = 4'd16;
@(posedge clk_i);
a_mant0 = 8'd132; a_mant1 = 8'd245; a_mant2 = 8'd53; a_mant3 = 8'd177;
b_mant0 = 8'd153; b_mant1 = 8'd35; b_mant2 = 8'd29; b_mant3 = 8'd3;
a_exp0 = 10'd400; a_exp1 = 10'd415; a_exp2 = 10'd118; a_exp3 = 10'd607;
b_exp0 = 10'd948; b_exp1 = 10'd208; b_exp2 = 10'd344; b_exp3 = 10'd106;
a_sign0 = 4'd5; a_sign1 = 4'd7; a_sign2 = 4'd0; a_sign3 = 4'd16;
b_sign0 = 4'd8; b_sign1 = 4'd7; b_sign2 = 4'd7; b_sign3 = 4'd4;
@(posedge clk_i);
shared_exps0 = 8'd77;
shared_exps1 = 8'd130;
a_mant0 = 8'd183; a_mant1 = 8'd139; a_mant2 = 8'd116; a_mant3 = 8'd186;
b_mant0 = 8'd162; b_mant1 = 8'd211; b_mant2 = 8'd219; b_mant3 = 8'd109;
a_exp0 = 10'd1022; a_exp1 = 10'd269; a_exp2 = 10'd74; a_exp3 = 10'd615;
b_exp0 = 10'd722; b_exp1 = 10'd457; b_exp2 = 10'd60; b_exp3 = 10'd984;
a_sign0 = 4'd7; a_sign1 = 4'd15; a_sign2 = 4'd12; a_sign3 = 4'd14;
b_sign0 = 4'd7; b_sign1 = 4'd4; b_sign2 = 4'd9; b_sign3 = 4'd13;
@(posedge clk_i);
a_mant0 = 8'd55; a_mant1 = 8'd69; a_mant2 = 8'd118; a_mant3 = 8'd95;
b_mant0 = 8'd81; b_mant1 = 8'd85; b_mant2 = 8'd253; b_mant3 = 8'd4;
a_exp0 = 10'd656; a_exp1 = 10'd233; a_exp2 = 10'd492; a_exp3 = 10'd693;
b_exp0 = 10'd542; b_exp1 = 10'd92; b_exp2 = 10'd518; b_exp3 = 10'd651;
a_sign0 = 4'd0; a_sign1 = 4'd11; a_sign2 = 4'd7; a_sign3 = 4'd7;
b_sign0 = 4'd4; b_sign1 = 4'd12; b_sign2 = 4'd4; b_sign3 = 4'd6;
@(posedge clk_i);
a_mant0 = 8'd118; a_mant1 = 8'd234; a_mant2 = 8'd21; a_mant3 = 8'd49;
b_mant0 = 8'd186; b_mant1 = 8'd178; b_mant2 = 8'd17; b_mant3 = 8'd166;
a_exp0 = 10'd458; a_exp1 = 10'd845; a_exp2 = 10'd267; a_exp3 = 10'd71;
b_exp0 = 10'd550; b_exp1 = 10'd154; b_exp2 = 10'd50; b_exp3 = 10'd533;
a_sign0 = 4'd4; a_sign1 = 4'd7; a_sign2 = 4'd11; a_sign3 = 4'd9;
b_sign0 = 4'd8; b_sign1 = 4'd9; b_sign2 = 4'd5; b_sign3 = 4'd11;
@(posedge clk_i);
a_mant0 = 8'd188; a_mant1 = 8'd173; a_mant2 = 8'd139; a_mant3 = 8'd78;
b_mant0 = 8'd205; b_mant1 = 8'd90; b_mant2 = 8'd153; b_mant3 = 8'd3;
a_exp0 = 10'd717; a_exp1 = 10'd677; a_exp2 = 10'd588; a_exp3 = 10'd245;
b_exp0 = 10'd187; b_exp1 = 10'd803; b_exp2 = 10'd939; b_exp3 = 10'd105;
a_sign0 = 4'd9; a_sign1 = 4'd3; a_sign2 = 4'd9; a_sign3 = 4'd7;
b_sign0 = 4'd1; b_sign1 = 4'd5; b_sign2 = 4'd4; b_sign3 = 4'd15;
@(posedge clk_i);
a_mant0 = 8'd219; a_mant1 = 8'd115; a_mant2 = 8'd92; a_mant3 = 8'd162;
b_mant0 = 8'd154; b_mant1 = 8'd95; b_mant2 = 8'd175; b_mant3 = 8'd242;
a_exp0 = 10'd635; a_exp1 = 10'd667; a_exp2 = 10'd723; a_exp3 = 10'd1017;
b_exp0 = 10'd69; b_exp1 = 10'd946; b_exp2 = 10'd781; b_exp3 = 10'd236;
a_sign0 = 4'd5; a_sign1 = 4'd0; a_sign2 = 4'd13; a_sign3 = 4'd12;
b_sign0 = 4'd5; b_sign1 = 4'd16; b_sign2 = 4'd3; b_sign3 = 4'd7;
@(posedge clk_i);
a_mant0 = 8'd250; a_mant1 = 8'd92; a_mant2 = 8'd232; a_mant3 = 8'd120;
b_mant0 = 8'd233; b_mant1 = 8'd124; b_mant2 = 8'd60; b_mant3 = 8'd2;
a_exp0 = 10'd461; a_exp1 = 10'd833; a_exp2 = 10'd565; a_exp3 = 10'd869;
b_exp0 = 10'd390; b_exp1 = 10'd665; b_exp2 = 10'd796; b_exp3 = 10'd34;
a_sign0 = 4'd14; a_sign1 = 4'd10; a_sign2 = 4'd5; a_sign3 = 4'd7;
b_sign0 = 4'd14; b_sign1 = 4'd16; b_sign2 = 4'd15; b_sign3 = 4'd12;
@(posedge clk_i);
a_mant0 = 8'd204; a_mant1 = 8'd37; a_mant2 = 8'd142; a_mant3 = 8'd226;
b_mant0 = 8'd159; b_mant1 = 8'd21; b_mant2 = 8'd79; b_mant3 = 8'd45;
a_exp0 = 10'd572; a_exp1 = 10'd97; a_exp2 = 10'd395; a_exp3 = 10'd175;
b_exp0 = 10'd109; b_exp1 = 10'd815; b_exp2 = 10'd30; b_exp3 = 10'd365;
a_sign0 = 4'd14; a_sign1 = 4'd11; a_sign2 = 4'd15; a_sign3 = 4'd14;
b_sign0 = 4'd12; b_sign1 = 4'd2; b_sign2 = 4'd3; b_sign3 = 4'd4;
@(posedge clk_i);
a_mant0 = 8'd123; a_mant1 = 8'd80; a_mant2 = 8'd78; a_mant3 = 8'd192;
b_mant0 = 8'd130; b_mant1 = 8'd83; b_mant2 = 8'd5; b_mant3 = 8'd211;
a_exp0 = 10'd158; a_exp1 = 10'd474; a_exp2 = 10'd371; a_exp3 = 10'd875;
b_exp0 = 10'd161; b_exp1 = 10'd166; b_exp2 = 10'd102; b_exp3 = 10'd293;
a_sign0 = 4'd9; a_sign1 = 4'd6; a_sign2 = 4'd5; a_sign3 = 4'd12;
b_sign0 = 4'd14; b_sign1 = 4'd1; b_sign2 = 4'd16; b_sign3 = 4'd4;
@(posedge clk_i);
shared_exps0 = 8'd130;
shared_exps1 = 8'd137;
rstn = 0;
@(posedge clk_i);
rstn = 1;
a_mant0 = 8'd21; a_mant1 = 8'd44; a_mant2 = 8'd192; a_mant3 = 8'd90;
b_mant0 = 8'd14; b_mant1 = 8'd6; b_mant2 = 8'd211; b_mant3 = 8'd171;
a_exp0 = 10'd900; a_exp1 = 10'd37; a_exp2 = 10'd516; a_exp3 = 10'd761;
b_exp0 = 10'd589; b_exp1 = 10'd253; b_exp2 = 10'd56; b_exp3 = 10'd411;
a_sign0 = 4'd11; a_sign1 = 4'd14; a_sign2 = 4'd10; a_sign3 = 4'd1;
b_sign0 = 4'd6; b_sign1 = 4'd9; b_sign2 = 4'd14; b_sign3 = 4'd12;
@(posedge clk_i);
a_mant0 = 8'd33; a_mant1 = 8'd0; a_mant2 = 8'd73; a_mant3 = 8'd156;
b_mant0 = 8'd216; b_mant1 = 8'd166; b_mant2 = 8'd70; b_mant3 = 8'd85;
a_exp0 = 10'd47; a_exp1 = 10'd646; a_exp2 = 10'd474; a_exp3 = 10'd817;
b_exp0 = 10'd224; b_exp1 = 10'd682; b_exp2 = 10'd929; b_exp3 = 10'd159;
a_sign0 = 4'd2; a_sign1 = 4'd8; a_sign2 = 4'd13; a_sign3 = 4'd16;
b_sign0 = 4'd3; b_sign1 = 4'd6; b_sign2 = 4'd13; b_sign3 = 4'd4;
@(posedge clk_i);
a_mant0 = 8'd0; a_mant1 = 8'd1; a_mant2 = 8'd86; a_mant3 = 8'd245;
b_mant0 = 8'd1; b_mant1 = 8'd159; b_mant2 = 8'd146; b_mant3 = 8'd96;
a_exp0 = 10'd165; a_exp1 = 10'd239; a_exp2 = 10'd880; a_exp3 = 10'd914;
b_exp0 = 10'd934; b_exp1 = 10'd349; b_exp2 = 10'd353; b_exp3 = 10'd511;
a_sign0 = 4'd11; a_sign1 = 4'd2; a_sign2 = 4'd4; a_sign3 = 4'd8;
b_sign0 = 4'd9; b_sign1 = 4'd7; b_sign2 = 4'd11; b_sign3 = 4'd14;
@(posedge clk_i);
a_mant0 = 8'd208; a_mant1 = 8'd32; a_mant2 = 8'd111; a_mant3 = 8'd87;
b_mant0 = 8'd33; b_mant1 = 8'd20; b_mant2 = 8'd185; b_mant3 = 8'd105;
a_exp0 = 10'd864; a_exp1 = 10'd750; a_exp2 = 10'd744; a_exp3 = 10'd116;
b_exp0 = 10'd840; b_exp1 = 10'd624; b_exp2 = 10'd659; b_exp3 = 10'd70;
a_sign0 = 4'd12; a_sign1 = 4'd14; a_sign2 = 4'd0; a_sign3 = 4'd15;
b_sign0 = 4'd4; b_sign1 = 4'd5; b_sign2 = 4'd15; b_sign3 = 4'd6;
@(posedge clk_i);
a_mant0 = 8'd183; a_mant1 = 8'd101; a_mant2 = 8'd226; a_mant3 = 8'd126;
b_mant0 = 8'd2; b_mant1 = 8'd81; b_mant2 = 8'd235; b_mant3 = 8'd103;
a_exp0 = 10'd893; a_exp1 = 10'd216; a_exp2 = 10'd844; a_exp3 = 10'd199;
b_exp0 = 10'd635; b_exp1 = 10'd390; b_exp2 = 10'd1; b_exp3 = 10'd16;
a_sign0 = 4'd7; a_sign1 = 4'd4; a_sign2 = 4'd6; a_sign3 = 4'd7;
b_sign0 = 4'd11; b_sign1 = 4'd8; b_sign2 = 4'd7; b_sign3 = 4'd11;
@(posedge clk_i);
a_mant0 = 8'd232; a_mant1 = 8'd92; a_mant2 = 8'd32; a_mant3 = 8'd218;
b_mant0 = 8'd31; b_mant1 = 8'd50; b_mant2 = 8'd189; b_mant3 = 8'd189;
a_exp0 = 10'd771; a_exp1 = 10'd643; a_exp2 = 10'd173; a_exp3 = 10'd125;
b_exp0 = 10'd37; b_exp1 = 10'd362; b_exp2 = 10'd250; b_exp3 = 10'd577;
a_sign0 = 4'd15; a_sign1 = 4'd14; a_sign2 = 4'd9; a_sign3 = 4'd0;
b_sign0 = 4'd15; b_sign1 = 4'd0; b_sign2 = 4'd14; b_sign3 = 4'd1;
@(posedge clk_i);
a_mant0 = 8'd163; a_mant1 = 8'd52; a_mant2 = 8'd90; a_mant3 = 8'd169;
b_mant0 = 8'd25; b_mant1 = 8'd132; b_mant2 = 8'd243; b_mant3 = 8'd9;
a_exp0 = 10'd494; a_exp1 = 10'd671; a_exp2 = 10'd702; a_exp3 = 10'd348;
b_exp0 = 10'd129; b_exp1 = 10'd423; b_exp2 = 10'd385; b_exp3 = 10'd873;
a_sign0 = 4'd10; a_sign1 = 4'd3; a_sign2 = 4'd1; a_sign3 = 4'd16;
b_sign0 = 4'd14; b_sign1 = 4'd5; b_sign2 = 4'd4; b_sign3 = 4'd7;
@(posedge clk_i);
shared_exps0 = 8'd132;
shared_exps1 = 8'd116;
a_mant0 = 8'd90; a_mant1 = 8'd4; a_mant2 = 8'd149; a_mant3 = 8'd176;
b_mant0 = 8'd227; b_mant1 = 8'd135; b_mant2 = 8'd136; b_mant3 = 8'd43;
a_exp0 = 10'd270; a_exp1 = 10'd481; a_exp2 = 10'd833; a_exp3 = 10'd152;
b_exp0 = 10'd810; b_exp1 = 10'd661; b_exp2 = 10'd986; b_exp3 = 10'd415;
a_sign0 = 4'd2; a_sign1 = 4'd3; a_sign2 = 4'd1; a_sign3 = 4'd6;
b_sign0 = 4'd10; b_sign1 = 4'd4; b_sign2 = 4'd12; b_sign3 = 4'd5;
@(posedge clk_i);
a_mant0 = 8'd80; a_mant1 = 8'd211; a_mant2 = 8'd127; a_mant3 = 8'd95;
b_mant0 = 8'd245; b_mant1 = 8'd201; b_mant2 = 8'd78; b_mant3 = 8'd170;
a_exp0 = 10'd388; a_exp1 = 10'd246; a_exp2 = 10'd729; a_exp3 = 10'd1022;
b_exp0 = 10'd975; b_exp1 = 10'd120; b_exp2 = 10'd14; b_exp3 = 10'd954;
a_sign0 = 4'd11; a_sign1 = 4'd11; a_sign2 = 4'd6; a_sign3 = 4'd12;
b_sign0 = 4'd11; b_sign1 = 4'd4; b_sign2 = 4'd7; b_sign3 = 4'd11;
@(posedge clk_i);
a_mant0 = 8'd175; a_mant1 = 8'd250; a_mant2 = 8'd59; a_mant3 = 8'd218;
b_mant0 = 8'd161; b_mant1 = 8'd137; b_mant2 = 8'd243; b_mant3 = 8'd158;
a_exp0 = 10'd490; a_exp1 = 10'd132; a_exp2 = 10'd323; a_exp3 = 10'd358;
b_exp0 = 10'd543; b_exp1 = 10'd933; b_exp2 = 10'd416; b_exp3 = 10'd912;
a_sign0 = 4'd10; a_sign1 = 4'd9; a_sign2 = 4'd4; a_sign3 = 4'd5;
b_sign0 = 4'd12; b_sign1 = 4'd15; b_sign2 = 4'd13; b_sign3 = 4'd15;
@(posedge clk_i);
a_mant0 = 8'd136; a_mant1 = 8'd94; a_mant2 = 8'd148; a_mant3 = 8'd119;
b_mant0 = 8'd223; b_mant1 = 8'd222; b_mant2 = 8'd65; b_mant3 = 8'd202;
a_exp0 = 10'd824; a_exp1 = 10'd736; a_exp2 = 10'd877; a_exp3 = 10'd46;
b_exp0 = 10'd899; b_exp1 = 10'd439; b_exp2 = 10'd219; b_exp3 = 10'd661;
a_sign0 = 4'd14; a_sign1 = 4'd5; a_sign2 = 4'd7; a_sign3 = 4'd4;
b_sign0 = 4'd10; b_sign1 = 4'd16; b_sign2 = 4'd10; b_sign3 = 4'd15;
@(posedge clk_i);
a_mant0 = 8'd77; a_mant1 = 8'd121; a_mant2 = 8'd68; a_mant3 = 8'd232;
b_mant0 = 8'd217; b_mant1 = 8'd119; b_mant2 = 8'd144; b_mant3 = 8'd51;
a_exp0 = 10'd869; a_exp1 = 10'd705; a_exp2 = 10'd618; a_exp3 = 10'd720;
b_exp0 = 10'd745; b_exp1 = 10'd554; b_exp2 = 10'd308; b_exp3 = 10'd625;
a_sign0 = 4'd8; a_sign1 = 4'd9; a_sign2 = 4'd6; a_sign3 = 4'd7;
b_sign0 = 4'd13; b_sign1 = 4'd4; b_sign2 = 4'd7; b_sign3 = 4'd11;
@(posedge clk_i);
a_mant0 = 8'd146; a_mant1 = 8'd187; a_mant2 = 8'd109; a_mant3 = 8'd146;
b_mant0 = 8'd74; b_mant1 = 8'd239; b_mant2 = 8'd157; b_mant3 = 8'd192;
a_exp0 = 10'd365; a_exp1 = 10'd13; a_exp2 = 10'd770; a_exp3 = 10'd583;
b_exp0 = 10'd431; b_exp1 = 10'd639; b_exp2 = 10'd946; b_exp3 = 10'd936;
a_sign0 = 4'd2; a_sign1 = 4'd13; a_sign2 = 4'd1; a_sign3 = 4'd12;
b_sign0 = 4'd13; b_sign1 = 4'd9; b_sign2 = 4'd12; b_sign3 = 4'd1;
@(posedge clk_i);
a_mant0 = 8'd105; a_mant1 = 8'd83; a_mant2 = 8'd61; a_mant3 = 8'd166;
b_mant0 = 8'd9; b_mant1 = 8'd168; b_mant2 = 8'd96; b_mant3 = 8'd27;
a_exp0 = 10'd884; a_exp1 = 10'd571; a_exp2 = 10'd804; a_exp3 = 10'd106;
b_exp0 = 10'd938; b_exp1 = 10'd649; b_exp2 = 10'd147; b_exp3 = 10'd180;
a_sign0 = 4'd4; a_sign1 = 4'd7; a_sign2 = 4'd12; a_sign3 = 4'd3;
b_sign0 = 4'd11; b_sign1 = 4'd0; b_sign2 = 4'd5; b_sign3 = 4'd16;
@(posedge clk_i);
a_mant0 = 8'd114; a_mant1 = 8'd39; a_mant2 = 8'd245; a_mant3 = 8'd21;
b_mant0 = 8'd136; b_mant1 = 8'd147; b_mant2 = 8'd167; b_mant3 = 8'd45;
a_exp0 = 10'd533; a_exp1 = 10'd551; a_exp2 = 10'd914; a_exp3 = 10'd77;
b_exp0 = 10'd274; b_exp1 = 10'd772; b_exp2 = 10'd731; b_exp3 = 10'd639;
a_sign0 = 4'd10; a_sign1 = 4'd7; a_sign2 = 4'd6; a_sign3 = 4'd14;
b_sign0 = 4'd14; b_sign1 = 4'd13; b_sign2 = 4'd10; b_sign3 = 4'd15;
@(posedge clk_i);
shared_exps0 = 8'd140;
shared_exps1 = 8'd117;
a_mant0 = 8'd41; a_mant1 = 8'd230; a_mant2 = 8'd139; a_mant3 = 8'd86;
b_mant0 = 8'd238; b_mant1 = 8'd209; b_mant2 = 8'd50; b_mant3 = 8'd51;
a_exp0 = 10'd462; a_exp1 = 10'd677; a_exp2 = 10'd515; a_exp3 = 10'd267;
b_exp0 = 10'd54; b_exp1 = 10'd223; b_exp2 = 10'd646; b_exp3 = 10'd470;
a_sign0 = 4'd14; a_sign1 = 4'd3; a_sign2 = 4'd10; a_sign3 = 4'd10;
b_sign0 = 4'd1; b_sign1 = 4'd2; b_sign2 = 4'd14; b_sign3 = 4'd16;
@(posedge clk_i);
a_mant0 = 8'd2; a_mant1 = 8'd229; a_mant2 = 8'd83; a_mant3 = 8'd92;
b_mant0 = 8'd143; b_mant1 = 8'd221; b_mant2 = 8'd105; b_mant3 = 8'd239;
a_exp0 = 10'd621; a_exp1 = 10'd114; a_exp2 = 10'd124; a_exp3 = 10'd750;
b_exp0 = 10'd845; b_exp1 = 10'd581; b_exp2 = 10'd805; b_exp3 = 10'd99;
a_sign0 = 4'd16; a_sign1 = 4'd11; a_sign2 = 4'd6; a_sign3 = 4'd4;
b_sign0 = 4'd5; b_sign1 = 4'd7; b_sign2 = 4'd14; b_sign3 = 4'd4;
@(posedge clk_i);
a_mant0 = 8'd165; a_mant1 = 8'd5; a_mant2 = 8'd204; a_mant3 = 8'd160;
b_mant0 = 8'd133; b_mant1 = 8'd251; b_mant2 = 8'd175; b_mant3 = 8'd37;
a_exp0 = 10'd692; a_exp1 = 10'd645; a_exp2 = 10'd882; a_exp3 = 10'd196;
b_exp0 = 10'd882; b_exp1 = 10'd52; b_exp2 = 10'd220; b_exp3 = 10'd203;
a_sign0 = 4'd13; a_sign1 = 4'd2; a_sign2 = 4'd9; a_sign3 = 4'd7;
b_sign0 = 4'd13; b_sign1 = 4'd12; b_sign2 = 4'd10; b_sign3 = 4'd14;
@(posedge clk_i);
a_mant0 = 8'd16; a_mant1 = 8'd66; a_mant2 = 8'd99; a_mant3 = 8'd173;
b_mant0 = 8'd121; b_mant1 = 8'd201; b_mant2 = 8'd42; b_mant3 = 8'd209;
a_exp0 = 10'd186; a_exp1 = 10'd65; a_exp2 = 10'd956; a_exp3 = 10'd191;
b_exp0 = 10'd98; b_exp1 = 10'd930; b_exp2 = 10'd382; b_exp3 = 10'd398;
a_sign0 = 4'd5; a_sign1 = 4'd13; a_sign2 = 4'd13; a_sign3 = 4'd9;
b_sign0 = 4'd9; b_sign1 = 4'd13; b_sign2 = 4'd11; b_sign3 = 4'd8;
@(posedge clk_i);
a_mant0 = 8'd235; a_mant1 = 8'd68; a_mant2 = 8'd120; a_mant3 = 8'd43;
b_mant0 = 8'd254; b_mant1 = 8'd255; b_mant2 = 8'd90; b_mant3 = 8'd172;
a_exp0 = 10'd990; a_exp1 = 10'd498; a_exp2 = 10'd999; a_exp3 = 10'd520;
b_exp0 = 10'd897; b_exp1 = 10'd439; b_exp2 = 10'd327; b_exp3 = 10'd300;
a_sign0 = 4'd3; a_sign1 = 4'd5; a_sign2 = 4'd13; a_sign3 = 4'd9;
b_sign0 = 4'd15; b_sign1 = 4'd3; b_sign2 = 4'd8; b_sign3 = 4'd3;
@(posedge clk_i);
a_mant0 = 8'd209; a_mant1 = 8'd113; a_mant2 = 8'd150; a_mant3 = 8'd45;
b_mant0 = 8'd129; b_mant1 = 8'd68; b_mant2 = 8'd86; b_mant3 = 8'd219;
a_exp0 = 10'd941; a_exp1 = 10'd382; a_exp2 = 10'd96; a_exp3 = 10'd962;
b_exp0 = 10'd84; b_exp1 = 10'd922; b_exp2 = 10'd108; b_exp3 = 10'd77;
a_sign0 = 4'd14; a_sign1 = 4'd6; a_sign2 = 4'd6; a_sign3 = 4'd5;
b_sign0 = 4'd7; b_sign1 = 4'd0; b_sign2 = 4'd6; b_sign3 = 4'd9;
@(posedge clk_i);
a_mant0 = 8'd182; a_mant1 = 8'd1; a_mant2 = 8'd93; a_mant3 = 8'd102;
b_mant0 = 8'd103; b_mant1 = 8'd42; b_mant2 = 8'd139; b_mant3 = 8'd210;
a_exp0 = 10'd291; a_exp1 = 10'd680; a_exp2 = 10'd824; a_exp3 = 10'd924;
b_exp0 = 10'd627; b_exp1 = 10'd903; b_exp2 = 10'd201; b_exp3 = 10'd409;
a_sign0 = 4'd14; a_sign1 = 4'd12; a_sign2 = 4'd14; a_sign3 = 4'd10;
b_sign0 = 4'd10; b_sign1 = 4'd14; b_sign2 = 4'd8; b_sign3 = 4'd8;
@(posedge clk_i);
a_mant0 = 8'd255; a_mant1 = 8'd36; a_mant2 = 8'd216; a_mant3 = 8'd179;
b_mant0 = 8'd252; b_mant1 = 8'd11; b_mant2 = 8'd20; b_mant3 = 8'd10;
a_exp0 = 10'd931; a_exp1 = 10'd550; a_exp2 = 10'd833; a_exp3 = 10'd304;
b_exp0 = 10'd876; b_exp1 = 10'd4; b_exp2 = 10'd408; b_exp3 = 10'd817;
a_sign0 = 4'd11; a_sign1 = 4'd15; a_sign2 = 4'd0; a_sign3 = 4'd9;
b_sign0 = 4'd16; b_sign1 = 4'd6; b_sign2 = 4'd10; b_sign3 = 4'd7;
@(posedge clk_i);
shared_exps0 = 8'd141;
shared_exps1 = 8'd152;
a_mant0 = 8'd209; a_mant1 = 8'd247; a_mant2 = 8'd38; a_mant3 = 8'd7;
b_mant0 = 8'd72; b_mant1 = 8'd29; b_mant2 = 8'd55; b_mant3 = 8'd35;
a_exp0 = 10'd373; a_exp1 = 10'd775; a_exp2 = 10'd488; a_exp3 = 10'd954;
b_exp0 = 10'd942; b_exp1 = 10'd983; b_exp2 = 10'd719; b_exp3 = 10'd944;
a_sign0 = 4'd5; a_sign1 = 4'd10; a_sign2 = 4'd6; a_sign3 = 4'd6;
b_sign0 = 4'd0; b_sign1 = 4'd7; b_sign2 = 4'd2; b_sign3 = 4'd1;
@(posedge clk_i);
a_mant0 = 8'd42; a_mant1 = 8'd40; a_mant2 = 8'd91; a_mant3 = 8'd135;
b_mant0 = 8'd246; b_mant1 = 8'd84; b_mant2 = 8'd207; b_mant3 = 8'd191;
a_exp0 = 10'd605; a_exp1 = 10'd967; a_exp2 = 10'd713; a_exp3 = 10'd729;
b_exp0 = 10'd375; b_exp1 = 10'd293; b_exp2 = 10'd602; b_exp3 = 10'd328;
a_sign0 = 4'd10; a_sign1 = 4'd15; a_sign2 = 4'd10; a_sign3 = 4'd3;
b_sign0 = 4'd5; b_sign1 = 4'd5; b_sign2 = 4'd3; b_sign3 = 4'd13;
@(posedge clk_i);
a_mant0 = 8'd116; a_mant1 = 8'd235; a_mant2 = 8'd15; a_mant3 = 8'd37;
b_mant0 = 8'd140; b_mant1 = 8'd96; b_mant2 = 8'd198; b_mant3 = 8'd46;
a_exp0 = 10'd770; a_exp1 = 10'd43; a_exp2 = 10'd145; a_exp3 = 10'd582;
b_exp0 = 10'd362; b_exp1 = 10'd892; b_exp2 = 10'd249; b_exp3 = 10'd1004;
a_sign0 = 4'd2; a_sign1 = 4'd10; a_sign2 = 4'd3; a_sign3 = 4'd10;
b_sign0 = 4'd15; b_sign1 = 4'd7; b_sign2 = 4'd16; b_sign3 = 4'd12;
@(posedge clk_i);
a_mant0 = 8'd141; a_mant1 = 8'd121; a_mant2 = 8'd137; a_mant3 = 8'd127;
b_mant0 = 8'd239; b_mant1 = 8'd148; b_mant2 = 8'd165; b_mant3 = 8'd185;
a_exp0 = 10'd267; a_exp1 = 10'd1020; a_exp2 = 10'd771; a_exp3 = 10'd11;
b_exp0 = 10'd825; b_exp1 = 10'd946; b_exp2 = 10'd571; b_exp3 = 10'd459;
a_sign0 = 4'd8; a_sign1 = 4'd1; a_sign2 = 4'd8; a_sign3 = 4'd1;
b_sign0 = 4'd12; b_sign1 = 4'd2; b_sign2 = 4'd2; b_sign3 = 4'd16;
@(posedge clk_i);
a_mant0 = 8'd91; a_mant1 = 8'd252; a_mant2 = 8'd237; a_mant3 = 8'd104;
b_mant0 = 8'd117; b_mant1 = 8'd24; b_mant2 = 8'd108; b_mant3 = 8'd221;
a_exp0 = 10'd743; a_exp1 = 10'd158; a_exp2 = 10'd129; a_exp3 = 10'd554;
b_exp0 = 10'd3; b_exp1 = 10'd77; b_exp2 = 10'd981; b_exp3 = 10'd104;
a_sign0 = 4'd11; a_sign1 = 4'd12; a_sign2 = 4'd7; a_sign3 = 4'd0;
b_sign0 = 4'd10; b_sign1 = 4'd7; b_sign2 = 4'd6; b_sign3 = 4'd6;
@(posedge clk_i);
a_mant0 = 8'd6; a_mant1 = 8'd253; a_mant2 = 8'd184; a_mant3 = 8'd8;
b_mant0 = 8'd210; b_mant1 = 8'd68; b_mant2 = 8'd230; b_mant3 = 8'd3;
a_exp0 = 10'd21; a_exp1 = 10'd605; a_exp2 = 10'd334; a_exp3 = 10'd945;
b_exp0 = 10'd323; b_exp1 = 10'd282; b_exp2 = 10'd976; b_exp3 = 10'd700;
a_sign0 = 4'd16; a_sign1 = 4'd16; a_sign2 = 4'd1; a_sign3 = 4'd2;
b_sign0 = 4'd10; b_sign1 = 4'd0; b_sign2 = 4'd15; b_sign3 = 4'd13;
@(posedge clk_i);
a_mant0 = 8'd204; a_mant1 = 8'd50; a_mant2 = 8'd149; a_mant3 = 8'd72;
b_mant0 = 8'd241; b_mant1 = 8'd17; b_mant2 = 8'd24; b_mant3 = 8'd134;
a_exp0 = 10'd217; a_exp1 = 10'd222; a_exp2 = 10'd129; a_exp3 = 10'd541;
b_exp0 = 10'd657; b_exp1 = 10'd666; b_exp2 = 10'd737; b_exp3 = 10'd826;
a_sign0 = 4'd11; a_sign1 = 4'd14; a_sign2 = 4'd15; a_sign3 = 4'd10;
b_sign0 = 4'd8; b_sign1 = 4'd3; b_sign2 = 4'd12; b_sign3 = 4'd5;
@(posedge clk_i);
a_mant0 = 8'd42; a_mant1 = 8'd50; a_mant2 = 8'd63; a_mant3 = 8'd89;
b_mant0 = 8'd10; b_mant1 = 8'd204; b_mant2 = 8'd135; b_mant3 = 8'd156;
a_exp0 = 10'd197; a_exp1 = 10'd469; a_exp2 = 10'd875; a_exp3 = 10'd865;
b_exp0 = 10'd509; b_exp1 = 10'd362; b_exp2 = 10'd810; b_exp3 = 10'd518;
a_sign0 = 4'd5; a_sign1 = 4'd16; a_sign2 = 4'd16; a_sign3 = 4'd7;
b_sign0 = 4'd3; b_sign1 = 4'd2; b_sign2 = 4'd10; b_sign3 = 4'd9;
@(posedge clk_i);
shared_exps0 = 8'd129;
shared_exps1 = 8'd107;
rstn = 0;
@(posedge clk_i);
rstn = 1;
a_mant0 = 8'd123; a_mant1 = 8'd78; a_mant2 = 8'd32; a_mant3 = 8'd188;
b_mant0 = 8'd183; b_mant1 = 8'd123; b_mant2 = 8'd150; b_mant3 = 8'd137;
a_exp0 = 10'd886; a_exp1 = 10'd901; a_exp2 = 10'd245; a_exp3 = 10'd816;
b_exp0 = 10'd698; b_exp1 = 10'd908; b_exp2 = 10'd520; b_exp3 = 10'd557;
a_sign0 = 4'd12; a_sign1 = 4'd6; a_sign2 = 4'd7; a_sign3 = 4'd8;
b_sign0 = 4'd3; b_sign1 = 4'd3; b_sign2 = 4'd5; b_sign3 = 4'd14;
@(posedge clk_i);
a_mant0 = 8'd47; a_mant1 = 8'd24; a_mant2 = 8'd188; a_mant3 = 8'd141;
b_mant0 = 8'd97; b_mant1 = 8'd65; b_mant2 = 8'd114; b_mant3 = 8'd182;
a_exp0 = 10'd982; a_exp1 = 10'd790; a_exp2 = 10'd446; a_exp3 = 10'd272;
b_exp0 = 10'd258; b_exp1 = 10'd839; b_exp2 = 10'd481; b_exp3 = 10'd407;
a_sign0 = 4'd9; a_sign1 = 4'd3; a_sign2 = 4'd0; a_sign3 = 4'd12;
b_sign0 = 4'd8; b_sign1 = 4'd7; b_sign2 = 4'd16; b_sign3 = 4'd1;
@(posedge clk_i);
a_mant0 = 8'd36; a_mant1 = 8'd172; a_mant2 = 8'd133; a_mant3 = 8'd242;
b_mant0 = 8'd94; b_mant1 = 8'd125; b_mant2 = 8'd63; b_mant3 = 8'd66;
a_exp0 = 10'd593; a_exp1 = 10'd907; a_exp2 = 10'd193; a_exp3 = 10'd129;
b_exp0 = 10'd579; b_exp1 = 10'd889; b_exp2 = 10'd700; b_exp3 = 10'd605;
a_sign0 = 4'd4; a_sign1 = 4'd14; a_sign2 = 4'd5; a_sign3 = 4'd14;
b_sign0 = 4'd6; b_sign1 = 4'd11; b_sign2 = 4'd9; b_sign3 = 4'd12;
@(posedge clk_i);
a_mant0 = 8'd14; a_mant1 = 8'd209; a_mant2 = 8'd210; a_mant3 = 8'd80;
b_mant0 = 8'd219; b_mant1 = 8'd153; b_mant2 = 8'd184; b_mant3 = 8'd70;
a_exp0 = 10'd944; a_exp1 = 10'd742; a_exp2 = 10'd781; a_exp3 = 10'd104;
b_exp0 = 10'd130; b_exp1 = 10'd453; b_exp2 = 10'd753; b_exp3 = 10'd869;
a_sign0 = 4'd10; a_sign1 = 4'd4; a_sign2 = 4'd13; a_sign3 = 4'd8;
b_sign0 = 4'd9; b_sign1 = 4'd1; b_sign2 = 4'd12; b_sign3 = 4'd5;
@(posedge clk_i);
a_mant0 = 8'd45; a_mant1 = 8'd24; a_mant2 = 8'd134; a_mant3 = 8'd16;
b_mant0 = 8'd82; b_mant1 = 8'd196; b_mant2 = 8'd132; b_mant3 = 8'd113;
a_exp0 = 10'd934; a_exp1 = 10'd757; a_exp2 = 10'd927; a_exp3 = 10'd809;
b_exp0 = 10'd154; b_exp1 = 10'd1021; b_exp2 = 10'd1019; b_exp3 = 10'd142;
a_sign0 = 4'd0; a_sign1 = 4'd1; a_sign2 = 4'd4; a_sign3 = 4'd13;
b_sign0 = 4'd4; b_sign1 = 4'd6; b_sign2 = 4'd5; b_sign3 = 4'd15;
@(posedge clk_i);
a_mant0 = 8'd246; a_mant1 = 8'd153; a_mant2 = 8'd233; a_mant3 = 8'd18;
b_mant0 = 8'd34; b_mant1 = 8'd97; b_mant2 = 8'd138; b_mant3 = 8'd152;
a_exp0 = 10'd913; a_exp1 = 10'd999; a_exp2 = 10'd890; a_exp3 = 10'd411;
b_exp0 = 10'd978; b_exp1 = 10'd385; b_exp2 = 10'd503; b_exp3 = 10'd945;
a_sign0 = 4'd8; a_sign1 = 4'd5; a_sign2 = 4'd7; a_sign3 = 4'd5;
b_sign0 = 4'd11; b_sign1 = 4'd13; b_sign2 = 4'd7; b_sign3 = 4'd9;
@(posedge clk_i);
a_mant0 = 8'd199; a_mant1 = 8'd87; a_mant2 = 8'd2; a_mant3 = 8'd188;
b_mant0 = 8'd64; b_mant1 = 8'd198; b_mant2 = 8'd251; b_mant3 = 8'd0;
a_exp0 = 10'd453; a_exp1 = 10'd226; a_exp2 = 10'd27; a_exp3 = 10'd837;
b_exp0 = 10'd873; b_exp1 = 10'd439; b_exp2 = 10'd209; b_exp3 = 10'd632;
a_sign0 = 4'd10; a_sign1 = 4'd11; a_sign2 = 4'd8; a_sign3 = 4'd2;
b_sign0 = 4'd8; b_sign1 = 4'd7; b_sign2 = 4'd12; b_sign3 = 4'd3;
@(posedge clk_i);
shared_exps0 = 8'd110;
shared_exps1 = 8'd135;
a_mant0 = 8'd42; a_mant1 = 8'd132; a_mant2 = 8'd103; a_mant3 = 8'd129;
b_mant0 = 8'd159; b_mant1 = 8'd41; b_mant2 = 8'd56; b_mant3 = 8'd68;
a_exp0 = 10'd928; a_exp1 = 10'd278; a_exp2 = 10'd1017; a_exp3 = 10'd359;
b_exp0 = 10'd371; b_exp1 = 10'd550; b_exp2 = 10'd555; b_exp3 = 10'd919;
a_sign0 = 4'd11; a_sign1 = 4'd2; a_sign2 = 4'd12; a_sign3 = 4'd12;
b_sign0 = 4'd0; b_sign1 = 4'd12; b_sign2 = 4'd14; b_sign3 = 4'd14;
@(posedge clk_i);
a_mant0 = 8'd40; a_mant1 = 8'd161; a_mant2 = 8'd184; a_mant3 = 8'd123;
b_mant0 = 8'd169; b_mant1 = 8'd206; b_mant2 = 8'd108; b_mant3 = 8'd255;
a_exp0 = 10'd1011; a_exp1 = 10'd335; a_exp2 = 10'd470; a_exp3 = 10'd599;
b_exp0 = 10'd580; b_exp1 = 10'd712; b_exp2 = 10'd990; b_exp3 = 10'd1015;
a_sign0 = 4'd14; a_sign1 = 4'd3; a_sign2 = 4'd6; a_sign3 = 4'd16;
b_sign0 = 4'd6; b_sign1 = 4'd4; b_sign2 = 4'd1; b_sign3 = 4'd7;
@(posedge clk_i);
a_mant0 = 8'd194; a_mant1 = 8'd39; a_mant2 = 8'd243; a_mant3 = 8'd104;
b_mant0 = 8'd35; b_mant1 = 8'd97; b_mant2 = 8'd25; b_mant3 = 8'd5;
a_exp0 = 10'd474; a_exp1 = 10'd1023; a_exp2 = 10'd20; a_exp3 = 10'd11;
b_exp0 = 10'd444; b_exp1 = 10'd296; b_exp2 = 10'd744; b_exp3 = 10'd942;
a_sign0 = 4'd7; a_sign1 = 4'd1; a_sign2 = 4'd5; a_sign3 = 4'd2;
b_sign0 = 4'd3; b_sign1 = 4'd8; b_sign2 = 4'd10; b_sign3 = 4'd9;
@(posedge clk_i);
a_mant0 = 8'd19; a_mant1 = 8'd152; a_mant2 = 8'd16; a_mant3 = 8'd182;
b_mant0 = 8'd235; b_mant1 = 8'd18; b_mant2 = 8'd138; b_mant3 = 8'd41;
a_exp0 = 10'd487; a_exp1 = 10'd861; a_exp2 = 10'd37; a_exp3 = 10'd195;
b_exp0 = 10'd524; b_exp1 = 10'd480; b_exp2 = 10'd369; b_exp3 = 10'd992;
a_sign0 = 4'd6; a_sign1 = 4'd1; a_sign2 = 4'd11; a_sign3 = 4'd13;
b_sign0 = 4'd1; b_sign1 = 4'd6; b_sign2 = 4'd12; b_sign3 = 4'd9;
@(posedge clk_i);
a_mant0 = 8'd188; a_mant1 = 8'd184; a_mant2 = 8'd236; a_mant3 = 8'd215;
b_mant0 = 8'd183; b_mant1 = 8'd7; b_mant2 = 8'd3; b_mant3 = 8'd95;
a_exp0 = 10'd659; a_exp1 = 10'd85; a_exp2 = 10'd78; a_exp3 = 10'd215;
b_exp0 = 10'd341; b_exp1 = 10'd93; b_exp2 = 10'd401; b_exp3 = 10'd56;
a_sign0 = 4'd13; a_sign1 = 4'd6; a_sign2 = 4'd5; a_sign3 = 4'd9;
b_sign0 = 4'd1; b_sign1 = 4'd10; b_sign2 = 4'd5; b_sign3 = 4'd2;
@(posedge clk_i);
a_mant0 = 8'd46; a_mant1 = 8'd106; a_mant2 = 8'd226; a_mant3 = 8'd63;
b_mant0 = 8'd3; b_mant1 = 8'd171; b_mant2 = 8'd39; b_mant3 = 8'd16;
a_exp0 = 10'd706; a_exp1 = 10'd590; a_exp2 = 10'd745; a_exp3 = 10'd534;
b_exp0 = 10'd761; b_exp1 = 10'd317; b_exp2 = 10'd179; b_exp3 = 10'd28;
a_sign0 = 4'd4; a_sign1 = 4'd3; a_sign2 = 4'd9; a_sign3 = 4'd14;
b_sign0 = 4'd9; b_sign1 = 4'd8; b_sign2 = 4'd6; b_sign3 = 4'd2;
@(posedge clk_i);
a_mant0 = 8'd24; a_mant1 = 8'd234; a_mant2 = 8'd199; a_mant3 = 8'd216;
b_mant0 = 8'd69; b_mant1 = 8'd27; b_mant2 = 8'd202; b_mant3 = 8'd10;
a_exp0 = 10'd216; a_exp1 = 10'd345; a_exp2 = 10'd463; a_exp3 = 10'd803;
b_exp0 = 10'd289; b_exp1 = 10'd202; b_exp2 = 10'd439; b_exp3 = 10'd590;
a_sign0 = 4'd6; a_sign1 = 4'd2; a_sign2 = 4'd10; a_sign3 = 4'd12;
b_sign0 = 4'd11; b_sign1 = 4'd4; b_sign2 = 4'd1; b_sign3 = 4'd10;
@(posedge clk_i);
a_mant0 = 8'd31; a_mant1 = 8'd83; a_mant2 = 8'd222; a_mant3 = 8'd156;
b_mant0 = 8'd253; b_mant1 = 8'd135; b_mant2 = 8'd19; b_mant3 = 8'd210;
a_exp0 = 10'd641; a_exp1 = 10'd708; a_exp2 = 10'd80; a_exp3 = 10'd645;
b_exp0 = 10'd432; b_exp1 = 10'd859; b_exp2 = 10'd803; b_exp3 = 10'd828;
a_sign0 = 4'd11; a_sign1 = 4'd10; a_sign2 = 4'd9; a_sign3 = 4'd3;
b_sign0 = 4'd3; b_sign1 = 4'd6; b_sign2 = 4'd15; b_sign3 = 4'd0;
@(posedge clk_i);
shared_exps0 = 8'd142;
shared_exps1 = 8'd126;
a_mant0 = 8'd141; a_mant1 = 8'd48; a_mant2 = 8'd248; a_mant3 = 8'd207;
b_mant0 = 8'd194; b_mant1 = 8'd26; b_mant2 = 8'd82; b_mant3 = 8'd192;
a_exp0 = 10'd533; a_exp1 = 10'd270; a_exp2 = 10'd986; a_exp3 = 10'd109;
b_exp0 = 10'd197; b_exp1 = 10'd81; b_exp2 = 10'd855; b_exp3 = 10'd637;
a_sign0 = 4'd7; a_sign1 = 4'd2; a_sign2 = 4'd5; a_sign3 = 4'd11;
b_sign0 = 4'd16; b_sign1 = 4'd3; b_sign2 = 4'd13; b_sign3 = 4'd12;
@(posedge clk_i);
a_mant0 = 8'd47; a_mant1 = 8'd135; a_mant2 = 8'd217; a_mant3 = 8'd75;
b_mant0 = 8'd99; b_mant1 = 8'd145; b_mant2 = 8'd13; b_mant3 = 8'd150;
a_exp0 = 10'd743; a_exp1 = 10'd380; a_exp2 = 10'd497; a_exp3 = 10'd483;
b_exp0 = 10'd485; b_exp1 = 10'd560; b_exp2 = 10'd980; b_exp3 = 10'd656;
a_sign0 = 4'd13; a_sign1 = 4'd8; a_sign2 = 4'd13; a_sign3 = 4'd7;
b_sign0 = 4'd7; b_sign1 = 4'd16; b_sign2 = 4'd6; b_sign3 = 4'd14;
@(posedge clk_i);
a_mant0 = 8'd162; a_mant1 = 8'd34; a_mant2 = 8'd205; a_mant3 = 8'd15;
b_mant0 = 8'd10; b_mant1 = 8'd30; b_mant2 = 8'd212; b_mant3 = 8'd9;
a_exp0 = 10'd208; a_exp1 = 10'd704; a_exp2 = 10'd436; a_exp3 = 10'd706;
b_exp0 = 10'd495; b_exp1 = 10'd577; b_exp2 = 10'd157; b_exp3 = 10'd806;
a_sign0 = 4'd1; a_sign1 = 4'd13; a_sign2 = 4'd4; a_sign3 = 4'd3;
b_sign0 = 4'd3; b_sign1 = 4'd2; b_sign2 = 4'd4; b_sign3 = 4'd15;
@(posedge clk_i);
a_mant0 = 8'd123; a_mant1 = 8'd31; a_mant2 = 8'd248; a_mant3 = 8'd44;
b_mant0 = 8'd60; b_mant1 = 8'd164; b_mant2 = 8'd147; b_mant3 = 8'd235;
a_exp0 = 10'd254; a_exp1 = 10'd975; a_exp2 = 10'd242; a_exp3 = 10'd733;
b_exp0 = 10'd661; b_exp1 = 10'd552; b_exp2 = 10'd376; b_exp3 = 10'd461;
a_sign0 = 4'd0; a_sign1 = 4'd0; a_sign2 = 4'd5; a_sign3 = 4'd8;
b_sign0 = 4'd9; b_sign1 = 4'd1; b_sign2 = 4'd6; b_sign3 = 4'd6;
@(posedge clk_i);
a_mant0 = 8'd96; a_mant1 = 8'd110; a_mant2 = 8'd68; a_mant3 = 8'd51;
b_mant0 = 8'd19; b_mant1 = 8'd180; b_mant2 = 8'd66; b_mant3 = 8'd228;
a_exp0 = 10'd109; a_exp1 = 10'd31; a_exp2 = 10'd707; a_exp3 = 10'd668;
b_exp0 = 10'd589; b_exp1 = 10'd517; b_exp2 = 10'd778; b_exp3 = 10'd129;
a_sign0 = 4'd3; a_sign1 = 4'd11; a_sign2 = 4'd4; a_sign3 = 4'd5;
b_sign0 = 4'd4; b_sign1 = 4'd14; b_sign2 = 4'd12; b_sign3 = 4'd9;
@(posedge clk_i);
a_mant0 = 8'd15; a_mant1 = 8'd40; a_mant2 = 8'd201; a_mant3 = 8'd111;
b_mant0 = 8'd10; b_mant1 = 8'd97; b_mant2 = 8'd190; b_mant3 = 8'd81;
a_exp0 = 10'd883; a_exp1 = 10'd188; a_exp2 = 10'd40; a_exp3 = 10'd478;
b_exp0 = 10'd162; b_exp1 = 10'd701; b_exp2 = 10'd992; b_exp3 = 10'd280;
a_sign0 = 4'd8; a_sign1 = 4'd0; a_sign2 = 4'd12; a_sign3 = 4'd3;
b_sign0 = 4'd14; b_sign1 = 4'd12; b_sign2 = 4'd5; b_sign3 = 4'd14;
@(posedge clk_i);
a_mant0 = 8'd42; a_mant1 = 8'd138; a_mant2 = 8'd48; a_mant3 = 8'd44;
b_mant0 = 8'd43; b_mant1 = 8'd117; b_mant2 = 8'd223; b_mant3 = 8'd59;
a_exp0 = 10'd643; a_exp1 = 10'd606; a_exp2 = 10'd623; a_exp3 = 10'd612;
b_exp0 = 10'd33; b_exp1 = 10'd252; b_exp2 = 10'd234; b_exp3 = 10'd207;
a_sign0 = 4'd0; a_sign1 = 4'd9; a_sign2 = 4'd1; a_sign3 = 4'd4;
b_sign0 = 4'd11; b_sign1 = 4'd4; b_sign2 = 4'd9; b_sign3 = 4'd6;
@(posedge clk_i);
a_mant0 = 8'd89; a_mant1 = 8'd52; a_mant2 = 8'd228; a_mant3 = 8'd130;
b_mant0 = 8'd88; b_mant1 = 8'd30; b_mant2 = 8'd153; b_mant3 = 8'd84;
a_exp0 = 10'd424; a_exp1 = 10'd400; a_exp2 = 10'd41; a_exp3 = 10'd497;
b_exp0 = 10'd342; b_exp1 = 10'd309; b_exp2 = 10'd914; b_exp3 = 10'd442;
a_sign0 = 4'd16; a_sign1 = 4'd4; a_sign2 = 4'd15; a_sign3 = 4'd2;
b_sign0 = 4'd1; b_sign1 = 4'd4; b_sign2 = 4'd6; b_sign3 = 4'd13;
@(posedge clk_i);
shared_exps0 = 8'd114;
shared_exps1 = 8'd127;
a_mant0 = 8'd57; a_mant1 = 8'd179; a_mant2 = 8'd41; a_mant3 = 8'd185;
b_mant0 = 8'd133; b_mant1 = 8'd41; b_mant2 = 8'd149; b_mant3 = 8'd6;
a_exp0 = 10'd610; a_exp1 = 10'd439; a_exp2 = 10'd90; a_exp3 = 10'd832;
b_exp0 = 10'd740; b_exp1 = 10'd515; b_exp2 = 10'd310; b_exp3 = 10'd464;
a_sign0 = 4'd3; a_sign1 = 4'd4; a_sign2 = 4'd11; a_sign3 = 4'd8;
b_sign0 = 4'd2; b_sign1 = 4'd11; b_sign2 = 4'd1; b_sign3 = 4'd9;
@(posedge clk_i);
a_mant0 = 8'd121; a_mant1 = 8'd91; a_mant2 = 8'd37; a_mant3 = 8'd109;
b_mant0 = 8'd120; b_mant1 = 8'd166; b_mant2 = 8'd251; b_mant3 = 8'd15;
a_exp0 = 10'd16; a_exp1 = 10'd432; a_exp2 = 10'd13; a_exp3 = 10'd74;
b_exp0 = 10'd414; b_exp1 = 10'd149; b_exp2 = 10'd601; b_exp3 = 10'd725;
a_sign0 = 4'd11; a_sign1 = 4'd7; a_sign2 = 4'd14; a_sign3 = 4'd15;
b_sign0 = 4'd16; b_sign1 = 4'd15; b_sign2 = 4'd0; b_sign3 = 4'd14;
@(posedge clk_i);
a_mant0 = 8'd111; a_mant1 = 8'd198; a_mant2 = 8'd45; a_mant3 = 8'd146;
b_mant0 = 8'd110; b_mant1 = 8'd234; b_mant2 = 8'd151; b_mant3 = 8'd131;
a_exp0 = 10'd575; a_exp1 = 10'd271; a_exp2 = 10'd180; a_exp3 = 10'd770;
b_exp0 = 10'd111; b_exp1 = 10'd715; b_exp2 = 10'd559; b_exp3 = 10'd792;
a_sign0 = 4'd13; a_sign1 = 4'd10; a_sign2 = 4'd7; a_sign3 = 4'd14;
b_sign0 = 4'd13; b_sign1 = 4'd4; b_sign2 = 4'd13; b_sign3 = 4'd5;
@(posedge clk_i);
a_mant0 = 8'd136; a_mant1 = 8'd42; a_mant2 = 8'd134; a_mant3 = 8'd207;
b_mant0 = 8'd243; b_mant1 = 8'd137; b_mant2 = 8'd188; b_mant3 = 8'd118;
a_exp0 = 10'd491; a_exp1 = 10'd84; a_exp2 = 10'd269; a_exp3 = 10'd534;
b_exp0 = 10'd591; b_exp1 = 10'd236; b_exp2 = 10'd207; b_exp3 = 10'd19;
a_sign0 = 4'd11; a_sign1 = 4'd6; a_sign2 = 4'd3; a_sign3 = 4'd16;
b_sign0 = 4'd12; b_sign1 = 4'd16; b_sign2 = 4'd9; b_sign3 = 4'd2;
@(posedge clk_i);
a_mant0 = 8'd142; a_mant1 = 8'd148; a_mant2 = 8'd31; a_mant3 = 8'd56;
b_mant0 = 8'd190; b_mant1 = 8'd29; b_mant2 = 8'd3; b_mant3 = 8'd223;
a_exp0 = 10'd64; a_exp1 = 10'd973; a_exp2 = 10'd159; a_exp3 = 10'd1017;
b_exp0 = 10'd338; b_exp1 = 10'd977; b_exp2 = 10'd643; b_exp3 = 10'd444;
a_sign0 = 4'd0; a_sign1 = 4'd9; a_sign2 = 4'd9; a_sign3 = 4'd13;
b_sign0 = 4'd15; b_sign1 = 4'd4; b_sign2 = 4'd9; b_sign3 = 4'd14;
@(posedge clk_i);
a_mant0 = 8'd93; a_mant1 = 8'd94; a_mant2 = 8'd11; a_mant3 = 8'd221;
b_mant0 = 8'd139; b_mant1 = 8'd2; b_mant2 = 8'd179; b_mant3 = 8'd66;
a_exp0 = 10'd1021; a_exp1 = 10'd798; a_exp2 = 10'd159; a_exp3 = 10'd714;
b_exp0 = 10'd869; b_exp1 = 10'd496; b_exp2 = 10'd777; b_exp3 = 10'd77;
a_sign0 = 4'd4; a_sign1 = 4'd3; a_sign2 = 4'd0; a_sign3 = 4'd16;
b_sign0 = 4'd2; b_sign1 = 4'd10; b_sign2 = 4'd14; b_sign3 = 4'd6;
@(posedge clk_i);
a_mant0 = 8'd34; a_mant1 = 8'd51; a_mant2 = 8'd41; a_mant3 = 8'd164;
b_mant0 = 8'd199; b_mant1 = 8'd144; b_mant2 = 8'd197; b_mant3 = 8'd184;
a_exp0 = 10'd418; a_exp1 = 10'd369; a_exp2 = 10'd464; a_exp3 = 10'd740;
b_exp0 = 10'd522; b_exp1 = 10'd612; b_exp2 = 10'd358; b_exp3 = 10'd756;
a_sign0 = 4'd3; a_sign1 = 4'd15; a_sign2 = 4'd14; a_sign3 = 4'd0;
b_sign0 = 4'd1; b_sign1 = 4'd16; b_sign2 = 4'd15; b_sign3 = 4'd0;
@(posedge clk_i);
a_mant0 = 8'd148; a_mant1 = 8'd10; a_mant2 = 8'd147; a_mant3 = 8'd179;
b_mant0 = 8'd183; b_mant1 = 8'd84; b_mant2 = 8'd20; b_mant3 = 8'd35;
a_exp0 = 10'd3; a_exp1 = 10'd922; a_exp2 = 10'd483; a_exp3 = 10'd698;
b_exp0 = 10'd1001; b_exp1 = 10'd541; b_exp2 = 10'd788; b_exp3 = 10'd210;
a_sign0 = 4'd12; a_sign1 = 4'd14; a_sign2 = 4'd16; a_sign3 = 4'd8;
b_sign0 = 4'd3; b_sign1 = 4'd16; b_sign2 = 4'd8; b_sign3 = 4'd15;
@(posedge clk_i);
shared_exps0 = 8'd135;
shared_exps1 = 8'd144;
rstn = 0;
@(posedge clk_i);
rstn = 1;
a_mant0 = 8'd188; a_mant1 = 8'd169; a_mant2 = 8'd255; a_mant3 = 8'd203;
b_mant0 = 8'd21; b_mant1 = 8'd57; b_mant2 = 8'd91; b_mant3 = 8'd218;
a_exp0 = 10'd335; a_exp1 = 10'd525; a_exp2 = 10'd318; a_exp3 = 10'd438;
b_exp0 = 10'd186; b_exp1 = 10'd701; b_exp2 = 10'd744; b_exp3 = 10'd1011;
a_sign0 = 4'd12; a_sign1 = 4'd11; a_sign2 = 4'd1; a_sign3 = 4'd13;
b_sign0 = 4'd3; b_sign1 = 4'd3; b_sign2 = 4'd1; b_sign3 = 4'd8;
@(posedge clk_i);
a_mant0 = 8'd72; a_mant1 = 8'd215; a_mant2 = 8'd96; a_mant3 = 8'd76;
b_mant0 = 8'd190; b_mant1 = 8'd165; b_mant2 = 8'd44; b_mant3 = 8'd167;
a_exp0 = 10'd156; a_exp1 = 10'd454; a_exp2 = 10'd8; a_exp3 = 10'd476;
b_exp0 = 10'd872; b_exp1 = 10'd81; b_exp2 = 10'd890; b_exp3 = 10'd930;
a_sign0 = 4'd6; a_sign1 = 4'd15; a_sign2 = 4'd13; a_sign3 = 4'd7;
b_sign0 = 4'd12; b_sign1 = 4'd15; b_sign2 = 4'd16; b_sign3 = 4'd16;
@(posedge clk_i);
a_mant0 = 8'd57; a_mant1 = 8'd171; a_mant2 = 8'd200; a_mant3 = 8'd141;
b_mant0 = 8'd126; b_mant1 = 8'd158; b_mant2 = 8'd7; b_mant3 = 8'd176;
a_exp0 = 10'd86; a_exp1 = 10'd271; a_exp2 = 10'd276; a_exp3 = 10'd988;
b_exp0 = 10'd332; b_exp1 = 10'd441; b_exp2 = 10'd867; b_exp3 = 10'd983;
a_sign0 = 4'd0; a_sign1 = 4'd11; a_sign2 = 4'd9; a_sign3 = 4'd6;
b_sign0 = 4'd4; b_sign1 = 4'd1; b_sign2 = 4'd14; b_sign3 = 4'd13;
@(posedge clk_i);
a_mant0 = 8'd93; a_mant1 = 8'd78; a_mant2 = 8'd186; a_mant3 = 8'd136;
b_mant0 = 8'd213; b_mant1 = 8'd254; b_mant2 = 8'd135; b_mant3 = 8'd57;
a_exp0 = 10'd888; a_exp1 = 10'd305; a_exp2 = 10'd659; a_exp3 = 10'd12;
b_exp0 = 10'd692; b_exp1 = 10'd360; b_exp2 = 10'd268; b_exp3 = 10'd468;
a_sign0 = 4'd2; a_sign1 = 4'd13; a_sign2 = 4'd5; a_sign3 = 4'd8;
b_sign0 = 4'd10; b_sign1 = 4'd6; b_sign2 = 4'd3; b_sign3 = 4'd12;
@(posedge clk_i);
a_mant0 = 8'd227; a_mant1 = 8'd218; a_mant2 = 8'd203; a_mant3 = 8'd238;
b_mant0 = 8'd52; b_mant1 = 8'd183; b_mant2 = 8'd67; b_mant3 = 8'd239;
a_exp0 = 10'd676; a_exp1 = 10'd813; a_exp2 = 10'd769; a_exp3 = 10'd846;
b_exp0 = 10'd555; b_exp1 = 10'd714; b_exp2 = 10'd852; b_exp3 = 10'd508;
a_sign0 = 4'd3; a_sign1 = 4'd5; a_sign2 = 4'd14; a_sign3 = 4'd12;
b_sign0 = 4'd10; b_sign1 = 4'd6; b_sign2 = 4'd4; b_sign3 = 4'd6;
@(posedge clk_i);
a_mant0 = 8'd184; a_mant1 = 8'd98; a_mant2 = 8'd105; a_mant3 = 8'd239;
b_mant0 = 8'd187; b_mant1 = 8'd1; b_mant2 = 8'd16; b_mant3 = 8'd64;
a_exp0 = 10'd780; a_exp1 = 10'd694; a_exp2 = 10'd819; a_exp3 = 10'd801;
b_exp0 = 10'd26; b_exp1 = 10'd348; b_exp2 = 10'd526; b_exp3 = 10'd688;
a_sign0 = 4'd7; a_sign1 = 4'd1; a_sign2 = 4'd1; a_sign3 = 4'd7;
b_sign0 = 4'd2; b_sign1 = 4'd9; b_sign2 = 4'd13; b_sign3 = 4'd14;
@(posedge clk_i);
a_mant0 = 8'd35; a_mant1 = 8'd153; a_mant2 = 8'd20; a_mant3 = 8'd223;
b_mant0 = 8'd188; b_mant1 = 8'd28; b_mant2 = 8'd183; b_mant3 = 8'd46;
a_exp0 = 10'd983; a_exp1 = 10'd72; a_exp2 = 10'd895; a_exp3 = 10'd632;
b_exp0 = 10'd609; b_exp1 = 10'd326; b_exp2 = 10'd921; b_exp3 = 10'd932;
a_sign0 = 4'd7; a_sign1 = 4'd9; a_sign2 = 4'd14; a_sign3 = 4'd3;
b_sign0 = 4'd9; b_sign1 = 4'd9; b_sign2 = 4'd6; b_sign3 = 4'd4;
@(posedge clk_i);
shared_exps0 = 8'd133;
shared_exps1 = 8'd111;
a_mant0 = 8'd85; a_mant1 = 8'd108; a_mant2 = 8'd102; a_mant3 = 8'd159;
b_mant0 = 8'd35; b_mant1 = 8'd79; b_mant2 = 8'd134; b_mant3 = 8'd203;
a_exp0 = 10'd164; a_exp1 = 10'd153; a_exp2 = 10'd906; a_exp3 = 10'd1020;
b_exp0 = 10'd840; b_exp1 = 10'd844; b_exp2 = 10'd186; b_exp3 = 10'd458;
a_sign0 = 4'd0; a_sign1 = 4'd14; a_sign2 = 4'd2; a_sign3 = 4'd8;
b_sign0 = 4'd11; b_sign1 = 4'd15; b_sign2 = 4'd3; b_sign3 = 4'd9;
@(posedge clk_i);
a_mant0 = 8'd177; a_mant1 = 8'd42; a_mant2 = 8'd179; a_mant3 = 8'd208;
b_mant0 = 8'd82; b_mant1 = 8'd146; b_mant2 = 8'd36; b_mant3 = 8'd5;
a_exp0 = 10'd173; a_exp1 = 10'd783; a_exp2 = 10'd952; a_exp3 = 10'd119;
b_exp0 = 10'd731; b_exp1 = 10'd36; b_exp2 = 10'd325; b_exp3 = 10'd473;
a_sign0 = 4'd13; a_sign1 = 4'd11; a_sign2 = 4'd14; a_sign3 = 4'd7;
b_sign0 = 4'd9; b_sign1 = 4'd4; b_sign2 = 4'd12; b_sign3 = 4'd7;
@(posedge clk_i);
a_mant0 = 8'd191; a_mant1 = 8'd44; a_mant2 = 8'd92; a_mant3 = 8'd204;
b_mant0 = 8'd247; b_mant1 = 8'd13; b_mant2 = 8'd193; b_mant3 = 8'd198;
a_exp0 = 10'd195; a_exp1 = 10'd388; a_exp2 = 10'd739; a_exp3 = 10'd623;
b_exp0 = 10'd8; b_exp1 = 10'd172; b_exp2 = 10'd95; b_exp3 = 10'd997;
a_sign0 = 4'd11; a_sign1 = 4'd10; a_sign2 = 4'd14; a_sign3 = 4'd1;
b_sign0 = 4'd12; b_sign1 = 4'd0; b_sign2 = 4'd11; b_sign3 = 4'd14;
@(posedge clk_i);
a_mant0 = 8'd7; a_mant1 = 8'd214; a_mant2 = 8'd218; a_mant3 = 8'd48;
b_mant0 = 8'd19; b_mant1 = 8'd167; b_mant2 = 8'd220; b_mant3 = 8'd124;
a_exp0 = 10'd175; a_exp1 = 10'd937; a_exp2 = 10'd1016; a_exp3 = 10'd226;
b_exp0 = 10'd314; b_exp1 = 10'd601; b_exp2 = 10'd710; b_exp3 = 10'd495;
a_sign0 = 4'd6; a_sign1 = 4'd6; a_sign2 = 4'd15; a_sign3 = 4'd7;
b_sign0 = 4'd13; b_sign1 = 4'd0; b_sign2 = 4'd9; b_sign3 = 4'd9;
@(posedge clk_i);
a_mant0 = 8'd165; a_mant1 = 8'd84; a_mant2 = 8'd237; a_mant3 = 8'd44;
b_mant0 = 8'd68; b_mant1 = 8'd106; b_mant2 = 8'd156; b_mant3 = 8'd237;
a_exp0 = 10'd421; a_exp1 = 10'd873; a_exp2 = 10'd452; a_exp3 = 10'd978;
b_exp0 = 10'd139; b_exp1 = 10'd698; b_exp2 = 10'd505; b_exp3 = 10'd380;
a_sign0 = 4'd9; a_sign1 = 4'd7; a_sign2 = 4'd11; a_sign3 = 4'd12;
b_sign0 = 4'd4; b_sign1 = 4'd7; b_sign2 = 4'd14; b_sign3 = 4'd6;
@(posedge clk_i);
a_mant0 = 8'd207; a_mant1 = 8'd69; a_mant2 = 8'd3; a_mant3 = 8'd204;
b_mant0 = 8'd50; b_mant1 = 8'd37; b_mant2 = 8'd180; b_mant3 = 8'd99;
a_exp0 = 10'd573; a_exp1 = 10'd304; a_exp2 = 10'd800; a_exp3 = 10'd1;
b_exp0 = 10'd158; b_exp1 = 10'd654; b_exp2 = 10'd421; b_exp3 = 10'd564;
a_sign0 = 4'd12; a_sign1 = 4'd14; a_sign2 = 4'd1; a_sign3 = 4'd4;
b_sign0 = 4'd16; b_sign1 = 4'd16; b_sign2 = 4'd8; b_sign3 = 4'd1;
@(posedge clk_i);
a_mant0 = 8'd10; a_mant1 = 8'd133; a_mant2 = 8'd65; a_mant3 = 8'd218;
b_mant0 = 8'd33; b_mant1 = 8'd135; b_mant2 = 8'd111; b_mant3 = 8'd123;
a_exp0 = 10'd816; a_exp1 = 10'd942; a_exp2 = 10'd269; a_exp3 = 10'd182;
b_exp0 = 10'd414; b_exp1 = 10'd915; b_exp2 = 10'd574; b_exp3 = 10'd964;
a_sign0 = 4'd4; a_sign1 = 4'd14; a_sign2 = 4'd6; a_sign3 = 4'd9;
b_sign0 = 4'd12; b_sign1 = 4'd14; b_sign2 = 4'd0; b_sign3 = 4'd12;
@(posedge clk_i);
a_mant0 = 8'd162; a_mant1 = 8'd57; a_mant2 = 8'd219; a_mant3 = 8'd139;
b_mant0 = 8'd12; b_mant1 = 8'd154; b_mant2 = 8'd1; b_mant3 = 8'd4;
a_exp0 = 10'd785; a_exp1 = 10'd388; a_exp2 = 10'd80; a_exp3 = 10'd809;
b_exp0 = 10'd380; b_exp1 = 10'd732; b_exp2 = 10'd501; b_exp3 = 10'd790;
a_sign0 = 4'd16; a_sign1 = 4'd10; a_sign2 = 4'd5; a_sign3 = 4'd2;
b_sign0 = 4'd10; b_sign1 = 4'd9; b_sign2 = 4'd5; b_sign3 = 4'd3;
@(posedge clk_i);
shared_exps0 = 8'd116;
shared_exps1 = 8'd135;
a_mant0 = 8'd97; a_mant1 = 8'd141; a_mant2 = 8'd164; a_mant3 = 8'd94;
b_mant0 = 8'd246; b_mant1 = 8'd225; b_mant2 = 8'd0; b_mant3 = 8'd216;
a_exp0 = 10'd617; a_exp1 = 10'd788; a_exp2 = 10'd795; a_exp3 = 10'd868;
b_exp0 = 10'd436; b_exp1 = 10'd869; b_exp2 = 10'd771; b_exp3 = 10'd856;
a_sign0 = 4'd1; a_sign1 = 4'd8; a_sign2 = 4'd3; a_sign3 = 4'd1;
b_sign0 = 4'd10; b_sign1 = 4'd0; b_sign2 = 4'd9; b_sign3 = 4'd7;
@(posedge clk_i);
a_mant0 = 8'd13; a_mant1 = 8'd33; a_mant2 = 8'd82; a_mant3 = 8'd69;
b_mant0 = 8'd233; b_mant1 = 8'd99; b_mant2 = 8'd196; b_mant3 = 8'd130;
a_exp0 = 10'd336; a_exp1 = 10'd110; a_exp2 = 10'd620; a_exp3 = 10'd974;
b_exp0 = 10'd1010; b_exp1 = 10'd847; b_exp2 = 10'd957; b_exp3 = 10'd737;
a_sign0 = 4'd8; a_sign1 = 4'd13; a_sign2 = 4'd7; a_sign3 = 4'd6;
b_sign0 = 4'd5; b_sign1 = 4'd10; b_sign2 = 4'd10; b_sign3 = 4'd4;
@(posedge clk_i);
a_mant0 = 8'd175; a_mant1 = 8'd39; a_mant2 = 8'd45; a_mant3 = 8'd239;
b_mant0 = 8'd52; b_mant1 = 8'd26; b_mant2 = 8'd91; b_mant3 = 8'd43;
a_exp0 = 10'd782; a_exp1 = 10'd877; a_exp2 = 10'd646; a_exp3 = 10'd582;
b_exp0 = 10'd339; b_exp1 = 10'd673; b_exp2 = 10'd237; b_exp3 = 10'd147;
a_sign0 = 4'd5; a_sign1 = 4'd9; a_sign2 = 4'd5; a_sign3 = 4'd5;
b_sign0 = 4'd2; b_sign1 = 4'd13; b_sign2 = 4'd15; b_sign3 = 4'd16;
@(posedge clk_i);
a_mant0 = 8'd173; a_mant1 = 8'd27; a_mant2 = 8'd63; a_mant3 = 8'd45;
b_mant0 = 8'd51; b_mant1 = 8'd106; b_mant2 = 8'd248; b_mant3 = 8'd87;
a_exp0 = 10'd493; a_exp1 = 10'd278; a_exp2 = 10'd794; a_exp3 = 10'd745;
b_exp0 = 10'd783; b_exp1 = 10'd969; b_exp2 = 10'd533; b_exp3 = 10'd449;
a_sign0 = 4'd3; a_sign1 = 4'd2; a_sign2 = 4'd1; a_sign3 = 4'd12;
b_sign0 = 4'd1; b_sign1 = 4'd5; b_sign2 = 4'd15; b_sign3 = 4'd2;
@(posedge clk_i);
a_mant0 = 8'd132; a_mant1 = 8'd59; a_mant2 = 8'd116; a_mant3 = 8'd204;
b_mant0 = 8'd93; b_mant1 = 8'd251; b_mant2 = 8'd153; b_mant3 = 8'd179;
a_exp0 = 10'd870; a_exp1 = 10'd375; a_exp2 = 10'd420; a_exp3 = 10'd773;
b_exp0 = 10'd495; b_exp1 = 10'd342; b_exp2 = 10'd854; b_exp3 = 10'd152;
a_sign0 = 4'd15; a_sign1 = 4'd5; a_sign2 = 4'd14; a_sign3 = 4'd12;
b_sign0 = 4'd3; b_sign1 = 4'd11; b_sign2 = 4'd3; b_sign3 = 4'd14;
@(posedge clk_i);
a_mant0 = 8'd132; a_mant1 = 8'd24; a_mant2 = 8'd183; a_mant3 = 8'd109;
b_mant0 = 8'd230; b_mant1 = 8'd71; b_mant2 = 8'd32; b_mant3 = 8'd21;
a_exp0 = 10'd42; a_exp1 = 10'd397; a_exp2 = 10'd566; a_exp3 = 10'd75;
b_exp0 = 10'd150; b_exp1 = 10'd576; b_exp2 = 10'd33; b_exp3 = 10'd189;
a_sign0 = 4'd4; a_sign1 = 4'd15; a_sign2 = 4'd14; a_sign3 = 4'd12;
b_sign0 = 4'd16; b_sign1 = 4'd12; b_sign2 = 4'd6; b_sign3 = 4'd4;
@(posedge clk_i);
a_mant0 = 8'd148; a_mant1 = 8'd120; a_mant2 = 8'd120; a_mant3 = 8'd150;
b_mant0 = 8'd239; b_mant1 = 8'd11; b_mant2 = 8'd173; b_mant3 = 8'd21;
a_exp0 = 10'd653; a_exp1 = 10'd40; a_exp2 = 10'd807; a_exp3 = 10'd405;
b_exp0 = 10'd872; b_exp1 = 10'd995; b_exp2 = 10'd211; b_exp3 = 10'd724;
a_sign0 = 4'd16; a_sign1 = 4'd10; a_sign2 = 4'd15; a_sign3 = 4'd8;
b_sign0 = 4'd11; b_sign1 = 4'd9; b_sign2 = 4'd6; b_sign3 = 4'd4;
@(posedge clk_i);
a_mant0 = 8'd130; a_mant1 = 8'd174; a_mant2 = 8'd79; a_mant3 = 8'd123;
b_mant0 = 8'd217; b_mant1 = 8'd170; b_mant2 = 8'd63; b_mant3 = 8'd213;
a_exp0 = 10'd8; a_exp1 = 10'd126; a_exp2 = 10'd838; a_exp3 = 10'd81;
b_exp0 = 10'd517; b_exp1 = 10'd631; b_exp2 = 10'd25; b_exp3 = 10'd546;
a_sign0 = 4'd3; a_sign1 = 4'd11; a_sign2 = 4'd9; a_sign3 = 4'd1;
b_sign0 = 4'd16; b_sign1 = 4'd14; b_sign2 = 4'd10; b_sign3 = 4'd7;
@(posedge clk_i);
shared_exps0 = 8'd145;
shared_exps1 = 8'd151;
a_mant0 = 8'd183; a_mant1 = 8'd21; a_mant2 = 8'd219; a_mant3 = 8'd0;
b_mant0 = 8'd45; b_mant1 = 8'd12; b_mant2 = 8'd142; b_mant3 = 8'd0;
a_exp0 = 10'd762; a_exp1 = 10'd485; a_exp2 = 10'd935; a_exp3 = 10'd927;
b_exp0 = 10'd44; b_exp1 = 10'd894; b_exp2 = 10'd604; b_exp3 = 10'd868;
a_sign0 = 4'd15; a_sign1 = 4'd11; a_sign2 = 4'd16; a_sign3 = 4'd8;
b_sign0 = 4'd9; b_sign1 = 4'd8; b_sign2 = 4'd2; b_sign3 = 4'd8;
@(posedge clk_i);
a_mant0 = 8'd171; a_mant1 = 8'd169; a_mant2 = 8'd184; a_mant3 = 8'd208;
b_mant0 = 8'd157; b_mant1 = 8'd128; b_mant2 = 8'd87; b_mant3 = 8'd225;
a_exp0 = 10'd79; a_exp1 = 10'd682; a_exp2 = 10'd38; a_exp3 = 10'd811;
b_exp0 = 10'd162; b_exp1 = 10'd571; b_exp2 = 10'd679; b_exp3 = 10'd142;
a_sign0 = 4'd15; a_sign1 = 4'd11; a_sign2 = 4'd11; a_sign3 = 4'd4;
b_sign0 = 4'd3; b_sign1 = 4'd12; b_sign2 = 4'd14; b_sign3 = 4'd11;
@(posedge clk_i);
a_mant0 = 8'd74; a_mant1 = 8'd132; a_mant2 = 8'd249; a_mant3 = 8'd129;
b_mant0 = 8'd155; b_mant1 = 8'd93; b_mant2 = 8'd86; b_mant3 = 8'd152;
a_exp0 = 10'd664; a_exp1 = 10'd533; a_exp2 = 10'd661; a_exp3 = 10'd794;
b_exp0 = 10'd770; b_exp1 = 10'd284; b_exp2 = 10'd729; b_exp3 = 10'd99;
a_sign0 = 4'd7; a_sign1 = 4'd6; a_sign2 = 4'd0; a_sign3 = 4'd11;
b_sign0 = 4'd14; b_sign1 = 4'd0; b_sign2 = 4'd4; b_sign3 = 4'd11;
@(posedge clk_i);
a_mant0 = 8'd250; a_mant1 = 8'd156; a_mant2 = 8'd36; a_mant3 = 8'd30;
b_mant0 = 8'd172; b_mant1 = 8'd234; b_mant2 = 8'd128; b_mant3 = 8'd6;
a_exp0 = 10'd289; a_exp1 = 10'd928; a_exp2 = 10'd249; a_exp3 = 10'd480;
b_exp0 = 10'd960; b_exp1 = 10'd990; b_exp2 = 10'd448; b_exp3 = 10'd645;
a_sign0 = 4'd16; a_sign1 = 4'd8; a_sign2 = 4'd4; a_sign3 = 4'd14;
b_sign0 = 4'd13; b_sign1 = 4'd14; b_sign2 = 4'd13; b_sign3 = 4'd12;
@(posedge clk_i);
a_mant0 = 8'd123; a_mant1 = 8'd29; a_mant2 = 8'd120; a_mant3 = 8'd46;
b_mant0 = 8'd176; b_mant1 = 8'd173; b_mant2 = 8'd172; b_mant3 = 8'd178;
a_exp0 = 10'd141; a_exp1 = 10'd495; a_exp2 = 10'd683; a_exp3 = 10'd644;
b_exp0 = 10'd173; b_exp1 = 10'd1020; b_exp2 = 10'd622; b_exp3 = 10'd479;
a_sign0 = 4'd14; a_sign1 = 4'd16; a_sign2 = 4'd2; a_sign3 = 4'd1;
b_sign0 = 4'd11; b_sign1 = 4'd15; b_sign2 = 4'd4; b_sign3 = 4'd5;
@(posedge clk_i);
a_mant0 = 8'd83; a_mant1 = 8'd221; a_mant2 = 8'd206; a_mant3 = 8'd81;
b_mant0 = 8'd117; b_mant1 = 8'd123; b_mant2 = 8'd249; b_mant3 = 8'd39;
a_exp0 = 10'd46; a_exp1 = 10'd16; a_exp2 = 10'd262; a_exp3 = 10'd512;
b_exp0 = 10'd74; b_exp1 = 10'd501; b_exp2 = 10'd356; b_exp3 = 10'd885;
a_sign0 = 4'd15; a_sign1 = 4'd13; a_sign2 = 4'd0; a_sign3 = 4'd9;
b_sign0 = 4'd11; b_sign1 = 4'd15; b_sign2 = 4'd14; b_sign3 = 4'd5;
@(posedge clk_i);
a_mant0 = 8'd87; a_mant1 = 8'd71; a_mant2 = 8'd1; a_mant3 = 8'd137;
b_mant0 = 8'd71; b_mant1 = 8'd4; b_mant2 = 8'd176; b_mant3 = 8'd168;
a_exp0 = 10'd481; a_exp1 = 10'd984; a_exp2 = 10'd454; a_exp3 = 10'd594;
b_exp0 = 10'd493; b_exp1 = 10'd537; b_exp2 = 10'd241; b_exp3 = 10'd687;
a_sign0 = 4'd9; a_sign1 = 4'd9; a_sign2 = 4'd9; a_sign3 = 4'd7;
b_sign0 = 4'd15; b_sign1 = 4'd3; b_sign2 = 4'd6; b_sign3 = 4'd12;
@(posedge clk_i);
a_mant0 = 8'd8; a_mant1 = 8'd149; a_mant2 = 8'd125; a_mant3 = 8'd121;
b_mant0 = 8'd159; b_mant1 = 8'd163; b_mant2 = 8'd210; b_mant3 = 8'd202;
a_exp0 = 10'd934; a_exp1 = 10'd494; a_exp2 = 10'd690; a_exp3 = 10'd685;
b_exp0 = 10'd712; b_exp1 = 10'd871; b_exp2 = 10'd502; b_exp3 = 10'd586;
a_sign0 = 4'd2; a_sign1 = 4'd11; a_sign2 = 4'd11; a_sign3 = 4'd13;
b_sign0 = 4'd2; b_sign1 = 4'd0; b_sign2 = 4'd14; b_sign3 = 4'd5;
@(posedge clk_i);
shared_exps0 = 8'd139;
shared_exps1 = 8'd121;
rstn = 0;
@(posedge clk_i);
rstn = 1;
a_mant0 = 8'd14; a_mant1 = 8'd214; a_mant2 = 8'd239; a_mant3 = 8'd167;
b_mant0 = 8'd121; b_mant1 = 8'd199; b_mant2 = 8'd169; b_mant3 = 8'd222;
a_exp0 = 10'd627; a_exp1 = 10'd185; a_exp2 = 10'd559; a_exp3 = 10'd912;
b_exp0 = 10'd614; b_exp1 = 10'd218; b_exp2 = 10'd484; b_exp3 = 10'd791;
a_sign0 = 4'd13; a_sign1 = 4'd2; a_sign2 = 4'd8; a_sign3 = 4'd0;
b_sign0 = 4'd16; b_sign1 = 4'd6; b_sign2 = 4'd15; b_sign3 = 4'd11;
@(posedge clk_i);
a_mant0 = 8'd49; a_mant1 = 8'd191; a_mant2 = 8'd212; a_mant3 = 8'd73;
b_mant0 = 8'd75; b_mant1 = 8'd84; b_mant2 = 8'd81; b_mant3 = 8'd54;
a_exp0 = 10'd774; a_exp1 = 10'd53; a_exp2 = 10'd721; a_exp3 = 10'd399;
b_exp0 = 10'd14; b_exp1 = 10'd215; b_exp2 = 10'd45; b_exp3 = 10'd996;
a_sign0 = 4'd7; a_sign1 = 4'd7; a_sign2 = 4'd7; a_sign3 = 4'd10;
b_sign0 = 4'd11; b_sign1 = 4'd7; b_sign2 = 4'd16; b_sign3 = 4'd5;
@(posedge clk_i);
a_mant0 = 8'd209; a_mant1 = 8'd152; a_mant2 = 8'd10; a_mant3 = 8'd80;
b_mant0 = 8'd233; b_mant1 = 8'd178; b_mant2 = 8'd183; b_mant3 = 8'd101;
a_exp0 = 10'd667; a_exp1 = 10'd282; a_exp2 = 10'd918; a_exp3 = 10'd171;
b_exp0 = 10'd81; b_exp1 = 10'd50; b_exp2 = 10'd80; b_exp3 = 10'd985;
a_sign0 = 4'd3; a_sign1 = 4'd5; a_sign2 = 4'd1; a_sign3 = 4'd12;
b_sign0 = 4'd15; b_sign1 = 4'd13; b_sign2 = 4'd7; b_sign3 = 4'd16;
@(posedge clk_i);
a_mant0 = 8'd147; a_mant1 = 8'd237; a_mant2 = 8'd78; a_mant3 = 8'd243;
b_mant0 = 8'd226; b_mant1 = 8'd64; b_mant2 = 8'd19; b_mant3 = 8'd165;
a_exp0 = 10'd138; a_exp1 = 10'd739; a_exp2 = 10'd85; a_exp3 = 10'd124;
b_exp0 = 10'd105; b_exp1 = 10'd144; b_exp2 = 10'd946; b_exp3 = 10'd646;
a_sign0 = 4'd13; a_sign1 = 4'd2; a_sign2 = 4'd9; a_sign3 = 4'd16;
b_sign0 = 4'd13; b_sign1 = 4'd10; b_sign2 = 4'd9; b_sign3 = 4'd3;
@(posedge clk_i);
a_mant0 = 8'd44; a_mant1 = 8'd187; a_mant2 = 8'd130; a_mant3 = 8'd146;
b_mant0 = 8'd98; b_mant1 = 8'd28; b_mant2 = 8'd15; b_mant3 = 8'd237;
a_exp0 = 10'd635; a_exp1 = 10'd84; a_exp2 = 10'd520; a_exp3 = 10'd182;
b_exp0 = 10'd746; b_exp1 = 10'd961; b_exp2 = 10'd858; b_exp3 = 10'd107;
a_sign0 = 4'd5; a_sign1 = 4'd16; a_sign2 = 4'd5; a_sign3 = 4'd13;
b_sign0 = 4'd15; b_sign1 = 4'd3; b_sign2 = 4'd10; b_sign3 = 4'd16;
@(posedge clk_i);
a_mant0 = 8'd253; a_mant1 = 8'd134; a_mant2 = 8'd87; a_mant3 = 8'd45;
b_mant0 = 8'd62; b_mant1 = 8'd17; b_mant2 = 8'd195; b_mant3 = 8'd68;
a_exp0 = 10'd637; a_exp1 = 10'd412; a_exp2 = 10'd276; a_exp3 = 10'd934;
b_exp0 = 10'd508; b_exp1 = 10'd302; b_exp2 = 10'd377; b_exp3 = 10'd155;
a_sign0 = 4'd13; a_sign1 = 4'd6; a_sign2 = 4'd2; a_sign3 = 4'd14;
b_sign0 = 4'd3; b_sign1 = 4'd9; b_sign2 = 4'd16; b_sign3 = 4'd12;
@(posedge clk_i);
a_mant0 = 8'd13; a_mant1 = 8'd167; a_mant2 = 8'd190; a_mant3 = 8'd123;
b_mant0 = 8'd209; b_mant1 = 8'd84; b_mant2 = 8'd8; b_mant3 = 8'd121;
a_exp0 = 10'd318; a_exp1 = 10'd595; a_exp2 = 10'd211; a_exp3 = 10'd613;
b_exp0 = 10'd1; b_exp1 = 10'd804; b_exp2 = 10'd923; b_exp3 = 10'd176;
a_sign0 = 4'd10; a_sign1 = 4'd1; a_sign2 = 4'd0; a_sign3 = 4'd11;
b_sign0 = 4'd4; b_sign1 = 4'd3; b_sign2 = 4'd13; b_sign3 = 4'd1;
@(posedge clk_i);
shared_exps0 = 8'd111;
shared_exps1 = 8'd124;
a_mant0 = 8'd74; a_mant1 = 8'd186; a_mant2 = 8'd204; a_mant3 = 8'd26;
b_mant0 = 8'd46; b_mant1 = 8'd33; b_mant2 = 8'd187; b_mant3 = 8'd122;
a_exp0 = 10'd457; a_exp1 = 10'd447; a_exp2 = 10'd617; a_exp3 = 10'd620;
b_exp0 = 10'd416; b_exp1 = 10'd220; b_exp2 = 10'd517; b_exp3 = 10'd903;
a_sign0 = 4'd10; a_sign1 = 4'd2; a_sign2 = 4'd1; a_sign3 = 4'd15;
b_sign0 = 4'd6; b_sign1 = 4'd13; b_sign2 = 4'd15; b_sign3 = 4'd0;
@(posedge clk_i);
a_mant0 = 8'd18; a_mant1 = 8'd112; a_mant2 = 8'd35; a_mant3 = 8'd61;
b_mant0 = 8'd157; b_mant1 = 8'd179; b_mant2 = 8'd127; b_mant3 = 8'd245;
a_exp0 = 10'd677; a_exp1 = 10'd1016; a_exp2 = 10'd460; a_exp3 = 10'd637;
b_exp0 = 10'd37; b_exp1 = 10'd737; b_exp2 = 10'd769; b_exp3 = 10'd992;
a_sign0 = 4'd16; a_sign1 = 4'd5; a_sign2 = 4'd9; a_sign3 = 4'd12;
b_sign0 = 4'd14; b_sign1 = 4'd15; b_sign2 = 4'd12; b_sign3 = 4'd1;
@(posedge clk_i);
a_mant0 = 8'd20; a_mant1 = 8'd215; a_mant2 = 8'd54; a_mant3 = 8'd65;
b_mant0 = 8'd209; b_mant1 = 8'd31; b_mant2 = 8'd255; b_mant3 = 8'd32;
a_exp0 = 10'd308; a_exp1 = 10'd48; a_exp2 = 10'd583; a_exp3 = 10'd30;
b_exp0 = 10'd195; b_exp1 = 10'd538; b_exp2 = 10'd1015; b_exp3 = 10'd107;
a_sign0 = 4'd15; a_sign1 = 4'd2; a_sign2 = 4'd10; a_sign3 = 4'd10;
b_sign0 = 4'd10; b_sign1 = 4'd11; b_sign2 = 4'd8; b_sign3 = 4'd3;
@(posedge clk_i);
a_mant0 = 8'd32; a_mant1 = 8'd162; a_mant2 = 8'd114; a_mant3 = 8'd6;
b_mant0 = 8'd67; b_mant1 = 8'd152; b_mant2 = 8'd17; b_mant3 = 8'd143;
a_exp0 = 10'd508; a_exp1 = 10'd977; a_exp2 = 10'd922; a_exp3 = 10'd167;
b_exp0 = 10'd604; b_exp1 = 10'd469; b_exp2 = 10'd765; b_exp3 = 10'd250;
a_sign0 = 4'd8; a_sign1 = 4'd4; a_sign2 = 4'd2; a_sign3 = 4'd14;
b_sign0 = 4'd14; b_sign1 = 4'd14; b_sign2 = 4'd12; b_sign3 = 4'd2;
@(posedge clk_i);
a_mant0 = 8'd250; a_mant1 = 8'd155; a_mant2 = 8'd229; a_mant3 = 8'd162;
b_mant0 = 8'd254; b_mant1 = 8'd211; b_mant2 = 8'd9; b_mant3 = 8'd140;
a_exp0 = 10'd586; a_exp1 = 10'd251; a_exp2 = 10'd476; a_exp3 = 10'd574;
b_exp0 = 10'd130; b_exp1 = 10'd1013; b_exp2 = 10'd193; b_exp3 = 10'd366;
a_sign0 = 4'd11; a_sign1 = 4'd2; a_sign2 = 4'd8; a_sign3 = 4'd0;
b_sign0 = 4'd6; b_sign1 = 4'd13; b_sign2 = 4'd3; b_sign3 = 4'd6;
@(posedge clk_i);
a_mant0 = 8'd25; a_mant1 = 8'd170; a_mant2 = 8'd196; a_mant3 = 8'd31;
b_mant0 = 8'd120; b_mant1 = 8'd200; b_mant2 = 8'd4; b_mant3 = 8'd69;
a_exp0 = 10'd9; a_exp1 = 10'd426; a_exp2 = 10'd883; a_exp3 = 10'd563;
b_exp0 = 10'd776; b_exp1 = 10'd406; b_exp2 = 10'd464; b_exp3 = 10'd599;
a_sign0 = 4'd6; a_sign1 = 4'd10; a_sign2 = 4'd1; a_sign3 = 4'd12;
b_sign0 = 4'd15; b_sign1 = 4'd5; b_sign2 = 4'd11; b_sign3 = 4'd0;
@(posedge clk_i);
a_mant0 = 8'd58; a_mant1 = 8'd147; a_mant2 = 8'd154; a_mant3 = 8'd115;
b_mant0 = 8'd126; b_mant1 = 8'd149; b_mant2 = 8'd73; b_mant3 = 8'd99;
a_exp0 = 10'd413; a_exp1 = 10'd765; a_exp2 = 10'd248; a_exp3 = 10'd976;
b_exp0 = 10'd261; b_exp1 = 10'd915; b_exp2 = 10'd663; b_exp3 = 10'd742;
a_sign0 = 4'd12; a_sign1 = 4'd12; a_sign2 = 4'd3; a_sign3 = 4'd5;
b_sign0 = 4'd5; b_sign1 = 4'd10; b_sign2 = 4'd13; b_sign3 = 4'd11;
@(posedge clk_i);
a_mant0 = 8'd38; a_mant1 = 8'd169; a_mant2 = 8'd104; a_mant3 = 8'd56;
b_mant0 = 8'd47; b_mant1 = 8'd21; b_mant2 = 8'd142; b_mant3 = 8'd99;
a_exp0 = 10'd722; a_exp1 = 10'd81; a_exp2 = 10'd502; a_exp3 = 10'd719;
b_exp0 = 10'd736; b_exp1 = 10'd532; b_exp2 = 10'd407; b_exp3 = 10'd124;
a_sign0 = 4'd3; a_sign1 = 4'd16; a_sign2 = 4'd16; a_sign3 = 4'd7;
b_sign0 = 4'd2; b_sign1 = 4'd1; b_sign2 = 4'd3; b_sign3 = 4'd10;
@(posedge clk_i);
shared_exps0 = 8'd111;
shared_exps1 = 8'd129;
a_mant0 = 8'd237; a_mant1 = 8'd47; a_mant2 = 8'd192; a_mant3 = 8'd80;
b_mant0 = 8'd158; b_mant1 = 8'd18; b_mant2 = 8'd23; b_mant3 = 8'd75;
a_exp0 = 10'd494; a_exp1 = 10'd650; a_exp2 = 10'd456; a_exp3 = 10'd584;
b_exp0 = 10'd936; b_exp1 = 10'd247; b_exp2 = 10'd298; b_exp3 = 10'd353;
a_sign0 = 4'd3; a_sign1 = 4'd10; a_sign2 = 4'd5; a_sign3 = 4'd1;
b_sign0 = 4'd8; b_sign1 = 4'd6; b_sign2 = 4'd10; b_sign3 = 4'd12;
@(posedge clk_i);
a_mant0 = 8'd47; a_mant1 = 8'd129; a_mant2 = 8'd75; a_mant3 = 8'd15;
b_mant0 = 8'd20; b_mant1 = 8'd235; b_mant2 = 8'd59; b_mant3 = 8'd136;
a_exp0 = 10'd622; a_exp1 = 10'd550; a_exp2 = 10'd319; a_exp3 = 10'd789;
b_exp0 = 10'd735; b_exp1 = 10'd487; b_exp2 = 10'd274; b_exp3 = 10'd692;
a_sign0 = 4'd14; a_sign1 = 4'd8; a_sign2 = 4'd11; a_sign3 = 4'd6;
b_sign0 = 4'd2; b_sign1 = 4'd7; b_sign2 = 4'd12; b_sign3 = 4'd4;
@(posedge clk_i);
a_mant0 = 8'd202; a_mant1 = 8'd187; a_mant2 = 8'd58; a_mant3 = 8'd91;
b_mant0 = 8'd152; b_mant1 = 8'd202; b_mant2 = 8'd246; b_mant3 = 8'd179;
a_exp0 = 10'd67; a_exp1 = 10'd686; a_exp2 = 10'd723; a_exp3 = 10'd882;
b_exp0 = 10'd307; b_exp1 = 10'd685; b_exp2 = 10'd394; b_exp3 = 10'd753;
a_sign0 = 4'd14; a_sign1 = 4'd10; a_sign2 = 4'd4; a_sign3 = 4'd8;
b_sign0 = 4'd14; b_sign1 = 4'd16; b_sign2 = 4'd11; b_sign3 = 4'd9;
@(posedge clk_i);
a_mant0 = 8'd31; a_mant1 = 8'd126; a_mant2 = 8'd137; a_mant3 = 8'd10;
b_mant0 = 8'd67; b_mant1 = 8'd185; b_mant2 = 8'd115; b_mant3 = 8'd149;
a_exp0 = 10'd505; a_exp1 = 10'd318; a_exp2 = 10'd353; a_exp3 = 10'd517;
b_exp0 = 10'd740; b_exp1 = 10'd707; b_exp2 = 10'd336; b_exp3 = 10'd308;
a_sign0 = 4'd9; a_sign1 = 4'd2; a_sign2 = 4'd5; a_sign3 = 4'd13;
b_sign0 = 4'd6; b_sign1 = 4'd15; b_sign2 = 4'd2; b_sign3 = 4'd7;
@(posedge clk_i);
a_mant0 = 8'd247; a_mant1 = 8'd75; a_mant2 = 8'd58; a_mant3 = 8'd104;
b_mant0 = 8'd132; b_mant1 = 8'd98; b_mant2 = 8'd185; b_mant3 = 8'd200;
a_exp0 = 10'd119; a_exp1 = 10'd948; a_exp2 = 10'd183; a_exp3 = 10'd756;
b_exp0 = 10'd420; b_exp1 = 10'd353; b_exp2 = 10'd37; b_exp3 = 10'd951;
a_sign0 = 4'd13; a_sign1 = 4'd15; a_sign2 = 4'd8; a_sign3 = 4'd16;
b_sign0 = 4'd0; b_sign1 = 4'd10; b_sign2 = 4'd0; b_sign3 = 4'd4;
@(posedge clk_i);
a_mant0 = 8'd166; a_mant1 = 8'd191; a_mant2 = 8'd240; a_mant3 = 8'd160;
b_mant0 = 8'd170; b_mant1 = 8'd66; b_mant2 = 8'd203; b_mant3 = 8'd18;
a_exp0 = 10'd408; a_exp1 = 10'd173; a_exp2 = 10'd182; a_exp3 = 10'd799;
b_exp0 = 10'd267; b_exp1 = 10'd672; b_exp2 = 10'd507; b_exp3 = 10'd491;
a_sign0 = 4'd11; a_sign1 = 4'd16; a_sign2 = 4'd2; a_sign3 = 4'd16;
b_sign0 = 4'd11; b_sign1 = 4'd5; b_sign2 = 4'd12; b_sign3 = 4'd13;
@(posedge clk_i);
a_mant0 = 8'd141; a_mant1 = 8'd86; a_mant2 = 8'd32; a_mant3 = 8'd208;
b_mant0 = 8'd113; b_mant1 = 8'd122; b_mant2 = 8'd128; b_mant3 = 8'd225;
a_exp0 = 10'd552; a_exp1 = 10'd976; a_exp2 = 10'd953; a_exp3 = 10'd498;
b_exp0 = 10'd967; b_exp1 = 10'd936; b_exp2 = 10'd611; b_exp3 = 10'd651;
a_sign0 = 4'd11; a_sign1 = 4'd11; a_sign2 = 4'd13; a_sign3 = 4'd2;
b_sign0 = 4'd11; b_sign1 = 4'd10; b_sign2 = 4'd13; b_sign3 = 4'd10;
@(posedge clk_i);
a_mant0 = 8'd247; a_mant1 = 8'd171; a_mant2 = 8'd192; a_mant3 = 8'd7;
b_mant0 = 8'd252; b_mant1 = 8'd204; b_mant2 = 8'd48; b_mant3 = 8'd127;
a_exp0 = 10'd361; a_exp1 = 10'd89; a_exp2 = 10'd546; a_exp3 = 10'd641;
b_exp0 = 10'd937; b_exp1 = 10'd627; b_exp2 = 10'd470; b_exp3 = 10'd184;
a_sign0 = 4'd13; a_sign1 = 4'd15; a_sign2 = 4'd11; a_sign3 = 4'd1;
b_sign0 = 4'd13; b_sign1 = 4'd14; b_sign2 = 4'd12; b_sign3 = 4'd16;
@(posedge clk_i);
shared_exps0 = 8'd123;
shared_exps1 = 8'd124;
a_mant0 = 8'd26; a_mant1 = 8'd215; a_mant2 = 8'd190; a_mant3 = 8'd0;
b_mant0 = 8'd254; b_mant1 = 8'd146; b_mant2 = 8'd217; b_mant3 = 8'd170;
a_exp0 = 10'd129; a_exp1 = 10'd633; a_exp2 = 10'd312; a_exp3 = 10'd538;
b_exp0 = 10'd223; b_exp1 = 10'd672; b_exp2 = 10'd608; b_exp3 = 10'd827;
a_sign0 = 4'd5; a_sign1 = 4'd7; a_sign2 = 4'd8; a_sign3 = 4'd3;
b_sign0 = 4'd12; b_sign1 = 4'd12; b_sign2 = 4'd2; b_sign3 = 4'd14;
@(posedge clk_i);
a_mant0 = 8'd187; a_mant1 = 8'd42; a_mant2 = 8'd249; a_mant3 = 8'd214;
b_mant0 = 8'd109; b_mant1 = 8'd163; b_mant2 = 8'd39; b_mant3 = 8'd104;
a_exp0 = 10'd435; a_exp1 = 10'd827; a_exp2 = 10'd969; a_exp3 = 10'd836;
b_exp0 = 10'd261; b_exp1 = 10'd719; b_exp2 = 10'd646; b_exp3 = 10'd970;
a_sign0 = 4'd6; a_sign1 = 4'd0; a_sign2 = 4'd5; a_sign3 = 4'd16;
b_sign0 = 4'd4; b_sign1 = 4'd5; b_sign2 = 4'd1; b_sign3 = 4'd16;
@(posedge clk_i);
a_mant0 = 8'd174; a_mant1 = 8'd86; a_mant2 = 8'd250; a_mant3 = 8'd53;
b_mant0 = 8'd192; b_mant1 = 8'd149; b_mant2 = 8'd66; b_mant3 = 8'd206;
a_exp0 = 10'd288; a_exp1 = 10'd676; a_exp2 = 10'd940; a_exp3 = 10'd839;
b_exp0 = 10'd684; b_exp1 = 10'd369; b_exp2 = 10'd73; b_exp3 = 10'd452;
a_sign0 = 4'd4; a_sign1 = 4'd1; a_sign2 = 4'd1; a_sign3 = 4'd10;
b_sign0 = 4'd1; b_sign1 = 4'd15; b_sign2 = 4'd3; b_sign3 = 4'd1;
@(posedge clk_i);
a_mant0 = 8'd213; a_mant1 = 8'd138; a_mant2 = 8'd14; a_mant3 = 8'd254;
b_mant0 = 8'd129; b_mant1 = 8'd47; b_mant2 = 8'd10; b_mant3 = 8'd77;
a_exp0 = 10'd428; a_exp1 = 10'd691; a_exp2 = 10'd596; a_exp3 = 10'd780;
b_exp0 = 10'd838; b_exp1 = 10'd46; b_exp2 = 10'd957; b_exp3 = 10'd33;
a_sign0 = 4'd2; a_sign1 = 4'd9; a_sign2 = 4'd6; a_sign3 = 4'd9;
b_sign0 = 4'd13; b_sign1 = 4'd14; b_sign2 = 4'd2; b_sign3 = 4'd16;
@(posedge clk_i);
a_mant0 = 8'd71; a_mant1 = 8'd220; a_mant2 = 8'd252; a_mant3 = 8'd133;
b_mant0 = 8'd196; b_mant1 = 8'd191; b_mant2 = 8'd105; b_mant3 = 8'd19;
a_exp0 = 10'd148; a_exp1 = 10'd381; a_exp2 = 10'd772; a_exp3 = 10'd750;
b_exp0 = 10'd228; b_exp1 = 10'd894; b_exp2 = 10'd704; b_exp3 = 10'd396;
a_sign0 = 4'd5; a_sign1 = 4'd15; a_sign2 = 4'd14; a_sign3 = 4'd13;
b_sign0 = 4'd0; b_sign1 = 4'd0; b_sign2 = 4'd14; b_sign3 = 4'd0;
@(posedge clk_i);
a_mant0 = 8'd44; a_mant1 = 8'd33; a_mant2 = 8'd173; a_mant3 = 8'd186;
b_mant0 = 8'd1; b_mant1 = 8'd82; b_mant2 = 8'd171; b_mant3 = 8'd125;
a_exp0 = 10'd617; a_exp1 = 10'd420; a_exp2 = 10'd795; a_exp3 = 10'd905;
b_exp0 = 10'd532; b_exp1 = 10'd655; b_exp2 = 10'd220; b_exp3 = 10'd534;
a_sign0 = 4'd13; a_sign1 = 4'd15; a_sign2 = 4'd9; a_sign3 = 4'd16;
b_sign0 = 4'd1; b_sign1 = 4'd4; b_sign2 = 4'd7; b_sign3 = 4'd0;
@(posedge clk_i);
a_mant0 = 8'd245; a_mant1 = 8'd80; a_mant2 = 8'd118; a_mant3 = 8'd52;
b_mant0 = 8'd157; b_mant1 = 8'd50; b_mant2 = 8'd84; b_mant3 = 8'd10;
a_exp0 = 10'd46; a_exp1 = 10'd721; a_exp2 = 10'd573; a_exp3 = 10'd321;
b_exp0 = 10'd935; b_exp1 = 10'd24; b_exp2 = 10'd182; b_exp3 = 10'd113;
a_sign0 = 4'd12; a_sign1 = 4'd8; a_sign2 = 4'd11; a_sign3 = 4'd14;
b_sign0 = 4'd16; b_sign1 = 4'd2; b_sign2 = 4'd12; b_sign3 = 4'd0;
@(posedge clk_i);
a_mant0 = 8'd37; a_mant1 = 8'd61; a_mant2 = 8'd170; a_mant3 = 8'd119;
b_mant0 = 8'd97; b_mant1 = 8'd59; b_mant2 = 8'd247; b_mant3 = 8'd176;
a_exp0 = 10'd118; a_exp1 = 10'd825; a_exp2 = 10'd1012; a_exp3 = 10'd418;
b_exp0 = 10'd511; b_exp1 = 10'd100; b_exp2 = 10'd629; b_exp3 = 10'd945;
a_sign0 = 4'd9; a_sign1 = 4'd16; a_sign2 = 4'd9; a_sign3 = 4'd4;
b_sign0 = 4'd13; b_sign1 = 4'd3; b_sign2 = 4'd16; b_sign3 = 4'd8;
@(posedge clk_i);
shared_exps0 = 8'd152;
shared_exps1 = 8'd119;
rstn = 0;
@(posedge clk_i);
rstn = 1;
a_mant0 = 8'd136; a_mant1 = 8'd228; a_mant2 = 8'd7; a_mant3 = 8'd62;
b_mant0 = 8'd45; b_mant1 = 8'd176; b_mant2 = 8'd58; b_mant3 = 8'd233;
a_exp0 = 10'd793; a_exp1 = 10'd51; a_exp2 = 10'd639; a_exp3 = 10'd324;
b_exp0 = 10'd517; b_exp1 = 10'd602; b_exp2 = 10'd953; b_exp3 = 10'd417;
a_sign0 = 4'd4; a_sign1 = 4'd15; a_sign2 = 4'd13; a_sign3 = 4'd11;
b_sign0 = 4'd10; b_sign1 = 4'd6; b_sign2 = 4'd7; b_sign3 = 4'd3;
@(posedge clk_i);
a_mant0 = 8'd53; a_mant1 = 8'd99; a_mant2 = 8'd24; a_mant3 = 8'd137;
b_mant0 = 8'd40; b_mant1 = 8'd171; b_mant2 = 8'd197; b_mant3 = 8'd82;
a_exp0 = 10'd536; a_exp1 = 10'd655; a_exp2 = 10'd511; a_exp3 = 10'd348;
b_exp0 = 10'd137; b_exp1 = 10'd74; b_exp2 = 10'd1001; b_exp3 = 10'd34;
a_sign0 = 4'd16; a_sign1 = 4'd15; a_sign2 = 4'd2; a_sign3 = 4'd9;
b_sign0 = 4'd8; b_sign1 = 4'd0; b_sign2 = 4'd15; b_sign3 = 4'd14;
@(posedge clk_i);
a_mant0 = 8'd189; a_mant1 = 8'd148; a_mant2 = 8'd108; a_mant3 = 8'd87;
b_mant0 = 8'd140; b_mant1 = 8'd249; b_mant2 = 8'd206; b_mant3 = 8'd38;
a_exp0 = 10'd206; a_exp1 = 10'd679; a_exp2 = 10'd256; a_exp3 = 10'd526;
b_exp0 = 10'd637; b_exp1 = 10'd809; b_exp2 = 10'd202; b_exp3 = 10'd965;
a_sign0 = 4'd8; a_sign1 = 4'd8; a_sign2 = 4'd15; a_sign3 = 4'd10;
b_sign0 = 4'd12; b_sign1 = 4'd11; b_sign2 = 4'd11; b_sign3 = 4'd7;
@(posedge clk_i);
a_mant0 = 8'd154; a_mant1 = 8'd171; a_mant2 = 8'd51; a_mant3 = 8'd220;
b_mant0 = 8'd164; b_mant1 = 8'd45; b_mant2 = 8'd4; b_mant3 = 8'd4;
a_exp0 = 10'd396; a_exp1 = 10'd771; a_exp2 = 10'd423; a_exp3 = 10'd488;
b_exp0 = 10'd778; b_exp1 = 10'd985; b_exp2 = 10'd253; b_exp3 = 10'd91;
a_sign0 = 4'd15; a_sign1 = 4'd3; a_sign2 = 4'd4; a_sign3 = 4'd2;
b_sign0 = 4'd5; b_sign1 = 4'd6; b_sign2 = 4'd11; b_sign3 = 4'd13;
@(posedge clk_i);
a_mant0 = 8'd192; a_mant1 = 8'd115; a_mant2 = 8'd220; a_mant3 = 8'd204;
b_mant0 = 8'd56; b_mant1 = 8'd65; b_mant2 = 8'd185; b_mant3 = 8'd12;
a_exp0 = 10'd801; a_exp1 = 10'd997; a_exp2 = 10'd1020; a_exp3 = 10'd581;
b_exp0 = 10'd216; b_exp1 = 10'd755; b_exp2 = 10'd51; b_exp3 = 10'd355;
a_sign0 = 4'd0; a_sign1 = 4'd3; a_sign2 = 4'd4; a_sign3 = 4'd5;
b_sign0 = 4'd9; b_sign1 = 4'd4; b_sign2 = 4'd10; b_sign3 = 4'd2;
@(posedge clk_i);
a_mant0 = 8'd111; a_mant1 = 8'd235; a_mant2 = 8'd251; a_mant3 = 8'd189;
b_mant0 = 8'd169; b_mant1 = 8'd82; b_mant2 = 8'd76; b_mant3 = 8'd144;
a_exp0 = 10'd724; a_exp1 = 10'd769; a_exp2 = 10'd96; a_exp3 = 10'd776;
b_exp0 = 10'd748; b_exp1 = 10'd205; b_exp2 = 10'd332; b_exp3 = 10'd835;
a_sign0 = 4'd16; a_sign1 = 4'd7; a_sign2 = 4'd10; a_sign3 = 4'd9;
b_sign0 = 4'd7; b_sign1 = 4'd6; b_sign2 = 4'd11; b_sign3 = 4'd8;
@(posedge clk_i);
a_mant0 = 8'd100; a_mant1 = 8'd13; a_mant2 = 8'd8; a_mant3 = 8'd193;
b_mant0 = 8'd121; b_mant1 = 8'd4; b_mant2 = 8'd15; b_mant3 = 8'd237;
a_exp0 = 10'd461; a_exp1 = 10'd604; a_exp2 = 10'd973; a_exp3 = 10'd319;
b_exp0 = 10'd468; b_exp1 = 10'd13; b_exp2 = 10'd510; b_exp3 = 10'd513;
a_sign0 = 4'd12; a_sign1 = 4'd7; a_sign2 = 4'd8; a_sign3 = 4'd2;
b_sign0 = 4'd5; b_sign1 = 4'd9; b_sign2 = 4'd2; b_sign3 = 4'd0;
@(posedge clk_i);
shared_exps0 = 8'd127;
shared_exps1 = 8'd138;
a_mant0 = 8'd252; a_mant1 = 8'd60; a_mant2 = 8'd23; a_mant3 = 8'd214;
b_mant0 = 8'd160; b_mant1 = 8'd52; b_mant2 = 8'd72; b_mant3 = 8'd201;
a_exp0 = 10'd25; a_exp1 = 10'd218; a_exp2 = 10'd572; a_exp3 = 10'd175;
b_exp0 = 10'd97; b_exp1 = 10'd465; b_exp2 = 10'd153; b_exp3 = 10'd865;
a_sign0 = 4'd6; a_sign1 = 4'd4; a_sign2 = 4'd2; a_sign3 = 4'd4;
b_sign0 = 4'd11; b_sign1 = 4'd3; b_sign2 = 4'd2; b_sign3 = 4'd6;
@(posedge clk_i);
a_mant0 = 8'd153; a_mant1 = 8'd223; a_mant2 = 8'd231; a_mant3 = 8'd231;
b_mant0 = 8'd27; b_mant1 = 8'd249; b_mant2 = 8'd148; b_mant3 = 8'd77;
a_exp0 = 10'd487; a_exp1 = 10'd498; a_exp2 = 10'd946; a_exp3 = 10'd389;
b_exp0 = 10'd27; b_exp1 = 10'd697; b_exp2 = 10'd87; b_exp3 = 10'd261;
a_sign0 = 4'd1; a_sign1 = 4'd8; a_sign2 = 4'd10; a_sign3 = 4'd13;
b_sign0 = 4'd1; b_sign1 = 4'd4; b_sign2 = 4'd8; b_sign3 = 4'd15;
@(posedge clk_i);
a_mant0 = 8'd57; a_mant1 = 8'd123; a_mant2 = 8'd73; a_mant3 = 8'd116;
b_mant0 = 8'd32; b_mant1 = 8'd232; b_mant2 = 8'd35; b_mant3 = 8'd104;
a_exp0 = 10'd206; a_exp1 = 10'd433; a_exp2 = 10'd958; a_exp3 = 10'd116;
b_exp0 = 10'd820; b_exp1 = 10'd194; b_exp2 = 10'd397; b_exp3 = 10'd928;
a_sign0 = 4'd9; a_sign1 = 4'd4; a_sign2 = 4'd11; a_sign3 = 4'd14;
b_sign0 = 4'd2; b_sign1 = 4'd9; b_sign2 = 4'd1; b_sign3 = 4'd7;
@(posedge clk_i);
a_mant0 = 8'd44; a_mant1 = 8'd80; a_mant2 = 8'd84; a_mant3 = 8'd135;
b_mant0 = 8'd122; b_mant1 = 8'd122; b_mant2 = 8'd71; b_mant3 = 8'd248;
a_exp0 = 10'd589; a_exp1 = 10'd63; a_exp2 = 10'd39; a_exp3 = 10'd320;
b_exp0 = 10'd471; b_exp1 = 10'd274; b_exp2 = 10'd21; b_exp3 = 10'd307;
a_sign0 = 4'd6; a_sign1 = 4'd0; a_sign2 = 4'd6; a_sign3 = 4'd9;
b_sign0 = 4'd4; b_sign1 = 4'd7; b_sign2 = 4'd7; b_sign3 = 4'd0;
@(posedge clk_i);
a_mant0 = 8'd145; a_mant1 = 8'd47; a_mant2 = 8'd128; a_mant3 = 8'd252;
b_mant0 = 8'd45; b_mant1 = 8'd37; b_mant2 = 8'd173; b_mant3 = 8'd156;
a_exp0 = 10'd496; a_exp1 = 10'd604; a_exp2 = 10'd796; a_exp3 = 10'd482;
b_exp0 = 10'd982; b_exp1 = 10'd143; b_exp2 = 10'd732; b_exp3 = 10'd374;
a_sign0 = 4'd14; a_sign1 = 4'd3; a_sign2 = 4'd11; a_sign3 = 4'd3;
b_sign0 = 4'd5; b_sign1 = 4'd1; b_sign2 = 4'd3; b_sign3 = 4'd11;
@(posedge clk_i);
a_mant0 = 8'd237; a_mant1 = 8'd100; a_mant2 = 8'd48; a_mant3 = 8'd124;
b_mant0 = 8'd91; b_mant1 = 8'd251; b_mant2 = 8'd185; b_mant3 = 8'd165;
a_exp0 = 10'd650; a_exp1 = 10'd433; a_exp2 = 10'd306; a_exp3 = 10'd620;
b_exp0 = 10'd405; b_exp1 = 10'd459; b_exp2 = 10'd315; b_exp3 = 10'd523;
a_sign0 = 4'd5; a_sign1 = 4'd0; a_sign2 = 4'd11; a_sign3 = 4'd7;
b_sign0 = 4'd5; b_sign1 = 4'd9; b_sign2 = 4'd1; b_sign3 = 4'd9;
@(posedge clk_i);
a_mant0 = 8'd181; a_mant1 = 8'd168; a_mant2 = 8'd148; a_mant3 = 8'd232;
b_mant0 = 8'd103; b_mant1 = 8'd168; b_mant2 = 8'd191; b_mant3 = 8'd171;
a_exp0 = 10'd119; a_exp1 = 10'd109; a_exp2 = 10'd920; a_exp3 = 10'd438;
b_exp0 = 10'd1; b_exp1 = 10'd394; b_exp2 = 10'd600; b_exp3 = 10'd167;
a_sign0 = 4'd4; a_sign1 = 4'd6; a_sign2 = 4'd12; a_sign3 = 4'd14;
b_sign0 = 4'd11; b_sign1 = 4'd13; b_sign2 = 4'd9; b_sign3 = 4'd16;
@(posedge clk_i);
a_mant0 = 8'd179; a_mant1 = 8'd17; a_mant2 = 8'd177; a_mant3 = 8'd222;
b_mant0 = 8'd65; b_mant1 = 8'd73; b_mant2 = 8'd44; b_mant3 = 8'd35;
a_exp0 = 10'd958; a_exp1 = 10'd807; a_exp2 = 10'd672; a_exp3 = 10'd915;
b_exp0 = 10'd743; b_exp1 = 10'd305; b_exp2 = 10'd129; b_exp3 = 10'd751;
a_sign0 = 4'd13; a_sign1 = 4'd11; a_sign2 = 4'd5; a_sign3 = 4'd10;
b_sign0 = 4'd2; b_sign1 = 4'd11; b_sign2 = 4'd5; b_sign3 = 4'd15;
@(posedge clk_i);
shared_exps0 = 8'd154;
shared_exps1 = 8'd120;
a_mant0 = 8'd234; a_mant1 = 8'd80; a_mant2 = 8'd55; a_mant3 = 8'd59;
b_mant0 = 8'd250; b_mant1 = 8'd232; b_mant2 = 8'd180; b_mant3 = 8'd199;
a_exp0 = 10'd228; a_exp1 = 10'd227; a_exp2 = 10'd120; a_exp3 = 10'd634;
b_exp0 = 10'd880; b_exp1 = 10'd42; b_exp2 = 10'd620; b_exp3 = 10'd646;
a_sign0 = 4'd12; a_sign1 = 4'd5; a_sign2 = 4'd9; a_sign3 = 4'd0;
b_sign0 = 4'd0; b_sign1 = 4'd9; b_sign2 = 4'd1; b_sign3 = 4'd14;
@(posedge clk_i);
a_mant0 = 8'd194; a_mant1 = 8'd66; a_mant2 = 8'd98; a_mant3 = 8'd171;
b_mant0 = 8'd28; b_mant1 = 8'd67; b_mant2 = 8'd37; b_mant3 = 8'd48;
a_exp0 = 10'd803; a_exp1 = 10'd396; a_exp2 = 10'd406; a_exp3 = 10'd318;
b_exp0 = 10'd732; b_exp1 = 10'd644; b_exp2 = 10'd190; b_exp3 = 10'd240;
a_sign0 = 4'd3; a_sign1 = 4'd1; a_sign2 = 4'd1; a_sign3 = 4'd2;
b_sign0 = 4'd6; b_sign1 = 4'd7; b_sign2 = 4'd8; b_sign3 = 4'd7;
@(posedge clk_i);
a_mant0 = 8'd56; a_mant1 = 8'd85; a_mant2 = 8'd166; a_mant3 = 8'd213;
b_mant0 = 8'd142; b_mant1 = 8'd49; b_mant2 = 8'd50; b_mant3 = 8'd62;
a_exp0 = 10'd230; a_exp1 = 10'd568; a_exp2 = 10'd843; a_exp3 = 10'd181;
b_exp0 = 10'd231; b_exp1 = 10'd36; b_exp2 = 10'd169; b_exp3 = 10'd974;
a_sign0 = 4'd7; a_sign1 = 4'd5; a_sign2 = 4'd10; a_sign3 = 4'd11;
b_sign0 = 4'd0; b_sign1 = 4'd1; b_sign2 = 4'd6; b_sign3 = 4'd5;
@(posedge clk_i);
a_mant0 = 8'd224; a_mant1 = 8'd98; a_mant2 = 8'd178; a_mant3 = 8'd254;
b_mant0 = 8'd133; b_mant1 = 8'd184; b_mant2 = 8'd221; b_mant3 = 8'd198;
a_exp0 = 10'd140; a_exp1 = 10'd399; a_exp2 = 10'd817; a_exp3 = 10'd378;
b_exp0 = 10'd615; b_exp1 = 10'd439; b_exp2 = 10'd849; b_exp3 = 10'd874;
a_sign0 = 4'd16; a_sign1 = 4'd2; a_sign2 = 4'd15; a_sign3 = 4'd16;
b_sign0 = 4'd1; b_sign1 = 4'd5; b_sign2 = 4'd8; b_sign3 = 4'd12;
@(posedge clk_i);
a_mant0 = 8'd138; a_mant1 = 8'd1; a_mant2 = 8'd233; a_mant3 = 8'd201;
b_mant0 = 8'd172; b_mant1 = 8'd106; b_mant2 = 8'd49; b_mant3 = 8'd173;
a_exp0 = 10'd584; a_exp1 = 10'd414; a_exp2 = 10'd911; a_exp3 = 10'd559;
b_exp0 = 10'd155; b_exp1 = 10'd805; b_exp2 = 10'd180; b_exp3 = 10'd666;
a_sign0 = 4'd8; a_sign1 = 4'd13; a_sign2 = 4'd7; a_sign3 = 4'd7;
b_sign0 = 4'd10; b_sign1 = 4'd16; b_sign2 = 4'd5; b_sign3 = 4'd12;
@(posedge clk_i);
a_mant0 = 8'd97; a_mant1 = 8'd246; a_mant2 = 8'd26; a_mant3 = 8'd248;
b_mant0 = 8'd231; b_mant1 = 8'd64; b_mant2 = 8'd112; b_mant3 = 8'd178;
a_exp0 = 10'd514; a_exp1 = 10'd825; a_exp2 = 10'd31; a_exp3 = 10'd232;
b_exp0 = 10'd5; b_exp1 = 10'd375; b_exp2 = 10'd676; b_exp3 = 10'd136;
a_sign0 = 4'd3; a_sign1 = 4'd6; a_sign2 = 4'd14; a_sign3 = 4'd8;
b_sign0 = 4'd8; b_sign1 = 4'd4; b_sign2 = 4'd8; b_sign3 = 4'd15;
@(posedge clk_i);
a_mant0 = 8'd94; a_mant1 = 8'd156; a_mant2 = 8'd179; a_mant3 = 8'd59;
b_mant0 = 8'd173; b_mant1 = 8'd168; b_mant2 = 8'd116; b_mant3 = 8'd52;
a_exp0 = 10'd105; a_exp1 = 10'd594; a_exp2 = 10'd140; a_exp3 = 10'd420;
b_exp0 = 10'd595; b_exp1 = 10'd540; b_exp2 = 10'd351; b_exp3 = 10'd191;
a_sign0 = 4'd6; a_sign1 = 4'd8; a_sign2 = 4'd9; a_sign3 = 4'd3;
b_sign0 = 4'd5; b_sign1 = 4'd10; b_sign2 = 4'd15; b_sign3 = 4'd16;
@(posedge clk_i);
a_mant0 = 8'd68; a_mant1 = 8'd50; a_mant2 = 8'd193; a_mant3 = 8'd210;
b_mant0 = 8'd158; b_mant1 = 8'd27; b_mant2 = 8'd148; b_mant3 = 8'd186;
a_exp0 = 10'd35; a_exp1 = 10'd411; a_exp2 = 10'd1004; a_exp3 = 10'd710;
b_exp0 = 10'd626; b_exp1 = 10'd417; b_exp2 = 10'd514; b_exp3 = 10'd421;
a_sign0 = 4'd15; a_sign1 = 4'd8; a_sign2 = 4'd1; a_sign3 = 4'd1;
b_sign0 = 4'd16; b_sign1 = 4'd4; b_sign2 = 4'd9; b_sign3 = 4'd8;
@(posedge clk_i);
shared_exps0 = 8'd91;
shared_exps1 = 8'd125;
a_mant0 = 8'd128; a_mant1 = 8'd214; a_mant2 = 8'd196; a_mant3 = 8'd208;
b_mant0 = 8'd160; b_mant1 = 8'd50; b_mant2 = 8'd14; b_mant3 = 8'd111;
a_exp0 = 10'd291; a_exp1 = 10'd7; a_exp2 = 10'd266; a_exp3 = 10'd491;
b_exp0 = 10'd461; b_exp1 = 10'd746; b_exp2 = 10'd509; b_exp3 = 10'd930;
a_sign0 = 4'd10; a_sign1 = 4'd9; a_sign2 = 4'd0; a_sign3 = 4'd14;
b_sign0 = 4'd16; b_sign1 = 4'd10; b_sign2 = 4'd15; b_sign3 = 4'd2;
@(posedge clk_i);
a_mant0 = 8'd155; a_mant1 = 8'd145; a_mant2 = 8'd55; a_mant3 = 8'd120;
b_mant0 = 8'd134; b_mant1 = 8'd179; b_mant2 = 8'd222; b_mant3 = 8'd190;
a_exp0 = 10'd923; a_exp1 = 10'd621; a_exp2 = 10'd590; a_exp3 = 10'd909;
b_exp0 = 10'd485; b_exp1 = 10'd179; b_exp2 = 10'd700; b_exp3 = 10'd87;
a_sign0 = 4'd11; a_sign1 = 4'd1; a_sign2 = 4'd15; a_sign3 = 4'd2;
b_sign0 = 4'd2; b_sign1 = 4'd9; b_sign2 = 4'd16; b_sign3 = 4'd10;
@(posedge clk_i);
a_mant0 = 8'd20; a_mant1 = 8'd62; a_mant2 = 8'd235; a_mant3 = 8'd74;
b_mant0 = 8'd2; b_mant1 = 8'd78; b_mant2 = 8'd209; b_mant3 = 8'd65;
a_exp0 = 10'd21; a_exp1 = 10'd2; a_exp2 = 10'd478; a_exp3 = 10'd361;
b_exp0 = 10'd818; b_exp1 = 10'd103; b_exp2 = 10'd866; b_exp3 = 10'd378;
a_sign0 = 4'd3; a_sign1 = 4'd16; a_sign2 = 4'd5; a_sign3 = 4'd0;
b_sign0 = 4'd12; b_sign1 = 4'd8; b_sign2 = 4'd9; b_sign3 = 4'd5;
@(posedge clk_i);
a_mant0 = 8'd168; a_mant1 = 8'd202; a_mant2 = 8'd207; a_mant3 = 8'd204;
b_mant0 = 8'd108; b_mant1 = 8'd210; b_mant2 = 8'd114; b_mant3 = 8'd35;
a_exp0 = 10'd668; a_exp1 = 10'd615; a_exp2 = 10'd373; a_exp3 = 10'd848;
b_exp0 = 10'd403; b_exp1 = 10'd155; b_exp2 = 10'd37; b_exp3 = 10'd357;
a_sign0 = 4'd16; a_sign1 = 4'd4; a_sign2 = 4'd0; a_sign3 = 4'd6;
b_sign0 = 4'd2; b_sign1 = 4'd12; b_sign2 = 4'd11; b_sign3 = 4'd13;
@(posedge clk_i);
a_mant0 = 8'd57; a_mant1 = 8'd29; a_mant2 = 8'd172; a_mant3 = 8'd247;
b_mant0 = 8'd81; b_mant1 = 8'd1; b_mant2 = 8'd231; b_mant3 = 8'd123;
a_exp0 = 10'd640; a_exp1 = 10'd162; a_exp2 = 10'd940; a_exp3 = 10'd919;
b_exp0 = 10'd102; b_exp1 = 10'd431; b_exp2 = 10'd131; b_exp3 = 10'd55;
a_sign0 = 4'd16; a_sign1 = 4'd16; a_sign2 = 4'd16; a_sign3 = 4'd7;
b_sign0 = 4'd0; b_sign1 = 4'd16; b_sign2 = 4'd15; b_sign3 = 4'd7;
@(posedge clk_i);
a_mant0 = 8'd197; a_mant1 = 8'd34; a_mant2 = 8'd246; a_mant3 = 8'd69;
b_mant0 = 8'd11; b_mant1 = 8'd23; b_mant2 = 8'd92; b_mant3 = 8'd119;
a_exp0 = 10'd981; a_exp1 = 10'd793; a_exp2 = 10'd189; a_exp3 = 10'd679;
b_exp0 = 10'd481; b_exp1 = 10'd295; b_exp2 = 10'd1001; b_exp3 = 10'd245;
a_sign0 = 4'd9; a_sign1 = 4'd14; a_sign2 = 4'd15; a_sign3 = 4'd13;
b_sign0 = 4'd6; b_sign1 = 4'd14; b_sign2 = 4'd12; b_sign3 = 4'd9;
@(posedge clk_i);
a_mant0 = 8'd176; a_mant1 = 8'd236; a_mant2 = 8'd221; a_mant3 = 8'd25;
b_mant0 = 8'd83; b_mant1 = 8'd118; b_mant2 = 8'd97; b_mant3 = 8'd144;
a_exp0 = 10'd926; a_exp1 = 10'd646; a_exp2 = 10'd263; a_exp3 = 10'd471;
b_exp0 = 10'd125; b_exp1 = 10'd244; b_exp2 = 10'd552; b_exp3 = 10'd541;
a_sign0 = 4'd12; a_sign1 = 4'd16; a_sign2 = 4'd16; a_sign3 = 4'd6;
b_sign0 = 4'd9; b_sign1 = 4'd9; b_sign2 = 4'd7; b_sign3 = 4'd1;
@(posedge clk_i);
a_mant0 = 8'd35; a_mant1 = 8'd89; a_mant2 = 8'd65; a_mant3 = 8'd153;
b_mant0 = 8'd42; b_mant1 = 8'd51; b_mant2 = 8'd147; b_mant3 = 8'd188;
a_exp0 = 10'd855; a_exp1 = 10'd291; a_exp2 = 10'd118; a_exp3 = 10'd596;
b_exp0 = 10'd201; b_exp1 = 10'd463; b_exp2 = 10'd699; b_exp3 = 10'd364;
a_sign0 = 4'd10; a_sign1 = 4'd1; a_sign2 = 4'd14; a_sign3 = 4'd10;
b_sign0 = 4'd3; b_sign1 = 4'd2; b_sign2 = 4'd7; b_sign3 = 4'd10;
@(posedge clk_i);
shared_exps0 = 8'd126;
shared_exps1 = 8'd124;
rstn = 0;
@(posedge clk_i);
rstn = 1;
a_mant0 = 8'd252; a_mant1 = 8'd139; a_mant2 = 8'd253; a_mant3 = 8'd199;
b_mant0 = 8'd51; b_mant1 = 8'd116; b_mant2 = 8'd231; b_mant3 = 8'd188;
a_exp0 = 10'd555; a_exp1 = 10'd805; a_exp2 = 10'd884; a_exp3 = 10'd417;
b_exp0 = 10'd25; b_exp1 = 10'd511; b_exp2 = 10'd639; b_exp3 = 10'd243;
a_sign0 = 4'd14; a_sign1 = 4'd12; a_sign2 = 4'd11; a_sign3 = 4'd0;
b_sign0 = 4'd13; b_sign1 = 4'd9; b_sign2 = 4'd2; b_sign3 = 4'd7;
@(posedge clk_i);
a_mant0 = 8'd26; a_mant1 = 8'd220; a_mant2 = 8'd57; a_mant3 = 8'd12;
b_mant0 = 8'd213; b_mant1 = 8'd134; b_mant2 = 8'd73; b_mant3 = 8'd118;
a_exp0 = 10'd1005; a_exp1 = 10'd185; a_exp2 = 10'd757; a_exp3 = 10'd953;
b_exp0 = 10'd677; b_exp1 = 10'd234; b_exp2 = 10'd682; b_exp3 = 10'd406;
a_sign0 = 4'd11; a_sign1 = 4'd4; a_sign2 = 4'd4; a_sign3 = 4'd10;
b_sign0 = 4'd13; b_sign1 = 4'd6; b_sign2 = 4'd2; b_sign3 = 4'd3;
@(posedge clk_i);
a_mant0 = 8'd126; a_mant1 = 8'd151; a_mant2 = 8'd60; a_mant3 = 8'd110;
b_mant0 = 8'd106; b_mant1 = 8'd113; b_mant2 = 8'd161; b_mant3 = 8'd26;
a_exp0 = 10'd801; a_exp1 = 10'd443; a_exp2 = 10'd789; a_exp3 = 10'd106;
b_exp0 = 10'd517; b_exp1 = 10'd312; b_exp2 = 10'd987; b_exp3 = 10'd1000;
a_sign0 = 4'd8; a_sign1 = 4'd1; a_sign2 = 4'd10; a_sign3 = 4'd12;
b_sign0 = 4'd13; b_sign1 = 4'd10; b_sign2 = 4'd0; b_sign3 = 4'd4;
@(posedge clk_i);
a_mant0 = 8'd140; a_mant1 = 8'd122; a_mant2 = 8'd47; a_mant3 = 8'd248;
b_mant0 = 8'd217; b_mant1 = 8'd192; b_mant2 = 8'd71; b_mant3 = 8'd121;
a_exp0 = 10'd470; a_exp1 = 10'd967; a_exp2 = 10'd823; a_exp3 = 10'd72;
b_exp0 = 10'd697; b_exp1 = 10'd981; b_exp2 = 10'd587; b_exp3 = 10'd697;
a_sign0 = 4'd14; a_sign1 = 4'd12; a_sign2 = 4'd13; a_sign3 = 4'd9;
b_sign0 = 4'd15; b_sign1 = 4'd1; b_sign2 = 4'd9; b_sign3 = 4'd16;
@(posedge clk_i);
a_mant0 = 8'd153; a_mant1 = 8'd222; a_mant2 = 8'd203; a_mant3 = 8'd77;
b_mant0 = 8'd207; b_mant1 = 8'd113; b_mant2 = 8'd188; b_mant3 = 8'd199;
a_exp0 = 10'd203; a_exp1 = 10'd407; a_exp2 = 10'd817; a_exp3 = 10'd188;
b_exp0 = 10'd574; b_exp1 = 10'd276; b_exp2 = 10'd981; b_exp3 = 10'd32;
a_sign0 = 4'd15; a_sign1 = 4'd13; a_sign2 = 4'd8; a_sign3 = 4'd5;
b_sign0 = 4'd10; b_sign1 = 4'd8; b_sign2 = 4'd16; b_sign3 = 4'd7;
@(posedge clk_i);
a_mant0 = 8'd250; a_mant1 = 8'd139; a_mant2 = 8'd110; a_mant3 = 8'd133;
b_mant0 = 8'd180; b_mant1 = 8'd162; b_mant2 = 8'd245; b_mant3 = 8'd35;
a_exp0 = 10'd977; a_exp1 = 10'd474; a_exp2 = 10'd485; a_exp3 = 10'd754;
b_exp0 = 10'd420; b_exp1 = 10'd902; b_exp2 = 10'd651; b_exp3 = 10'd43;
a_sign0 = 4'd16; a_sign1 = 4'd0; a_sign2 = 4'd0; a_sign3 = 4'd15;
b_sign0 = 4'd2; b_sign1 = 4'd3; b_sign2 = 4'd15; b_sign3 = 4'd16;
@(posedge clk_i);
a_mant0 = 8'd149; a_mant1 = 8'd240; a_mant2 = 8'd168; a_mant3 = 8'd0;
b_mant0 = 8'd182; b_mant1 = 8'd166; b_mant2 = 8'd187; b_mant3 = 8'd248;
a_exp0 = 10'd331; a_exp1 = 10'd277; a_exp2 = 10'd388; a_exp3 = 10'd733;
b_exp0 = 10'd779; b_exp1 = 10'd407; b_exp2 = 10'd863; b_exp3 = 10'd959;
a_sign0 = 4'd7; a_sign1 = 4'd2; a_sign2 = 4'd6; a_sign3 = 4'd5;
b_sign0 = 4'd16; b_sign1 = 4'd8; b_sign2 = 4'd15; b_sign3 = 4'd3;
@(posedge clk_i);
shared_exps0 = 8'd138;
shared_exps1 = 8'd150;
a_mant0 = 8'd71; a_mant1 = 8'd164; a_mant2 = 8'd231; a_mant3 = 8'd96;
b_mant0 = 8'd59; b_mant1 = 8'd37; b_mant2 = 8'd232; b_mant3 = 8'd7;
a_exp0 = 10'd172; a_exp1 = 10'd80; a_exp2 = 10'd745; a_exp3 = 10'd466;
b_exp0 = 10'd837; b_exp1 = 10'd316; b_exp2 = 10'd319; b_exp3 = 10'd807;
a_sign0 = 4'd0; a_sign1 = 4'd12; a_sign2 = 4'd2; a_sign3 = 4'd16;
b_sign0 = 4'd4; b_sign1 = 4'd8; b_sign2 = 4'd7; b_sign3 = 4'd10;
@(posedge clk_i);
a_mant0 = 8'd215; a_mant1 = 8'd22; a_mant2 = 8'd12; a_mant3 = 8'd206;
b_mant0 = 8'd214; b_mant1 = 8'd60; b_mant2 = 8'd107; b_mant3 = 8'd109;
a_exp0 = 10'd51; a_exp1 = 10'd815; a_exp2 = 10'd38; a_exp3 = 10'd788;
b_exp0 = 10'd829; b_exp1 = 10'd212; b_exp2 = 10'd182; b_exp3 = 10'd666;
a_sign0 = 4'd13; a_sign1 = 4'd16; a_sign2 = 4'd8; a_sign3 = 4'd13;
b_sign0 = 4'd7; b_sign1 = 4'd0; b_sign2 = 4'd13; b_sign3 = 4'd4;
@(posedge clk_i);
a_mant0 = 8'd182; a_mant1 = 8'd45; a_mant2 = 8'd179; a_mant3 = 8'd124;
b_mant0 = 8'd195; b_mant1 = 8'd98; b_mant2 = 8'd86; b_mant3 = 8'd123;
a_exp0 = 10'd816; a_exp1 = 10'd144; a_exp2 = 10'd237; a_exp3 = 10'd169;
b_exp0 = 10'd888; b_exp1 = 10'd868; b_exp2 = 10'd777; b_exp3 = 10'd655;
a_sign0 = 4'd9; a_sign1 = 4'd7; a_sign2 = 4'd12; a_sign3 = 4'd5;
b_sign0 = 4'd5; b_sign1 = 4'd16; b_sign2 = 4'd1; b_sign3 = 4'd14;
@(posedge clk_i);
a_mant0 = 8'd31; a_mant1 = 8'd69; a_mant2 = 8'd190; a_mant3 = 8'd158;
b_mant0 = 8'd165; b_mant1 = 8'd78; b_mant2 = 8'd239; b_mant3 = 8'd197;
a_exp0 = 10'd882; a_exp1 = 10'd402; a_exp2 = 10'd293; a_exp3 = 10'd420;
b_exp0 = 10'd541; b_exp1 = 10'd297; b_exp2 = 10'd494; b_exp3 = 10'd937;
a_sign0 = 4'd16; a_sign1 = 4'd0; a_sign2 = 4'd0; a_sign3 = 4'd9;
b_sign0 = 4'd7; b_sign1 = 4'd0; b_sign2 = 4'd14; b_sign3 = 4'd15;
@(posedge clk_i);
a_mant0 = 8'd44; a_mant1 = 8'd44; a_mant2 = 8'd74; a_mant3 = 8'd142;
b_mant0 = 8'd145; b_mant1 = 8'd163; b_mant2 = 8'd5; b_mant3 = 8'd250;
a_exp0 = 10'd653; a_exp1 = 10'd804; a_exp2 = 10'd391; a_exp3 = 10'd586;
b_exp0 = 10'd195; b_exp1 = 10'd997; b_exp2 = 10'd1; b_exp3 = 10'd886;
a_sign0 = 4'd5; a_sign1 = 4'd9; a_sign2 = 4'd9; a_sign3 = 4'd8;
b_sign0 = 4'd4; b_sign1 = 4'd14; b_sign2 = 4'd10; b_sign3 = 4'd9;
@(posedge clk_i);
a_mant0 = 8'd170; a_mant1 = 8'd165; a_mant2 = 8'd233; a_mant3 = 8'd249;
b_mant0 = 8'd146; b_mant1 = 8'd26; b_mant2 = 8'd240; b_mant3 = 8'd159;
a_exp0 = 10'd497; a_exp1 = 10'd738; a_exp2 = 10'd41; a_exp3 = 10'd726;
b_exp0 = 10'd963; b_exp1 = 10'd762; b_exp2 = 10'd880; b_exp3 = 10'd379;
a_sign0 = 4'd3; a_sign1 = 4'd6; a_sign2 = 4'd14; a_sign3 = 4'd10;
b_sign0 = 4'd15; b_sign1 = 4'd15; b_sign2 = 4'd3; b_sign3 = 4'd1;
@(posedge clk_i);
a_mant0 = 8'd153; a_mant1 = 8'd249; a_mant2 = 8'd102; a_mant3 = 8'd94;
b_mant0 = 8'd227; b_mant1 = 8'd1; b_mant2 = 8'd41; b_mant3 = 8'd197;
a_exp0 = 10'd455; a_exp1 = 10'd537; a_exp2 = 10'd221; a_exp3 = 10'd116;
b_exp0 = 10'd846; b_exp1 = 10'd879; b_exp2 = 10'd289; b_exp3 = 10'd653;
a_sign0 = 4'd1; a_sign1 = 4'd0; a_sign2 = 4'd15; a_sign3 = 4'd3;
b_sign0 = 4'd1; b_sign1 = 4'd11; b_sign2 = 4'd15; b_sign3 = 4'd10;
@(posedge clk_i);
a_mant0 = 8'd36; a_mant1 = 8'd167; a_mant2 = 8'd16; a_mant3 = 8'd36;
b_mant0 = 8'd12; b_mant1 = 8'd137; b_mant2 = 8'd122; b_mant3 = 8'd210;
a_exp0 = 10'd501; a_exp1 = 10'd245; a_exp2 = 10'd808; a_exp3 = 10'd488;
b_exp0 = 10'd640; b_exp1 = 10'd660; b_exp2 = 10'd1; b_exp3 = 10'd252;
a_sign0 = 4'd10; a_sign1 = 4'd10; a_sign2 = 4'd14; a_sign3 = 4'd6;
b_sign0 = 4'd13; b_sign1 = 4'd13; b_sign2 = 4'd2; b_sign3 = 4'd10;
@(posedge clk_i);
shared_exps0 = 8'd116;
shared_exps1 = 8'd133;
a_mant0 = 8'd162; a_mant1 = 8'd171; a_mant2 = 8'd33; a_mant3 = 8'd179;
b_mant0 = 8'd140; b_mant1 = 8'd83; b_mant2 = 8'd126; b_mant3 = 8'd193;
a_exp0 = 10'd852; a_exp1 = 10'd409; a_exp2 = 10'd930; a_exp3 = 10'd838;
b_exp0 = 10'd200; b_exp1 = 10'd211; b_exp2 = 10'd252; b_exp3 = 10'd18;
a_sign0 = 4'd0; a_sign1 = 4'd12; a_sign2 = 4'd4; a_sign3 = 4'd13;
b_sign0 = 4'd10; b_sign1 = 4'd0; b_sign2 = 4'd5; b_sign3 = 4'd11;
@(posedge clk_i);
a_mant0 = 8'd65; a_mant1 = 8'd244; a_mant2 = 8'd249; a_mant3 = 8'd93;
b_mant0 = 8'd97; b_mant1 = 8'd89; b_mant2 = 8'd13; b_mant3 = 8'd83;
a_exp0 = 10'd347; a_exp1 = 10'd1023; a_exp2 = 10'd925; a_exp3 = 10'd974;
b_exp0 = 10'd864; b_exp1 = 10'd485; b_exp2 = 10'd892; b_exp3 = 10'd587;
a_sign0 = 4'd0; a_sign1 = 4'd9; a_sign2 = 4'd16; a_sign3 = 4'd0;
b_sign0 = 4'd5; b_sign1 = 4'd1; b_sign2 = 4'd13; b_sign3 = 4'd6;
@(posedge clk_i);
a_mant0 = 8'd32; a_mant1 = 8'd141; a_mant2 = 8'd138; a_mant3 = 8'd50;
b_mant0 = 8'd28; b_mant1 = 8'd11; b_mant2 = 8'd70; b_mant3 = 8'd105;
a_exp0 = 10'd704; a_exp1 = 10'd6; a_exp2 = 10'd325; a_exp3 = 10'd903;
b_exp0 = 10'd305; b_exp1 = 10'd505; b_exp2 = 10'd220; b_exp3 = 10'd153;
a_sign0 = 4'd0; a_sign1 = 4'd4; a_sign2 = 4'd3; a_sign3 = 4'd9;
b_sign0 = 4'd1; b_sign1 = 4'd14; b_sign2 = 4'd10; b_sign3 = 4'd6;
@(posedge clk_i);
a_mant0 = 8'd241; a_mant1 = 8'd225; a_mant2 = 8'd201; a_mant3 = 8'd160;
b_mant0 = 8'd136; b_mant1 = 8'd126; b_mant2 = 8'd135; b_mant3 = 8'd82;
a_exp0 = 10'd959; a_exp1 = 10'd734; a_exp2 = 10'd48; a_exp3 = 10'd650;
b_exp0 = 10'd996; b_exp1 = 10'd269; b_exp2 = 10'd350; b_exp3 = 10'd991;
a_sign0 = 4'd7; a_sign1 = 4'd9; a_sign2 = 4'd15; a_sign3 = 4'd6;
b_sign0 = 4'd1; b_sign1 = 4'd5; b_sign2 = 4'd16; b_sign3 = 4'd11;
@(posedge clk_i);
a_mant0 = 8'd61; a_mant1 = 8'd221; a_mant2 = 8'd234; a_mant3 = 8'd124;
b_mant0 = 8'd81; b_mant1 = 8'd97; b_mant2 = 8'd36; b_mant3 = 8'd231;
a_exp0 = 10'd337; a_exp1 = 10'd103; a_exp2 = 10'd58; a_exp3 = 10'd341;
b_exp0 = 10'd759; b_exp1 = 10'd13; b_exp2 = 10'd166; b_exp3 = 10'd570;
a_sign0 = 4'd1; a_sign1 = 4'd4; a_sign2 = 4'd16; a_sign3 = 4'd6;
b_sign0 = 4'd2; b_sign1 = 4'd4; b_sign2 = 4'd7; b_sign3 = 4'd2;
@(posedge clk_i);
a_mant0 = 8'd223; a_mant1 = 8'd176; a_mant2 = 8'd54; a_mant3 = 8'd141;
b_mant0 = 8'd61; b_mant1 = 8'd129; b_mant2 = 8'd234; b_mant3 = 8'd44;
a_exp0 = 10'd113; a_exp1 = 10'd953; a_exp2 = 10'd696; a_exp3 = 10'd187;
b_exp0 = 10'd155; b_exp1 = 10'd157; b_exp2 = 10'd141; b_exp3 = 10'd58;
a_sign0 = 4'd11; a_sign1 = 4'd14; a_sign2 = 4'd5; a_sign3 = 4'd9;
b_sign0 = 4'd13; b_sign1 = 4'd13; b_sign2 = 4'd9; b_sign3 = 4'd12;
@(posedge clk_i);
a_mant0 = 8'd119; a_mant1 = 8'd42; a_mant2 = 8'd60; a_mant3 = 8'd213;
b_mant0 = 8'd28; b_mant1 = 8'd41; b_mant2 = 8'd6; b_mant3 = 8'd124;
a_exp0 = 10'd458; a_exp1 = 10'd911; a_exp2 = 10'd798; a_exp3 = 10'd184;
b_exp0 = 10'd735; b_exp1 = 10'd82; b_exp2 = 10'd768; b_exp3 = 10'd782;
a_sign0 = 4'd0; a_sign1 = 4'd12; a_sign2 = 4'd7; a_sign3 = 4'd7;
b_sign0 = 4'd3; b_sign1 = 4'd12; b_sign2 = 4'd1; b_sign3 = 4'd11;
@(posedge clk_i);
a_mant0 = 8'd150; a_mant1 = 8'd127; a_mant2 = 8'd38; a_mant3 = 8'd164;
b_mant0 = 8'd199; b_mant1 = 8'd231; b_mant2 = 8'd255; b_mant3 = 8'd124;
a_exp0 = 10'd188; a_exp1 = 10'd168; a_exp2 = 10'd946; a_exp3 = 10'd636;
b_exp0 = 10'd919; b_exp1 = 10'd975; b_exp2 = 10'd645; b_exp3 = 10'd206;
a_sign0 = 4'd5; a_sign1 = 4'd14; a_sign2 = 4'd7; a_sign3 = 4'd10;
b_sign0 = 4'd7; b_sign1 = 4'd16; b_sign2 = 4'd15; b_sign3 = 4'd16;
@(posedge clk_i);
shared_exps0 = 8'd110;
shared_exps1 = 8'd124;
a_mant0 = 8'd54; a_mant1 = 8'd202; a_mant2 = 8'd149; a_mant3 = 8'd27;
b_mant0 = 8'd48; b_mant1 = 8'd0; b_mant2 = 8'd196; b_mant3 = 8'd13;
a_exp0 = 10'd124; a_exp1 = 10'd84; a_exp2 = 10'd267; a_exp3 = 10'd722;
b_exp0 = 10'd311; b_exp1 = 10'd193; b_exp2 = 10'd931; b_exp3 = 10'd314;
a_sign0 = 4'd16; a_sign1 = 4'd10; a_sign2 = 4'd16; a_sign3 = 4'd15;
b_sign0 = 4'd7; b_sign1 = 4'd1; b_sign2 = 4'd9; b_sign3 = 4'd0;
@(posedge clk_i);
a_mant0 = 8'd116; a_mant1 = 8'd242; a_mant2 = 8'd207; a_mant3 = 8'd155;
b_mant0 = 8'd131; b_mant1 = 8'd219; b_mant2 = 8'd204; b_mant3 = 8'd109;
a_exp0 = 10'd817; a_exp1 = 10'd231; a_exp2 = 10'd195; a_exp3 = 10'd115;
b_exp0 = 10'd755; b_exp1 = 10'd9; b_exp2 = 10'd322; b_exp3 = 10'd550;
a_sign0 = 4'd0; a_sign1 = 4'd2; a_sign2 = 4'd15; a_sign3 = 4'd5;
b_sign0 = 4'd6; b_sign1 = 4'd0; b_sign2 = 4'd14; b_sign3 = 4'd1;
@(posedge clk_i);
a_mant0 = 8'd88; a_mant1 = 8'd185; a_mant2 = 8'd148; a_mant3 = 8'd48;
b_mant0 = 8'd123; b_mant1 = 8'd150; b_mant2 = 8'd125; b_mant3 = 8'd167;
a_exp0 = 10'd814; a_exp1 = 10'd895; a_exp2 = 10'd629; a_exp3 = 10'd151;
b_exp0 = 10'd14; b_exp1 = 10'd653; b_exp2 = 10'd217; b_exp3 = 10'd3;
a_sign0 = 4'd13; a_sign1 = 4'd4; a_sign2 = 4'd15; a_sign3 = 4'd7;
b_sign0 = 4'd15; b_sign1 = 4'd0; b_sign2 = 4'd1; b_sign3 = 4'd0;
@(posedge clk_i);
a_mant0 = 8'd158; a_mant1 = 8'd2; a_mant2 = 8'd241; a_mant3 = 8'd49;
b_mant0 = 8'd132; b_mant1 = 8'd180; b_mant2 = 8'd85; b_mant3 = 8'd115;
a_exp0 = 10'd486; a_exp1 = 10'd514; a_exp2 = 10'd243; a_exp3 = 10'd111;
b_exp0 = 10'd841; b_exp1 = 10'd770; b_exp2 = 10'd939; b_exp3 = 10'd356;
a_sign0 = 4'd9; a_sign1 = 4'd13; a_sign2 = 4'd12; a_sign3 = 4'd16;
b_sign0 = 4'd4; b_sign1 = 4'd9; b_sign2 = 4'd13; b_sign3 = 4'd4;
@(posedge clk_i);
a_mant0 = 8'd174; a_mant1 = 8'd41; a_mant2 = 8'd181; a_mant3 = 8'd162;
b_mant0 = 8'd87; b_mant1 = 8'd174; b_mant2 = 8'd12; b_mant3 = 8'd110;
a_exp0 = 10'd497; a_exp1 = 10'd287; a_exp2 = 10'd295; a_exp3 = 10'd190;
b_exp0 = 10'd401; b_exp1 = 10'd541; b_exp2 = 10'd484; b_exp3 = 10'd351;
a_sign0 = 4'd15; a_sign1 = 4'd9; a_sign2 = 4'd3; a_sign3 = 4'd8;
b_sign0 = 4'd4; b_sign1 = 4'd8; b_sign2 = 4'd15; b_sign3 = 4'd13;
@(posedge clk_i);
a_mant0 = 8'd131; a_mant1 = 8'd145; a_mant2 = 8'd134; a_mant3 = 8'd248;
b_mant0 = 8'd82; b_mant1 = 8'd155; b_mant2 = 8'd180; b_mant3 = 8'd229;
a_exp0 = 10'd367; a_exp1 = 10'd959; a_exp2 = 10'd10; a_exp3 = 10'd957;
b_exp0 = 10'd887; b_exp1 = 10'd926; b_exp2 = 10'd387; b_exp3 = 10'd908;
a_sign0 = 4'd7; a_sign1 = 4'd8; a_sign2 = 4'd7; a_sign3 = 4'd0;
b_sign0 = 4'd7; b_sign1 = 4'd1; b_sign2 = 4'd2; b_sign3 = 4'd5;
@(posedge clk_i);
a_mant0 = 8'd160; a_mant1 = 8'd95; a_mant2 = 8'd59; a_mant3 = 8'd201;
b_mant0 = 8'd100; b_mant1 = 8'd104; b_mant2 = 8'd69; b_mant3 = 8'd2;
a_exp0 = 10'd490; a_exp1 = 10'd770; a_exp2 = 10'd856; a_exp3 = 10'd530;
b_exp0 = 10'd107; b_exp1 = 10'd71; b_exp2 = 10'd270; b_exp3 = 10'd766;
a_sign0 = 4'd4; a_sign1 = 4'd1; a_sign2 = 4'd5; a_sign3 = 4'd1;
b_sign0 = 4'd0; b_sign1 = 4'd14; b_sign2 = 4'd10; b_sign3 = 4'd8;
@(posedge clk_i);
a_mant0 = 8'd85; a_mant1 = 8'd90; a_mant2 = 8'd139; a_mant3 = 8'd239;
b_mant0 = 8'd136; b_mant1 = 8'd133; b_mant2 = 8'd109; b_mant3 = 8'd183;
a_exp0 = 10'd340; a_exp1 = 10'd39; a_exp2 = 10'd635; a_exp3 = 10'd166;
b_exp0 = 10'd97; b_exp1 = 10'd516; b_exp2 = 10'd806; b_exp3 = 10'd534;
a_sign0 = 4'd13; a_sign1 = 4'd6; a_sign2 = 4'd5; a_sign3 = 4'd12;
b_sign0 = 4'd7; b_sign1 = 4'd9; b_sign2 = 4'd16; b_sign3 = 4'd6;
@(posedge clk_i);
shared_exps0 = 8'd124;
shared_exps1 = 8'd82;
rstn = 0;
@(posedge clk_i);
rstn = 1;
a_mant0 = 8'd47; a_mant1 = 8'd129; a_mant2 = 8'd168; a_mant3 = 8'd70;
b_mant0 = 8'd162; b_mant1 = 8'd64; b_mant2 = 8'd26; b_mant3 = 8'd55;
a_exp0 = 10'd649; a_exp1 = 10'd814; a_exp2 = 10'd755; a_exp3 = 10'd869;
b_exp0 = 10'd434; b_exp1 = 10'd617; b_exp2 = 10'd721; b_exp3 = 10'd168;
a_sign0 = 4'd12; a_sign1 = 4'd10; a_sign2 = 4'd3; a_sign3 = 4'd6;
b_sign0 = 4'd7; b_sign1 = 4'd15; b_sign2 = 4'd13; b_sign3 = 4'd8;
@(posedge clk_i);
a_mant0 = 8'd32; a_mant1 = 8'd220; a_mant2 = 8'd53; a_mant3 = 8'd193;
b_mant0 = 8'd165; b_mant1 = 8'd59; b_mant2 = 8'd206; b_mant3 = 8'd112;
a_exp0 = 10'd623; a_exp1 = 10'd318; a_exp2 = 10'd200; a_exp3 = 10'd880;
b_exp0 = 10'd687; b_exp1 = 10'd678; b_exp2 = 10'd381; b_exp3 = 10'd661;
a_sign0 = 4'd3; a_sign1 = 4'd13; a_sign2 = 4'd14; a_sign3 = 4'd4;
b_sign0 = 4'd9; b_sign1 = 4'd5; b_sign2 = 4'd0; b_sign3 = 4'd5;
@(posedge clk_i);
a_mant0 = 8'd201; a_mant1 = 8'd64; a_mant2 = 8'd142; a_mant3 = 8'd201;
b_mant0 = 8'd181; b_mant1 = 8'd117; b_mant2 = 8'd187; b_mant3 = 8'd223;
a_exp0 = 10'd130; a_exp1 = 10'd907; a_exp2 = 10'd510; a_exp3 = 10'd854;
b_exp0 = 10'd361; b_exp1 = 10'd509; b_exp2 = 10'd630; b_exp3 = 10'd722;
a_sign0 = 4'd5; a_sign1 = 4'd16; a_sign2 = 4'd9; a_sign3 = 4'd14;
b_sign0 = 4'd12; b_sign1 = 4'd15; b_sign2 = 4'd3; b_sign3 = 4'd5;
@(posedge clk_i);
a_mant0 = 8'd87; a_mant1 = 8'd111; a_mant2 = 8'd161; a_mant3 = 8'd40;
b_mant0 = 8'd92; b_mant1 = 8'd130; b_mant2 = 8'd44; b_mant3 = 8'd195;
a_exp0 = 10'd493; a_exp1 = 10'd519; a_exp2 = 10'd522; a_exp3 = 10'd181;
b_exp0 = 10'd620; b_exp1 = 10'd569; b_exp2 = 10'd536; b_exp3 = 10'd1005;
a_sign0 = 4'd5; a_sign1 = 4'd7; a_sign2 = 4'd4; a_sign3 = 4'd4;
b_sign0 = 4'd1; b_sign1 = 4'd2; b_sign2 = 4'd9; b_sign3 = 4'd14;
@(posedge clk_i);
a_mant0 = 8'd80; a_mant1 = 8'd226; a_mant2 = 8'd166; a_mant3 = 8'd226;
b_mant0 = 8'd144; b_mant1 = 8'd95; b_mant2 = 8'd208; b_mant3 = 8'd226;
a_exp0 = 10'd212; a_exp1 = 10'd95; a_exp2 = 10'd790; a_exp3 = 10'd921;
b_exp0 = 10'd152; b_exp1 = 10'd459; b_exp2 = 10'd38; b_exp3 = 10'd999;
a_sign0 = 4'd13; a_sign1 = 4'd10; a_sign2 = 4'd16; a_sign3 = 4'd7;
b_sign0 = 4'd4; b_sign1 = 4'd14; b_sign2 = 4'd11; b_sign3 = 4'd4;
@(posedge clk_i);
a_mant0 = 8'd33; a_mant1 = 8'd181; a_mant2 = 8'd6; a_mant3 = 8'd246;
b_mant0 = 8'd218; b_mant1 = 8'd232; b_mant2 = 8'd105; b_mant3 = 8'd179;
a_exp0 = 10'd978; a_exp1 = 10'd121; a_exp2 = 10'd494; a_exp3 = 10'd863;
b_exp0 = 10'd768; b_exp1 = 10'd838; b_exp2 = 10'd666; b_exp3 = 10'd305;
a_sign0 = 4'd8; a_sign1 = 4'd14; a_sign2 = 4'd12; a_sign3 = 4'd8;
b_sign0 = 4'd10; b_sign1 = 4'd12; b_sign2 = 4'd3; b_sign3 = 4'd11;
@(posedge clk_i);
a_mant0 = 8'd79; a_mant1 = 8'd190; a_mant2 = 8'd65; a_mant3 = 8'd58;
b_mant0 = 8'd147; b_mant1 = 8'd181; b_mant2 = 8'd180; b_mant3 = 8'd12;
a_exp0 = 10'd723; a_exp1 = 10'd764; a_exp2 = 10'd941; a_exp3 = 10'd943;
b_exp0 = 10'd1019; b_exp1 = 10'd862; b_exp2 = 10'd254; b_exp3 = 10'd243;
a_sign0 = 4'd15; a_sign1 = 4'd6; a_sign2 = 4'd14; a_sign3 = 4'd14;
b_sign0 = 4'd6; b_sign1 = 4'd16; b_sign2 = 4'd16; b_sign3 = 4'd16;
@(posedge clk_i);
shared_exps0 = 8'd136;
shared_exps1 = 8'd126;
a_mant0 = 8'd40; a_mant1 = 8'd149; a_mant2 = 8'd16; a_mant3 = 8'd117;
b_mant0 = 8'd159; b_mant1 = 8'd76; b_mant2 = 8'd50; b_mant3 = 8'd231;
a_exp0 = 10'd812; a_exp1 = 10'd74; a_exp2 = 10'd391; a_exp3 = 10'd536;
b_exp0 = 10'd600; b_exp1 = 10'd64; b_exp2 = 10'd790; b_exp3 = 10'd659;
a_sign0 = 4'd2; a_sign1 = 4'd4; a_sign2 = 4'd2; a_sign3 = 4'd14;
b_sign0 = 4'd13; b_sign1 = 4'd14; b_sign2 = 4'd13; b_sign3 = 4'd6;
@(posedge clk_i);
a_mant0 = 8'd78; a_mant1 = 8'd222; a_mant2 = 8'd221; a_mant3 = 8'd204;
b_mant0 = 8'd30; b_mant1 = 8'd91; b_mant2 = 8'd151; b_mant3 = 8'd0;
a_exp0 = 10'd802; a_exp1 = 10'd978; a_exp2 = 10'd469; a_exp3 = 10'd267;
b_exp0 = 10'd97; b_exp1 = 10'd62; b_exp2 = 10'd480; b_exp3 = 10'd915;
a_sign0 = 4'd10; a_sign1 = 4'd7; a_sign2 = 4'd16; a_sign3 = 4'd5;
b_sign0 = 4'd13; b_sign1 = 4'd5; b_sign2 = 4'd3; b_sign3 = 4'd2;
@(posedge clk_i);
a_mant0 = 8'd220; a_mant1 = 8'd1; a_mant2 = 8'd246; a_mant3 = 8'd177;
b_mant0 = 8'd173; b_mant1 = 8'd38; b_mant2 = 8'd246; b_mant3 = 8'd118;
a_exp0 = 10'd190; a_exp1 = 10'd954; a_exp2 = 10'd1000; a_exp3 = 10'd1004;
b_exp0 = 10'd237; b_exp1 = 10'd344; b_exp2 = 10'd70; b_exp3 = 10'd751;
a_sign0 = 4'd14; a_sign1 = 4'd12; a_sign2 = 4'd5; a_sign3 = 4'd0;
b_sign0 = 4'd13; b_sign1 = 4'd0; b_sign2 = 4'd3; b_sign3 = 4'd16;
@(posedge clk_i);
a_mant0 = 8'd112; a_mant1 = 8'd30; a_mant2 = 8'd210; a_mant3 = 8'd24;
b_mant0 = 8'd208; b_mant1 = 8'd16; b_mant2 = 8'd36; b_mant3 = 8'd163;
a_exp0 = 10'd269; a_exp1 = 10'd461; a_exp2 = 10'd735; a_exp3 = 10'd81;
b_exp0 = 10'd932; b_exp1 = 10'd778; b_exp2 = 10'd847; b_exp3 = 10'd572;
a_sign0 = 4'd13; a_sign1 = 4'd11; a_sign2 = 4'd10; a_sign3 = 4'd9;
b_sign0 = 4'd7; b_sign1 = 4'd13; b_sign2 = 4'd11; b_sign3 = 4'd8;
@(posedge clk_i);
a_mant0 = 8'd180; a_mant1 = 8'd178; a_mant2 = 8'd41; a_mant3 = 8'd177;
b_mant0 = 8'd109; b_mant1 = 8'd219; b_mant2 = 8'd31; b_mant3 = 8'd82;
a_exp0 = 10'd750; a_exp1 = 10'd708; a_exp2 = 10'd764; a_exp3 = 10'd76;
b_exp0 = 10'd147; b_exp1 = 10'd824; b_exp2 = 10'd868; b_exp3 = 10'd724;
a_sign0 = 4'd6; a_sign1 = 4'd1; a_sign2 = 4'd9; a_sign3 = 4'd7;
b_sign0 = 4'd13; b_sign1 = 4'd15; b_sign2 = 4'd5; b_sign3 = 4'd10;
@(posedge clk_i);
a_mant0 = 8'd163; a_mant1 = 8'd253; a_mant2 = 8'd200; a_mant3 = 8'd247;
b_mant0 = 8'd200; b_mant1 = 8'd51; b_mant2 = 8'd176; b_mant3 = 8'd120;
a_exp0 = 10'd516; a_exp1 = 10'd101; a_exp2 = 10'd221; a_exp3 = 10'd691;
b_exp0 = 10'd564; b_exp1 = 10'd587; b_exp2 = 10'd107; b_exp3 = 10'd667;
a_sign0 = 4'd15; a_sign1 = 4'd4; a_sign2 = 4'd8; a_sign3 = 4'd1;
b_sign0 = 4'd8; b_sign1 = 4'd5; b_sign2 = 4'd2; b_sign3 = 4'd1;
@(posedge clk_i);
a_mant0 = 8'd249; a_mant1 = 8'd70; a_mant2 = 8'd162; a_mant3 = 8'd227;
b_mant0 = 8'd135; b_mant1 = 8'd60; b_mant2 = 8'd193; b_mant3 = 8'd67;
a_exp0 = 10'd1002; a_exp1 = 10'd831; a_exp2 = 10'd711; a_exp3 = 10'd914;
b_exp0 = 10'd237; b_exp1 = 10'd662; b_exp2 = 10'd753; b_exp3 = 10'd642;
a_sign0 = 4'd11; a_sign1 = 4'd7; a_sign2 = 4'd11; a_sign3 = 4'd5;
b_sign0 = 4'd5; b_sign1 = 4'd1; b_sign2 = 4'd5; b_sign3 = 4'd0;
@(posedge clk_i);
a_mant0 = 8'd234; a_mant1 = 8'd141; a_mant2 = 8'd72; a_mant3 = 8'd186;
b_mant0 = 8'd18; b_mant1 = 8'd195; b_mant2 = 8'd224; b_mant3 = 8'd182;
a_exp0 = 10'd398; a_exp1 = 10'd1000; a_exp2 = 10'd41; a_exp3 = 10'd476;
b_exp0 = 10'd20; b_exp1 = 10'd40; b_exp2 = 10'd370; b_exp3 = 10'd626;
a_sign0 = 4'd9; a_sign1 = 4'd11; a_sign2 = 4'd10; a_sign3 = 4'd9;
b_sign0 = 4'd0; b_sign1 = 4'd1; b_sign2 = 4'd13; b_sign3 = 4'd12;
@(posedge clk_i);
shared_exps0 = 8'd138;
shared_exps1 = 8'd95;
a_mant0 = 8'd15; a_mant1 = 8'd136; a_mant2 = 8'd79; a_mant3 = 8'd48;
b_mant0 = 8'd250; b_mant1 = 8'd90; b_mant2 = 8'd252; b_mant3 = 8'd117;
a_exp0 = 10'd68; a_exp1 = 10'd658; a_exp2 = 10'd302; a_exp3 = 10'd994;
b_exp0 = 10'd422; b_exp1 = 10'd169; b_exp2 = 10'd538; b_exp3 = 10'd541;
a_sign0 = 4'd4; a_sign1 = 4'd12; a_sign2 = 4'd14; a_sign3 = 4'd13;
b_sign0 = 4'd7; b_sign1 = 4'd12; b_sign2 = 4'd16; b_sign3 = 4'd1;
@(posedge clk_i);
a_mant0 = 8'd132; a_mant1 = 8'd28; a_mant2 = 8'd78; a_mant3 = 8'd209;
b_mant0 = 8'd242; b_mant1 = 8'd91; b_mant2 = 8'd153; b_mant3 = 8'd23;
a_exp0 = 10'd928; a_exp1 = 10'd395; a_exp2 = 10'd844; a_exp3 = 10'd593;
b_exp0 = 10'd498; b_exp1 = 10'd918; b_exp2 = 10'd39; b_exp3 = 10'd68;
a_sign0 = 4'd12; a_sign1 = 4'd1; a_sign2 = 4'd2; a_sign3 = 4'd8;
b_sign0 = 4'd6; b_sign1 = 4'd11; b_sign2 = 4'd8; b_sign3 = 4'd4;
@(posedge clk_i);
a_mant0 = 8'd172; a_mant1 = 8'd233; a_mant2 = 8'd64; a_mant3 = 8'd137;
b_mant0 = 8'd89; b_mant1 = 8'd142; b_mant2 = 8'd235; b_mant3 = 8'd188;
a_exp0 = 10'd116; a_exp1 = 10'd160; a_exp2 = 10'd151; a_exp3 = 10'd273;
b_exp0 = 10'd750; b_exp1 = 10'd840; b_exp2 = 10'd906; b_exp3 = 10'd815;
a_sign0 = 4'd14; a_sign1 = 4'd2; a_sign2 = 4'd2; a_sign3 = 4'd13;
b_sign0 = 4'd15; b_sign1 = 4'd3; b_sign2 = 4'd10; b_sign3 = 4'd1;
@(posedge clk_i);
a_mant0 = 8'd47; a_mant1 = 8'd37; a_mant2 = 8'd16; a_mant3 = 8'd252;
b_mant0 = 8'd53; b_mant1 = 8'd2; b_mant2 = 8'd151; b_mant3 = 8'd220;
a_exp0 = 10'd865; a_exp1 = 10'd740; a_exp2 = 10'd349; a_exp3 = 10'd836;
b_exp0 = 10'd317; b_exp1 = 10'd169; b_exp2 = 10'd554; b_exp3 = 10'd170;
a_sign0 = 4'd11; a_sign1 = 4'd14; a_sign2 = 4'd15; a_sign3 = 4'd12;
b_sign0 = 4'd14; b_sign1 = 4'd9; b_sign2 = 4'd11; b_sign3 = 4'd9;
@(posedge clk_i);
a_mant0 = 8'd89; a_mant1 = 8'd190; a_mant2 = 8'd143; a_mant3 = 8'd58;
b_mant0 = 8'd231; b_mant1 = 8'd97; b_mant2 = 8'd42; b_mant3 = 8'd146;
a_exp0 = 10'd562; a_exp1 = 10'd742; a_exp2 = 10'd769; a_exp3 = 10'd123;
b_exp0 = 10'd188; b_exp1 = 10'd95; b_exp2 = 10'd80; b_exp3 = 10'd997;
a_sign0 = 4'd10; a_sign1 = 4'd11; a_sign2 = 4'd14; a_sign3 = 4'd15;
b_sign0 = 4'd8; b_sign1 = 4'd1; b_sign2 = 4'd15; b_sign3 = 4'd4;
@(posedge clk_i);
a_mant0 = 8'd83; a_mant1 = 8'd125; a_mant2 = 8'd109; a_mant3 = 8'd50;
b_mant0 = 8'd194; b_mant1 = 8'd138; b_mant2 = 8'd186; b_mant3 = 8'd1;
a_exp0 = 10'd778; a_exp1 = 10'd3; a_exp2 = 10'd309; a_exp3 = 10'd526;
b_exp0 = 10'd857; b_exp1 = 10'd605; b_exp2 = 10'd762; b_exp3 = 10'd667;
a_sign0 = 4'd16; a_sign1 = 4'd16; a_sign2 = 4'd10; a_sign3 = 4'd8;
b_sign0 = 4'd7; b_sign1 = 4'd7; b_sign2 = 4'd3; b_sign3 = 4'd5;
@(posedge clk_i);
a_mant0 = 8'd28; a_mant1 = 8'd93; a_mant2 = 8'd198; a_mant3 = 8'd76;
b_mant0 = 8'd20; b_mant1 = 8'd134; b_mant2 = 8'd100; b_mant3 = 8'd157;
a_exp0 = 10'd749; a_exp1 = 10'd469; a_exp2 = 10'd175; a_exp3 = 10'd341;
b_exp0 = 10'd125; b_exp1 = 10'd384; b_exp2 = 10'd606; b_exp3 = 10'd756;
a_sign0 = 4'd14; a_sign1 = 4'd8; a_sign2 = 4'd14; a_sign3 = 4'd3;
b_sign0 = 4'd8; b_sign1 = 4'd12; b_sign2 = 4'd3; b_sign3 = 4'd0;
@(posedge clk_i);
a_mant0 = 8'd77; a_mant1 = 8'd185; a_mant2 = 8'd3; a_mant3 = 8'd144;
b_mant0 = 8'd105; b_mant1 = 8'd38; b_mant2 = 8'd163; b_mant3 = 8'd39;
a_exp0 = 10'd88; a_exp1 = 10'd987; a_exp2 = 10'd517; a_exp3 = 10'd906;
b_exp0 = 10'd976; b_exp1 = 10'd795; b_exp2 = 10'd601; b_exp3 = 10'd796;
a_sign0 = 4'd10; a_sign1 = 4'd14; a_sign2 = 4'd5; a_sign3 = 4'd14;
b_sign0 = 4'd0; b_sign1 = 4'd16; b_sign2 = 4'd2; b_sign3 = 4'd7;
@(posedge clk_i);
shared_exps0 = 8'd109;
shared_exps1 = 8'd143;
a_mant0 = 8'd158; a_mant1 = 8'd211; a_mant2 = 8'd153; a_mant3 = 8'd208;
b_mant0 = 8'd8; b_mant1 = 8'd16; b_mant2 = 8'd186; b_mant3 = 8'd19;
a_exp0 = 10'd323; a_exp1 = 10'd821; a_exp2 = 10'd306; a_exp3 = 10'd123;
b_exp0 = 10'd157; b_exp1 = 10'd523; b_exp2 = 10'd326; b_exp3 = 10'd261;
a_sign0 = 4'd0; a_sign1 = 4'd15; a_sign2 = 4'd9; a_sign3 = 4'd13;
b_sign0 = 4'd2; b_sign1 = 4'd4; b_sign2 = 4'd0; b_sign3 = 4'd7;
@(posedge clk_i);
a_mant0 = 8'd165; a_mant1 = 8'd223; a_mant2 = 8'd177; a_mant3 = 8'd230;
b_mant0 = 8'd148; b_mant1 = 8'd72; b_mant2 = 8'd0; b_mant3 = 8'd174;
a_exp0 = 10'd678; a_exp1 = 10'd124; a_exp2 = 10'd259; a_exp3 = 10'd518;
b_exp0 = 10'd951; b_exp1 = 10'd149; b_exp2 = 10'd875; b_exp3 = 10'd375;
a_sign0 = 4'd3; a_sign1 = 4'd8; a_sign2 = 4'd14; a_sign3 = 4'd16;
b_sign0 = 4'd10; b_sign1 = 4'd7; b_sign2 = 4'd9; b_sign3 = 4'd9;
@(posedge clk_i);
a_mant0 = 8'd130; a_mant1 = 8'd125; a_mant2 = 8'd91; a_mant3 = 8'd203;
b_mant0 = 8'd91; b_mant1 = 8'd150; b_mant2 = 8'd169; b_mant3 = 8'd148;
a_exp0 = 10'd334; a_exp1 = 10'd219; a_exp2 = 10'd852; a_exp3 = 10'd354;
b_exp0 = 10'd24; b_exp1 = 10'd396; b_exp2 = 10'd310; b_exp3 = 10'd915;
a_sign0 = 4'd14; a_sign1 = 4'd6; a_sign2 = 4'd7; a_sign3 = 4'd12;
b_sign0 = 4'd6; b_sign1 = 4'd4; b_sign2 = 4'd13; b_sign3 = 4'd10;
@(posedge clk_i);
a_mant0 = 8'd30; a_mant1 = 8'd139; a_mant2 = 8'd18; a_mant3 = 8'd169;
b_mant0 = 8'd78; b_mant1 = 8'd82; b_mant2 = 8'd94; b_mant3 = 8'd126;
a_exp0 = 10'd719; a_exp1 = 10'd210; a_exp2 = 10'd696; a_exp3 = 10'd964;
b_exp0 = 10'd666; b_exp1 = 10'd980; b_exp2 = 10'd51; b_exp3 = 10'd629;
a_sign0 = 4'd4; a_sign1 = 4'd10; a_sign2 = 4'd13; a_sign3 = 4'd7;
b_sign0 = 4'd7; b_sign1 = 4'd7; b_sign2 = 4'd2; b_sign3 = 4'd11;
@(posedge clk_i);
a_mant0 = 8'd53; a_mant1 = 8'd216; a_mant2 = 8'd105; a_mant3 = 8'd216;
b_mant0 = 8'd104; b_mant1 = 8'd69; b_mant2 = 8'd113; b_mant3 = 8'd139;
a_exp0 = 10'd83; a_exp1 = 10'd664; a_exp2 = 10'd14; a_exp3 = 10'd794;
b_exp0 = 10'd655; b_exp1 = 10'd214; b_exp2 = 10'd870; b_exp3 = 10'd410;
a_sign0 = 4'd3; a_sign1 = 4'd7; a_sign2 = 4'd11; a_sign3 = 4'd0;
b_sign0 = 4'd3; b_sign1 = 4'd2; b_sign2 = 4'd11; b_sign3 = 4'd3;
@(posedge clk_i);
a_mant0 = 8'd155; a_mant1 = 8'd2; a_mant2 = 8'd14; a_mant3 = 8'd7;
b_mant0 = 8'd70; b_mant1 = 8'd4; b_mant2 = 8'd84; b_mant3 = 8'd168;
a_exp0 = 10'd910; a_exp1 = 10'd822; a_exp2 = 10'd310; a_exp3 = 10'd898;
b_exp0 = 10'd91; b_exp1 = 10'd552; b_exp2 = 10'd276; b_exp3 = 10'd133;
a_sign0 = 4'd14; a_sign1 = 4'd6; a_sign2 = 4'd6; a_sign3 = 4'd13;
b_sign0 = 4'd12; b_sign1 = 4'd3; b_sign2 = 4'd8; b_sign3 = 4'd9;
@(posedge clk_i);
a_mant0 = 8'd129; a_mant1 = 8'd57; a_mant2 = 8'd145; a_mant3 = 8'd163;
b_mant0 = 8'd40; b_mant1 = 8'd63; b_mant2 = 8'd166; b_mant3 = 8'd238;
a_exp0 = 10'd283; a_exp1 = 10'd391; a_exp2 = 10'd111; a_exp3 = 10'd418;
b_exp0 = 10'd612; b_exp1 = 10'd226; b_exp2 = 10'd1003; b_exp3 = 10'd932;
a_sign0 = 4'd13; a_sign1 = 4'd4; a_sign2 = 4'd10; a_sign3 = 4'd0;
b_sign0 = 4'd4; b_sign1 = 4'd4; b_sign2 = 4'd15; b_sign3 = 4'd2;
@(posedge clk_i);
a_mant0 = 8'd149; a_mant1 = 8'd198; a_mant2 = 8'd186; a_mant3 = 8'd111;
b_mant0 = 8'd172; b_mant1 = 8'd216; b_mant2 = 8'd251; b_mant3 = 8'd132;
a_exp0 = 10'd786; a_exp1 = 10'd700; a_exp2 = 10'd1010; a_exp3 = 10'd463;
b_exp0 = 10'd97; b_exp1 = 10'd653; b_exp2 = 10'd964; b_exp3 = 10'd425;
a_sign0 = 4'd12; a_sign1 = 4'd10; a_sign2 = 4'd11; a_sign3 = 4'd10;
b_sign0 = 4'd15; b_sign1 = 4'd13; b_sign2 = 4'd16; b_sign3 = 4'd7;
@(posedge clk_i);
shared_exps0 = 8'd133;
shared_exps1 = 8'd79;
rstn = 0;
@(posedge clk_i);
rstn = 1;
a_mant0 = 8'd243; a_mant1 = 8'd172; a_mant2 = 8'd154; a_mant3 = 8'd211;
b_mant0 = 8'd182; b_mant1 = 8'd99; b_mant2 = 8'd14; b_mant3 = 8'd117;
a_exp0 = 10'd625; a_exp1 = 10'd539; a_exp2 = 10'd350; a_exp3 = 10'd343;
b_exp0 = 10'd760; b_exp1 = 10'd188; b_exp2 = 10'd312; b_exp3 = 10'd390;
a_sign0 = 4'd5; a_sign1 = 4'd15; a_sign2 = 4'd1; a_sign3 = 4'd13;
b_sign0 = 4'd12; b_sign1 = 4'd15; b_sign2 = 4'd4; b_sign3 = 4'd6;
@(posedge clk_i);
a_mant0 = 8'd196; a_mant1 = 8'd160; a_mant2 = 8'd7; a_mant3 = 8'd108;
b_mant0 = 8'd139; b_mant1 = 8'd16; b_mant2 = 8'd35; b_mant3 = 8'd128;
a_exp0 = 10'd956; a_exp1 = 10'd723; a_exp2 = 10'd408; a_exp3 = 10'd456;
b_exp0 = 10'd409; b_exp1 = 10'd265; b_exp2 = 10'd468; b_exp3 = 10'd782;
a_sign0 = 4'd10; a_sign1 = 4'd1; a_sign2 = 4'd3; a_sign3 = 4'd0;
b_sign0 = 4'd4; b_sign1 = 4'd13; b_sign2 = 4'd16; b_sign3 = 4'd9;
@(posedge clk_i);
a_mant0 = 8'd194; a_mant1 = 8'd199; a_mant2 = 8'd201; a_mant3 = 8'd198;
b_mant0 = 8'd200; b_mant1 = 8'd73; b_mant2 = 8'd14; b_mant3 = 8'd146;
a_exp0 = 10'd720; a_exp1 = 10'd879; a_exp2 = 10'd378; a_exp3 = 10'd930;
b_exp0 = 10'd743; b_exp1 = 10'd528; b_exp2 = 10'd138; b_exp3 = 10'd486;
a_sign0 = 4'd5; a_sign1 = 4'd11; a_sign2 = 4'd4; a_sign3 = 4'd3;
b_sign0 = 4'd7; b_sign1 = 4'd4; b_sign2 = 4'd6; b_sign3 = 4'd11;
@(posedge clk_i);
a_mant0 = 8'd121; a_mant1 = 8'd142; a_mant2 = 8'd190; a_mant3 = 8'd50;
b_mant0 = 8'd183; b_mant1 = 8'd186; b_mant2 = 8'd238; b_mant3 = 8'd82;
a_exp0 = 10'd823; a_exp1 = 10'd470; a_exp2 = 10'd186; a_exp3 = 10'd882;
b_exp0 = 10'd39; b_exp1 = 10'd48; b_exp2 = 10'd965; b_exp3 = 10'd433;
a_sign0 = 4'd2; a_sign1 = 4'd4; a_sign2 = 4'd3; a_sign3 = 4'd6;
b_sign0 = 4'd1; b_sign1 = 4'd16; b_sign2 = 4'd6; b_sign3 = 4'd1;
@(posedge clk_i);
a_mant0 = 8'd28; a_mant1 = 8'd10; a_mant2 = 8'd244; a_mant3 = 8'd44;
b_mant0 = 8'd191; b_mant1 = 8'd154; b_mant2 = 8'd253; b_mant3 = 8'd168;
a_exp0 = 10'd442; a_exp1 = 10'd1016; a_exp2 = 10'd35; a_exp3 = 10'd631;
b_exp0 = 10'd347; b_exp1 = 10'd73; b_exp2 = 10'd686; b_exp3 = 10'd33;
a_sign0 = 4'd8; a_sign1 = 4'd6; a_sign2 = 4'd12; a_sign3 = 4'd10;
b_sign0 = 4'd1; b_sign1 = 4'd4; b_sign2 = 4'd7; b_sign3 = 4'd7;
@(posedge clk_i);
a_mant0 = 8'd216; a_mant1 = 8'd18; a_mant2 = 8'd72; a_mant3 = 8'd213;
b_mant0 = 8'd201; b_mant1 = 8'd199; b_mant2 = 8'd105; b_mant3 = 8'd196;
a_exp0 = 10'd624; a_exp1 = 10'd709; a_exp2 = 10'd813; a_exp3 = 10'd914;
b_exp0 = 10'd374; b_exp1 = 10'd697; b_exp2 = 10'd879; b_exp3 = 10'd482;
a_sign0 = 4'd16; a_sign1 = 4'd13; a_sign2 = 4'd7; a_sign3 = 4'd5;
b_sign0 = 4'd13; b_sign1 = 4'd4; b_sign2 = 4'd4; b_sign3 = 4'd1;
@(posedge clk_i);
a_mant0 = 8'd168; a_mant1 = 8'd196; a_mant2 = 8'd199; a_mant3 = 8'd129;
b_mant0 = 8'd93; b_mant1 = 8'd64; b_mant2 = 8'd73; b_mant3 = 8'd114;
a_exp0 = 10'd139; a_exp1 = 10'd782; a_exp2 = 10'd427; a_exp3 = 10'd319;
b_exp0 = 10'd306; b_exp1 = 10'd603; b_exp2 = 10'd324; b_exp3 = 10'd248;
a_sign0 = 4'd7; a_sign1 = 4'd8; a_sign2 = 4'd11; a_sign3 = 4'd2;
b_sign0 = 4'd10; b_sign1 = 4'd3; b_sign2 = 4'd9; b_sign3 = 4'd10;
@(posedge clk_i);
shared_exps0 = 8'd149;
shared_exps1 = 8'd111;
a_mant0 = 8'd209; a_mant1 = 8'd116; a_mant2 = 8'd116; a_mant3 = 8'd175;
b_mant0 = 8'd5; b_mant1 = 8'd237; b_mant2 = 8'd15; b_mant3 = 8'd40;
a_exp0 = 10'd207; a_exp1 = 10'd778; a_exp2 = 10'd456; a_exp3 = 10'd411;
b_exp0 = 10'd693; b_exp1 = 10'd24; b_exp2 = 10'd192; b_exp3 = 10'd421;
a_sign0 = 4'd7; a_sign1 = 4'd14; a_sign2 = 4'd4; a_sign3 = 4'd4;
b_sign0 = 4'd16; b_sign1 = 4'd5; b_sign2 = 4'd4; b_sign3 = 4'd6;
@(posedge clk_i);
a_mant0 = 8'd51; a_mant1 = 8'd86; a_mant2 = 8'd228; a_mant3 = 8'd233;
b_mant0 = 8'd137; b_mant1 = 8'd153; b_mant2 = 8'd212; b_mant3 = 8'd32;
a_exp0 = 10'd725; a_exp1 = 10'd735; a_exp2 = 10'd924; a_exp3 = 10'd185;
b_exp0 = 10'd311; b_exp1 = 10'd782; b_exp2 = 10'd5; b_exp3 = 10'd621;
a_sign0 = 4'd12; a_sign1 = 4'd2; a_sign2 = 4'd9; a_sign3 = 4'd12;
b_sign0 = 4'd5; b_sign1 = 4'd9; b_sign2 = 4'd8; b_sign3 = 4'd11;
@(posedge clk_i);
a_mant0 = 8'd108; a_mant1 = 8'd186; a_mant2 = 8'd129; a_mant3 = 8'd185;
b_mant0 = 8'd250; b_mant1 = 8'd98; b_mant2 = 8'd182; b_mant3 = 8'd24;
a_exp0 = 10'd350; a_exp1 = 10'd536; a_exp2 = 10'd548; a_exp3 = 10'd826;
b_exp0 = 10'd483; b_exp1 = 10'd374; b_exp2 = 10'd641; b_exp3 = 10'd550;
a_sign0 = 4'd4; a_sign1 = 4'd15; a_sign2 = 4'd3; a_sign3 = 4'd0;
b_sign0 = 4'd1; b_sign1 = 4'd12; b_sign2 = 4'd13; b_sign3 = 4'd7;
@(posedge clk_i);
a_mant0 = 8'd77; a_mant1 = 8'd170; a_mant2 = 8'd144; a_mant3 = 8'd218;
b_mant0 = 8'd117; b_mant1 = 8'd108; b_mant2 = 8'd226; b_mant3 = 8'd75;
a_exp0 = 10'd583; a_exp1 = 10'd369; a_exp2 = 10'd131; a_exp3 = 10'd844;
b_exp0 = 10'd641; b_exp1 = 10'd27; b_exp2 = 10'd958; b_exp3 = 10'd293;
a_sign0 = 4'd9; a_sign1 = 4'd3; a_sign2 = 4'd7; a_sign3 = 4'd16;
b_sign0 = 4'd14; b_sign1 = 4'd13; b_sign2 = 4'd5; b_sign3 = 4'd13;
@(posedge clk_i);
a_mant0 = 8'd145; a_mant1 = 8'd81; a_mant2 = 8'd235; a_mant3 = 8'd237;
b_mant0 = 8'd231; b_mant1 = 8'd29; b_mant2 = 8'd194; b_mant3 = 8'd64;
a_exp0 = 10'd120; a_exp1 = 10'd534; a_exp2 = 10'd932; a_exp3 = 10'd685;
b_exp0 = 10'd907; b_exp1 = 10'd374; b_exp2 = 10'd296; b_exp3 = 10'd493;
a_sign0 = 4'd11; a_sign1 = 4'd10; a_sign2 = 4'd1; a_sign3 = 4'd15;
b_sign0 = 4'd10; b_sign1 = 4'd9; b_sign2 = 4'd2; b_sign3 = 4'd8;
@(posedge clk_i);
a_mant0 = 8'd122; a_mant1 = 8'd22; a_mant2 = 8'd67; a_mant3 = 8'd197;
b_mant0 = 8'd201; b_mant1 = 8'd205; b_mant2 = 8'd28; b_mant3 = 8'd245;
a_exp0 = 10'd467; a_exp1 = 10'd909; a_exp2 = 10'd1011; a_exp3 = 10'd172;
b_exp0 = 10'd401; b_exp1 = 10'd231; b_exp2 = 10'd259; b_exp3 = 10'd778;
a_sign0 = 4'd8; a_sign1 = 4'd12; a_sign2 = 4'd8; a_sign3 = 4'd8;
b_sign0 = 4'd3; b_sign1 = 4'd15; b_sign2 = 4'd9; b_sign3 = 4'd10;
@(posedge clk_i);
a_mant0 = 8'd102; a_mant1 = 8'd30; a_mant2 = 8'd166; a_mant3 = 8'd215;
b_mant0 = 8'd173; b_mant1 = 8'd137; b_mant2 = 8'd50; b_mant3 = 8'd128;
a_exp0 = 10'd85; a_exp1 = 10'd440; a_exp2 = 10'd641; a_exp3 = 10'd580;
b_exp0 = 10'd315; b_exp1 = 10'd505; b_exp2 = 10'd97; b_exp3 = 10'd116;
a_sign0 = 4'd7; a_sign1 = 4'd4; a_sign2 = 4'd10; a_sign3 = 4'd2;
b_sign0 = 4'd10; b_sign1 = 4'd15; b_sign2 = 4'd0; b_sign3 = 4'd8;
@(posedge clk_i);
a_mant0 = 8'd159; a_mant1 = 8'd47; a_mant2 = 8'd148; a_mant3 = 8'd76;
b_mant0 = 8'd232; b_mant1 = 8'd99; b_mant2 = 8'd80; b_mant3 = 8'd70;
a_exp0 = 10'd224; a_exp1 = 10'd331; a_exp2 = 10'd773; a_exp3 = 10'd983;
b_exp0 = 10'd860; b_exp1 = 10'd186; b_exp2 = 10'd156; b_exp3 = 10'd869;
a_sign0 = 4'd13; a_sign1 = 4'd4; a_sign2 = 4'd7; a_sign3 = 4'd16;
b_sign0 = 4'd11; b_sign1 = 4'd7; b_sign2 = 4'd4; b_sign3 = 4'd0;
@(posedge clk_i);
shared_exps0 = 8'd125;
shared_exps1 = 8'd141;
a_mant0 = 8'd248; a_mant1 = 8'd48; a_mant2 = 8'd19; a_mant3 = 8'd20;
b_mant0 = 8'd64; b_mant1 = 8'd90; b_mant2 = 8'd187; b_mant3 = 8'd68;
a_exp0 = 10'd345; a_exp1 = 10'd762; a_exp2 = 10'd785; a_exp3 = 10'd174;
b_exp0 = 10'd623; b_exp1 = 10'd819; b_exp2 = 10'd267; b_exp3 = 10'd973;
a_sign0 = 4'd14; a_sign1 = 4'd2; a_sign2 = 4'd2; a_sign3 = 4'd3;
b_sign0 = 4'd10; b_sign1 = 4'd10; b_sign2 = 4'd1; b_sign3 = 4'd4;
@(posedge clk_i);
a_mant0 = 8'd52; a_mant1 = 8'd199; a_mant2 = 8'd95; a_mant3 = 8'd75;
b_mant0 = 8'd125; b_mant1 = 8'd241; b_mant2 = 8'd103; b_mant3 = 8'd48;
a_exp0 = 10'd286; a_exp1 = 10'd734; a_exp2 = 10'd994; a_exp3 = 10'd637;
b_exp0 = 10'd201; b_exp1 = 10'd580; b_exp2 = 10'd898; b_exp3 = 10'd2;
a_sign0 = 4'd6; a_sign1 = 4'd7; a_sign2 = 4'd0; a_sign3 = 4'd16;
b_sign0 = 4'd6; b_sign1 = 4'd11; b_sign2 = 4'd16; b_sign3 = 4'd16;
@(posedge clk_i);
a_mant0 = 8'd187; a_mant1 = 8'd102; a_mant2 = 8'd164; a_mant3 = 8'd156;
b_mant0 = 8'd36; b_mant1 = 8'd247; b_mant2 = 8'd55; b_mant3 = 8'd22;
a_exp0 = 10'd21; a_exp1 = 10'd140; a_exp2 = 10'd485; a_exp3 = 10'd396;
b_exp0 = 10'd991; b_exp1 = 10'd577; b_exp2 = 10'd315; b_exp3 = 10'd985;
a_sign0 = 4'd7; a_sign1 = 4'd13; a_sign2 = 4'd10; a_sign3 = 4'd3;
b_sign0 = 4'd1; b_sign1 = 4'd11; b_sign2 = 4'd4; b_sign3 = 4'd8;
@(posedge clk_i);
a_mant0 = 8'd94; a_mant1 = 8'd31; a_mant2 = 8'd8; a_mant3 = 8'd206;
b_mant0 = 8'd99; b_mant1 = 8'd205; b_mant2 = 8'd37; b_mant3 = 8'd39;
a_exp0 = 10'd988; a_exp1 = 10'd806; a_exp2 = 10'd800; a_exp3 = 10'd687;
b_exp0 = 10'd843; b_exp1 = 10'd27; b_exp2 = 10'd743; b_exp3 = 10'd882;
a_sign0 = 4'd13; a_sign1 = 4'd8; a_sign2 = 4'd16; a_sign3 = 4'd8;
b_sign0 = 4'd2; b_sign1 = 4'd1; b_sign2 = 4'd2; b_sign3 = 4'd14;
@(posedge clk_i);
a_mant0 = 8'd57; a_mant1 = 8'd63; a_mant2 = 8'd230; a_mant3 = 8'd249;
b_mant0 = 8'd37; b_mant1 = 8'd165; b_mant2 = 8'd155; b_mant3 = 8'd230;
a_exp0 = 10'd877; a_exp1 = 10'd46; a_exp2 = 10'd975; a_exp3 = 10'd766;
b_exp0 = 10'd50; b_exp1 = 10'd369; b_exp2 = 10'd673; b_exp3 = 10'd976;
a_sign0 = 4'd2; a_sign1 = 4'd13; a_sign2 = 4'd11; a_sign3 = 4'd1;
b_sign0 = 4'd0; b_sign1 = 4'd10; b_sign2 = 4'd10; b_sign3 = 4'd16;
@(posedge clk_i);
a_mant0 = 8'd115; a_mant1 = 8'd31; a_mant2 = 8'd64; a_mant3 = 8'd180;
b_mant0 = 8'd29; b_mant1 = 8'd183; b_mant2 = 8'd121; b_mant3 = 8'd1;
a_exp0 = 10'd276; a_exp1 = 10'd460; a_exp2 = 10'd304; a_exp3 = 10'd216;
b_exp0 = 10'd439; b_exp1 = 10'd583; b_exp2 = 10'd424; b_exp3 = 10'd469;
a_sign0 = 4'd2; a_sign1 = 4'd2; a_sign2 = 4'd2; a_sign3 = 4'd10;
b_sign0 = 4'd1; b_sign1 = 4'd2; b_sign2 = 4'd11; b_sign3 = 4'd16;
@(posedge clk_i);
a_mant0 = 8'd161; a_mant1 = 8'd93; a_mant2 = 8'd66; a_mant3 = 8'd203;
b_mant0 = 8'd102; b_mant1 = 8'd105; b_mant2 = 8'd153; b_mant3 = 8'd134;
a_exp0 = 10'd951; a_exp1 = 10'd371; a_exp2 = 10'd594; a_exp3 = 10'd385;
b_exp0 = 10'd502; b_exp1 = 10'd797; b_exp2 = 10'd155; b_exp3 = 10'd383;
a_sign0 = 4'd12; a_sign1 = 4'd9; a_sign2 = 4'd9; a_sign3 = 4'd10;
b_sign0 = 4'd1; b_sign1 = 4'd2; b_sign2 = 4'd5; b_sign3 = 4'd8;
@(posedge clk_i);
a_mant0 = 8'd171; a_mant1 = 8'd140; a_mant2 = 8'd222; a_mant3 = 8'd62;
b_mant0 = 8'd248; b_mant1 = 8'd126; b_mant2 = 8'd144; b_mant3 = 8'd195;
a_exp0 = 10'd105; a_exp1 = 10'd354; a_exp2 = 10'd805; a_exp3 = 10'd102;
b_exp0 = 10'd23; b_exp1 = 10'd393; b_exp2 = 10'd412; b_exp3 = 10'd758;
a_sign0 = 4'd3; a_sign1 = 4'd0; a_sign2 = 4'd14; a_sign3 = 4'd8;
b_sign0 = 4'd5; b_sign1 = 4'd0; b_sign2 = 4'd10; b_sign3 = 4'd9;
@(posedge clk_i);
shared_exps0 = 8'd146;
shared_exps1 = 8'd115;
a_mant0 = 8'd216; a_mant1 = 8'd87; a_mant2 = 8'd185; a_mant3 = 8'd196;
b_mant0 = 8'd236; b_mant1 = 8'd95; b_mant2 = 8'd98; b_mant3 = 8'd224;
a_exp0 = 10'd571; a_exp1 = 10'd58; a_exp2 = 10'd633; a_exp3 = 10'd126;
b_exp0 = 10'd645; b_exp1 = 10'd154; b_exp2 = 10'd358; b_exp3 = 10'd777;
a_sign0 = 4'd9; a_sign1 = 4'd9; a_sign2 = 4'd16; a_sign3 = 4'd13;
b_sign0 = 4'd11; b_sign1 = 4'd15; b_sign2 = 4'd7; b_sign3 = 4'd5;
@(posedge clk_i);
a_mant0 = 8'd148; a_mant1 = 8'd252; a_mant2 = 8'd21; a_mant3 = 8'd122;
b_mant0 = 8'd88; b_mant1 = 8'd30; b_mant2 = 8'd75; b_mant3 = 8'd44;
a_exp0 = 10'd506; a_exp1 = 10'd660; a_exp2 = 10'd105; a_exp3 = 10'd455;
b_exp0 = 10'd389; b_exp1 = 10'd64; b_exp2 = 10'd734; b_exp3 = 10'd446;
a_sign0 = 4'd6; a_sign1 = 4'd2; a_sign2 = 4'd1; a_sign3 = 4'd11;
b_sign0 = 4'd2; b_sign1 = 4'd14; b_sign2 = 4'd2; b_sign3 = 4'd2;
@(posedge clk_i);
a_mant0 = 8'd75; a_mant1 = 8'd28; a_mant2 = 8'd185; a_mant3 = 8'd64;
b_mant0 = 8'd219; b_mant1 = 8'd215; b_mant2 = 8'd239; b_mant3 = 8'd86;
a_exp0 = 10'd945; a_exp1 = 10'd927; a_exp2 = 10'd241; a_exp3 = 10'd938;
b_exp0 = 10'd725; b_exp1 = 10'd184; b_exp2 = 10'd1000; b_exp3 = 10'd517;
a_sign0 = 4'd15; a_sign1 = 4'd3; a_sign2 = 4'd4; a_sign3 = 4'd3;
b_sign0 = 4'd9; b_sign1 = 4'd0; b_sign2 = 4'd0; b_sign3 = 4'd8;
@(posedge clk_i);
a_mant0 = 8'd71; a_mant1 = 8'd112; a_mant2 = 8'd85; a_mant3 = 8'd164;
b_mant0 = 8'd21; b_mant1 = 8'd33; b_mant2 = 8'd133; b_mant3 = 8'd199;
a_exp0 = 10'd626; a_exp1 = 10'd529; a_exp2 = 10'd324; a_exp3 = 10'd67;
b_exp0 = 10'd535; b_exp1 = 10'd637; b_exp2 = 10'd401; b_exp3 = 10'd718;
a_sign0 = 4'd6; a_sign1 = 4'd4; a_sign2 = 4'd9; a_sign3 = 4'd4;
b_sign0 = 4'd13; b_sign1 = 4'd16; b_sign2 = 4'd9; b_sign3 = 4'd8;
@(posedge clk_i);
a_mant0 = 8'd67; a_mant1 = 8'd113; a_mant2 = 8'd231; a_mant3 = 8'd28;
b_mant0 = 8'd50; b_mant1 = 8'd191; b_mant2 = 8'd169; b_mant3 = 8'd250;
a_exp0 = 10'd273; a_exp1 = 10'd867; a_exp2 = 10'd427; a_exp3 = 10'd562;
b_exp0 = 10'd188; b_exp1 = 10'd985; b_exp2 = 10'd931; b_exp3 = 10'd426;
a_sign0 = 4'd3; a_sign1 = 4'd13; a_sign2 = 4'd10; a_sign3 = 4'd6;
b_sign0 = 4'd11; b_sign1 = 4'd2; b_sign2 = 4'd14; b_sign3 = 4'd5;
@(posedge clk_i);
a_mant0 = 8'd236; a_mant1 = 8'd220; a_mant2 = 8'd47; a_mant3 = 8'd251;
b_mant0 = 8'd44; b_mant1 = 8'd48; b_mant2 = 8'd114; b_mant3 = 8'd17;
a_exp0 = 10'd752; a_exp1 = 10'd830; a_exp2 = 10'd353; a_exp3 = 10'd287;
b_exp0 = 10'd343; b_exp1 = 10'd811; b_exp2 = 10'd746; b_exp3 = 10'd590;
a_sign0 = 4'd10; a_sign1 = 4'd6; a_sign2 = 4'd0; a_sign3 = 4'd0;
b_sign0 = 4'd13; b_sign1 = 4'd5; b_sign2 = 4'd12; b_sign3 = 4'd6;
@(posedge clk_i);
a_mant0 = 8'd4; a_mant1 = 8'd179; a_mant2 = 8'd235; a_mant3 = 8'd117;
b_mant0 = 8'd141; b_mant1 = 8'd31; b_mant2 = 8'd184; b_mant3 = 8'd143;
a_exp0 = 10'd453; a_exp1 = 10'd955; a_exp2 = 10'd64; a_exp3 = 10'd355;
b_exp0 = 10'd938; b_exp1 = 10'd997; b_exp2 = 10'd63; b_exp3 = 10'd69;
a_sign0 = 4'd0; a_sign1 = 4'd10; a_sign2 = 4'd3; a_sign3 = 4'd12;
b_sign0 = 4'd2; b_sign1 = 4'd12; b_sign2 = 4'd0; b_sign3 = 4'd14;
@(posedge clk_i);
a_mant0 = 8'd199; a_mant1 = 8'd183; a_mant2 = 8'd75; a_mant3 = 8'd225;
b_mant0 = 8'd45; b_mant1 = 8'd38; b_mant2 = 8'd123; b_mant3 = 8'd93;
a_exp0 = 10'd618; a_exp1 = 10'd471; a_exp2 = 10'd1017; a_exp3 = 10'd790;
b_exp0 = 10'd513; b_exp1 = 10'd165; b_exp2 = 10'd21; b_exp3 = 10'd733;
a_sign0 = 4'd12; a_sign1 = 4'd16; a_sign2 = 4'd12; a_sign3 = 4'd7;
b_sign0 = 4'd13; b_sign1 = 4'd7; b_sign2 = 4'd11; b_sign3 = 4'd10;
@(posedge clk_i);
shared_exps0 = 8'd104;
shared_exps1 = 8'd115;
rstn = 0;
@(posedge clk_i);
rstn = 1;
a_mant0 = 8'd176; a_mant1 = 8'd0; a_mant2 = 8'd142; a_mant3 = 8'd2;
b_mant0 = 8'd164; b_mant1 = 8'd206; b_mant2 = 8'd136; b_mant3 = 8'd16;
a_exp0 = 10'd464; a_exp1 = 10'd53; a_exp2 = 10'd375; a_exp3 = 10'd798;
b_exp0 = 10'd804; b_exp1 = 10'd405; b_exp2 = 10'd778; b_exp3 = 10'd602;
a_sign0 = 4'd8; a_sign1 = 4'd7; a_sign2 = 4'd14; a_sign3 = 4'd7;
b_sign0 = 4'd13; b_sign1 = 4'd3; b_sign2 = 4'd12; b_sign3 = 4'd0;
@(posedge clk_i);
a_mant0 = 8'd157; a_mant1 = 8'd112; a_mant2 = 8'd161; a_mant3 = 8'd26;
b_mant0 = 8'd144; b_mant1 = 8'd80; b_mant2 = 8'd164; b_mant3 = 8'd122;
a_exp0 = 10'd340; a_exp1 = 10'd247; a_exp2 = 10'd623; a_exp3 = 10'd690;
b_exp0 = 10'd302; b_exp1 = 10'd755; b_exp2 = 10'd904; b_exp3 = 10'd1011;
a_sign0 = 4'd2; a_sign1 = 4'd16; a_sign2 = 4'd5; a_sign3 = 4'd9;
b_sign0 = 4'd16; b_sign1 = 4'd0; b_sign2 = 4'd1; b_sign3 = 4'd0;
@(posedge clk_i);
a_mant0 = 8'd19; a_mant1 = 8'd162; a_mant2 = 8'd191; a_mant3 = 8'd120;
b_mant0 = 8'd182; b_mant1 = 8'd87; b_mant2 = 8'd159; b_mant3 = 8'd219;
a_exp0 = 10'd322; a_exp1 = 10'd670; a_exp2 = 10'd45; a_exp3 = 10'd1018;
b_exp0 = 10'd680; b_exp1 = 10'd147; b_exp2 = 10'd601; b_exp3 = 10'd810;
a_sign0 = 4'd5; a_sign1 = 4'd3; a_sign2 = 4'd12; a_sign3 = 4'd12;
b_sign0 = 4'd4; b_sign1 = 4'd3; b_sign2 = 4'd9; b_sign3 = 4'd4;
@(posedge clk_i);
a_mant0 = 8'd48; a_mant1 = 8'd193; a_mant2 = 8'd56; a_mant3 = 8'd81;
b_mant0 = 8'd14; b_mant1 = 8'd227; b_mant2 = 8'd3; b_mant3 = 8'd127;
a_exp0 = 10'd132; a_exp1 = 10'd980; a_exp2 = 10'd398; a_exp3 = 10'd670;
b_exp0 = 10'd76; b_exp1 = 10'd464; b_exp2 = 10'd278; b_exp3 = 10'd410;
a_sign0 = 4'd8; a_sign1 = 4'd2; a_sign2 = 4'd15; a_sign3 = 4'd3;
b_sign0 = 4'd12; b_sign1 = 4'd10; b_sign2 = 4'd9; b_sign3 = 4'd12;
@(posedge clk_i);
a_mant0 = 8'd86; a_mant1 = 8'd21; a_mant2 = 8'd1; a_mant3 = 8'd160;
b_mant0 = 8'd125; b_mant1 = 8'd235; b_mant2 = 8'd189; b_mant3 = 8'd254;
a_exp0 = 10'd668; a_exp1 = 10'd393; a_exp2 = 10'd689; a_exp3 = 10'd832;
b_exp0 = 10'd118; b_exp1 = 10'd500; b_exp2 = 10'd357; b_exp3 = 10'd721;
a_sign0 = 4'd13; a_sign1 = 4'd8; a_sign2 = 4'd0; a_sign3 = 4'd16;
b_sign0 = 4'd0; b_sign1 = 4'd15; b_sign2 = 4'd8; b_sign3 = 4'd3;
@(posedge clk_i);
a_mant0 = 8'd139; a_mant1 = 8'd237; a_mant2 = 8'd108; a_mant3 = 8'd62;
b_mant0 = 8'd25; b_mant1 = 8'd60; b_mant2 = 8'd186; b_mant3 = 8'd115;
a_exp0 = 10'd402; a_exp1 = 10'd155; a_exp2 = 10'd249; a_exp3 = 10'd560;
b_exp0 = 10'd346; b_exp1 = 10'd559; b_exp2 = 10'd56; b_exp3 = 10'd742;
a_sign0 = 4'd11; a_sign1 = 4'd1; a_sign2 = 4'd9; a_sign3 = 4'd11;
b_sign0 = 4'd1; b_sign1 = 4'd0; b_sign2 = 4'd8; b_sign3 = 4'd14;
@(posedge clk_i);
a_mant0 = 8'd28; a_mant1 = 8'd165; a_mant2 = 8'd8; a_mant3 = 8'd225;
b_mant0 = 8'd119; b_mant1 = 8'd23; b_mant2 = 8'd171; b_mant3 = 8'd185;
a_exp0 = 10'd553; a_exp1 = 10'd282; a_exp2 = 10'd609; a_exp3 = 10'd476;
b_exp0 = 10'd1011; b_exp1 = 10'd269; b_exp2 = 10'd765; b_exp3 = 10'd394;
a_sign0 = 4'd6; a_sign1 = 4'd4; a_sign2 = 4'd9; a_sign3 = 4'd11;
b_sign0 = 4'd5; b_sign1 = 4'd4; b_sign2 = 4'd6; b_sign3 = 4'd11;
@(posedge clk_i);
shared_exps0 = 8'd141;
shared_exps1 = 8'd101;
a_mant0 = 8'd195; a_mant1 = 8'd13; a_mant2 = 8'd168; a_mant3 = 8'd96;
b_mant0 = 8'd133; b_mant1 = 8'd42; b_mant2 = 8'd32; b_mant3 = 8'd106;
a_exp0 = 10'd389; a_exp1 = 10'd944; a_exp2 = 10'd901; a_exp3 = 10'd907;
b_exp0 = 10'd583; b_exp1 = 10'd346; b_exp2 = 10'd349; b_exp3 = 10'd552;
a_sign0 = 4'd2; a_sign1 = 4'd10; a_sign2 = 4'd6; a_sign3 = 4'd12;
b_sign0 = 4'd8; b_sign1 = 4'd2; b_sign2 = 4'd3; b_sign3 = 4'd4;
@(posedge clk_i);
a_mant0 = 8'd169; a_mant1 = 8'd207; a_mant2 = 8'd73; a_mant3 = 8'd119;
b_mant0 = 8'd130; b_mant1 = 8'd49; b_mant2 = 8'd219; b_mant3 = 8'd52;
a_exp0 = 10'd630; a_exp1 = 10'd102; a_exp2 = 10'd741; a_exp3 = 10'd625;
b_exp0 = 10'd218; b_exp1 = 10'd422; b_exp2 = 10'd57; b_exp3 = 10'd831;
a_sign0 = 4'd15; a_sign1 = 4'd16; a_sign2 = 4'd9; a_sign3 = 4'd0;
b_sign0 = 4'd11; b_sign1 = 4'd10; b_sign2 = 4'd7; b_sign3 = 4'd3;
@(posedge clk_i);
a_mant0 = 8'd73; a_mant1 = 8'd45; a_mant2 = 8'd99; a_mant3 = 8'd81;
b_mant0 = 8'd10; b_mant1 = 8'd243; b_mant2 = 8'd50; b_mant3 = 8'd13;
a_exp0 = 10'd843; a_exp1 = 10'd552; a_exp2 = 10'd487; a_exp3 = 10'd994;
b_exp0 = 10'd11; b_exp1 = 10'd969; b_exp2 = 10'd503; b_exp3 = 10'd181;
a_sign0 = 4'd8; a_sign1 = 4'd5; a_sign2 = 4'd15; a_sign3 = 4'd3;
b_sign0 = 4'd6; b_sign1 = 4'd12; b_sign2 = 4'd13; b_sign3 = 4'd0;
@(posedge clk_i);
a_mant0 = 8'd59; a_mant1 = 8'd17; a_mant2 = 8'd112; a_mant3 = 8'd9;
b_mant0 = 8'd209; b_mant1 = 8'd62; b_mant2 = 8'd51; b_mant3 = 8'd242;
a_exp0 = 10'd64; a_exp1 = 10'd118; a_exp2 = 10'd34; a_exp3 = 10'd822;
b_exp0 = 10'd766; b_exp1 = 10'd719; b_exp2 = 10'd471; b_exp3 = 10'd100;
a_sign0 = 4'd11; a_sign1 = 4'd6; a_sign2 = 4'd12; a_sign3 = 4'd3;
b_sign0 = 4'd10; b_sign1 = 4'd10; b_sign2 = 4'd11; b_sign3 = 4'd5;
@(posedge clk_i);
a_mant0 = 8'd38; a_mant1 = 8'd161; a_mant2 = 8'd235; a_mant3 = 8'd117;
b_mant0 = 8'd242; b_mant1 = 8'd8; b_mant2 = 8'd142; b_mant3 = 8'd55;
a_exp0 = 10'd163; a_exp1 = 10'd994; a_exp2 = 10'd562; a_exp3 = 10'd886;
b_exp0 = 10'd482; b_exp1 = 10'd650; b_exp2 = 10'd446; b_exp3 = 10'd838;
a_sign0 = 4'd7; a_sign1 = 4'd10; a_sign2 = 4'd13; a_sign3 = 4'd1;
b_sign0 = 4'd8; b_sign1 = 4'd7; b_sign2 = 4'd11; b_sign3 = 4'd9;
@(posedge clk_i);
a_mant0 = 8'd53; a_mant1 = 8'd124; a_mant2 = 8'd229; a_mant3 = 8'd11;
b_mant0 = 8'd219; b_mant1 = 8'd200; b_mant2 = 8'd68; b_mant3 = 8'd9;
a_exp0 = 10'd325; a_exp1 = 10'd522; a_exp2 = 10'd345; a_exp3 = 10'd58;
b_exp0 = 10'd592; b_exp1 = 10'd692; b_exp2 = 10'd250; b_exp3 = 10'd774;
a_sign0 = 4'd15; a_sign1 = 4'd2; a_sign2 = 4'd12; a_sign3 = 4'd10;
b_sign0 = 4'd5; b_sign1 = 4'd14; b_sign2 = 4'd5; b_sign3 = 4'd11;
@(posedge clk_i);
a_mant0 = 8'd199; a_mant1 = 8'd163; a_mant2 = 8'd212; a_mant3 = 8'd154;
b_mant0 = 8'd36; b_mant1 = 8'd208; b_mant2 = 8'd239; b_mant3 = 8'd62;
a_exp0 = 10'd931; a_exp1 = 10'd381; a_exp2 = 10'd1016; a_exp3 = 10'd52;
b_exp0 = 10'd682; b_exp1 = 10'd762; b_exp2 = 10'd984; b_exp3 = 10'd451;
a_sign0 = 4'd1; a_sign1 = 4'd2; a_sign2 = 4'd2; a_sign3 = 4'd5;
b_sign0 = 4'd0; b_sign1 = 4'd3; b_sign2 = 4'd4; b_sign3 = 4'd4;
@(posedge clk_i);
a_mant0 = 8'd173; a_mant1 = 8'd139; a_mant2 = 8'd39; a_mant3 = 8'd168;
b_mant0 = 8'd13; b_mant1 = 8'd253; b_mant2 = 8'd41; b_mant3 = 8'd78;
a_exp0 = 10'd49; a_exp1 = 10'd113; a_exp2 = 10'd491; a_exp3 = 10'd74;
b_exp0 = 10'd220; b_exp1 = 10'd94; b_exp2 = 10'd826; b_exp3 = 10'd326;
a_sign0 = 4'd12; a_sign1 = 4'd4; a_sign2 = 4'd8; a_sign3 = 4'd13;
b_sign0 = 4'd3; b_sign1 = 4'd0; b_sign2 = 4'd5; b_sign3 = 4'd3;
@(posedge clk_i);
shared_exps0 = 8'd143;
shared_exps1 = 8'd143;
a_mant0 = 8'd211; a_mant1 = 8'd145; a_mant2 = 8'd75; a_mant3 = 8'd147;
b_mant0 = 8'd198; b_mant1 = 8'd158; b_mant2 = 8'd171; b_mant3 = 8'd18;
a_exp0 = 10'd792; a_exp1 = 10'd478; a_exp2 = 10'd287; a_exp3 = 10'd962;
b_exp0 = 10'd372; b_exp1 = 10'd562; b_exp2 = 10'd477; b_exp3 = 10'd331;
a_sign0 = 4'd12; a_sign1 = 4'd10; a_sign2 = 4'd1; a_sign3 = 4'd1;
b_sign0 = 4'd9; b_sign1 = 4'd2; b_sign2 = 4'd13; b_sign3 = 4'd2;
@(posedge clk_i);
a_mant0 = 8'd209; a_mant1 = 8'd109; a_mant2 = 8'd155; a_mant3 = 8'd243;
b_mant0 = 8'd51; b_mant1 = 8'd71; b_mant2 = 8'd108; b_mant3 = 8'd93;
a_exp0 = 10'd665; a_exp1 = 10'd949; a_exp2 = 10'd353; a_exp3 = 10'd488;
b_exp0 = 10'd640; b_exp1 = 10'd494; b_exp2 = 10'd329; b_exp3 = 10'd817;
a_sign0 = 4'd1; a_sign1 = 4'd12; a_sign2 = 4'd14; a_sign3 = 4'd12;
b_sign0 = 4'd7; b_sign1 = 4'd13; b_sign2 = 4'd1; b_sign3 = 4'd5;
@(posedge clk_i);
a_mant0 = 8'd232; a_mant1 = 8'd176; a_mant2 = 8'd80; a_mant3 = 8'd54;
b_mant0 = 8'd123; b_mant1 = 8'd121; b_mant2 = 8'd130; b_mant3 = 8'd138;
a_exp0 = 10'd445; a_exp1 = 10'd203; a_exp2 = 10'd863; a_exp3 = 10'd51;
b_exp0 = 10'd482; b_exp1 = 10'd1020; b_exp2 = 10'd592; b_exp3 = 10'd64;
a_sign0 = 4'd11; a_sign1 = 4'd14; a_sign2 = 4'd1; a_sign3 = 4'd5;
b_sign0 = 4'd3; b_sign1 = 4'd4; b_sign2 = 4'd11; b_sign3 = 4'd4;
@(posedge clk_i);
a_mant0 = 8'd118; a_mant1 = 8'd27; a_mant2 = 8'd187; a_mant3 = 8'd138;
b_mant0 = 8'd123; b_mant1 = 8'd75; b_mant2 = 8'd84; b_mant3 = 8'd239;
a_exp0 = 10'd601; a_exp1 = 10'd90; a_exp2 = 10'd653; a_exp3 = 10'd458;
b_exp0 = 10'd691; b_exp1 = 10'd536; b_exp2 = 10'd198; b_exp3 = 10'd731;
a_sign0 = 4'd13; a_sign1 = 4'd0; a_sign2 = 4'd5; a_sign3 = 4'd4;
b_sign0 = 4'd5; b_sign1 = 4'd3; b_sign2 = 4'd15; b_sign3 = 4'd3;
@(posedge clk_i);
a_mant0 = 8'd105; a_mant1 = 8'd74; a_mant2 = 8'd78; a_mant3 = 8'd236;
b_mant0 = 8'd106; b_mant1 = 8'd136; b_mant2 = 8'd48; b_mant3 = 8'd244;
a_exp0 = 10'd197; a_exp1 = 10'd481; a_exp2 = 10'd495; a_exp3 = 10'd223;
b_exp0 = 10'd1019; b_exp1 = 10'd253; b_exp2 = 10'd527; b_exp3 = 10'd600;
a_sign0 = 4'd0; a_sign1 = 4'd1; a_sign2 = 4'd6; a_sign3 = 4'd10;
b_sign0 = 4'd1; b_sign1 = 4'd4; b_sign2 = 4'd8; b_sign3 = 4'd6;
@(posedge clk_i);
a_mant0 = 8'd238; a_mant1 = 8'd174; a_mant2 = 8'd65; a_mant3 = 8'd223;
b_mant0 = 8'd241; b_mant1 = 8'd122; b_mant2 = 8'd181; b_mant3 = 8'd3;
a_exp0 = 10'd81; a_exp1 = 10'd176; a_exp2 = 10'd780; a_exp3 = 10'd462;
b_exp0 = 10'd427; b_exp1 = 10'd857; b_exp2 = 10'd171; b_exp3 = 10'd140;
a_sign0 = 4'd1; a_sign1 = 4'd10; a_sign2 = 4'd7; a_sign3 = 4'd11;
b_sign0 = 4'd8; b_sign1 = 4'd16; b_sign2 = 4'd13; b_sign3 = 4'd10;
@(posedge clk_i);
a_mant0 = 8'd249; a_mant1 = 8'd158; a_mant2 = 8'd32; a_mant3 = 8'd134;
b_mant0 = 8'd159; b_mant1 = 8'd80; b_mant2 = 8'd13; b_mant3 = 8'd148;
a_exp0 = 10'd917; a_exp1 = 10'd267; a_exp2 = 10'd482; a_exp3 = 10'd183;
b_exp0 = 10'd435; b_exp1 = 10'd324; b_exp2 = 10'd552; b_exp3 = 10'd355;
a_sign0 = 4'd16; a_sign1 = 4'd7; a_sign2 = 4'd2; a_sign3 = 4'd6;
b_sign0 = 4'd0; b_sign1 = 4'd10; b_sign2 = 4'd1; b_sign3 = 4'd8;
@(posedge clk_i);
a_mant0 = 8'd193; a_mant1 = 8'd25; a_mant2 = 8'd19; a_mant3 = 8'd32;
b_mant0 = 8'd184; b_mant1 = 8'd30; b_mant2 = 8'd197; b_mant3 = 8'd216;
a_exp0 = 10'd680; a_exp1 = 10'd614; a_exp2 = 10'd75; a_exp3 = 10'd72;
b_exp0 = 10'd462; b_exp1 = 10'd479; b_exp2 = 10'd823; b_exp3 = 10'd149;
a_sign0 = 4'd15; a_sign1 = 4'd13; a_sign2 = 4'd3; a_sign3 = 4'd8;
b_sign0 = 4'd6; b_sign1 = 4'd0; b_sign2 = 4'd11; b_sign3 = 4'd16;
@(posedge clk_i);
shared_exps0 = 8'd124;
shared_exps1 = 8'd131;
a_mant0 = 8'd233; a_mant1 = 8'd159; a_mant2 = 8'd13; a_mant3 = 8'd195;
b_mant0 = 8'd82; b_mant1 = 8'd160; b_mant2 = 8'd252; b_mant3 = 8'd26;
a_exp0 = 10'd969; a_exp1 = 10'd679; a_exp2 = 10'd219; a_exp3 = 10'd442;
b_exp0 = 10'd492; b_exp1 = 10'd635; b_exp2 = 10'd893; b_exp3 = 10'd937;
a_sign0 = 4'd2; a_sign1 = 4'd7; a_sign2 = 4'd8; a_sign3 = 4'd11;
b_sign0 = 4'd1; b_sign1 = 4'd1; b_sign2 = 4'd10; b_sign3 = 4'd3;
@(posedge clk_i);
a_mant0 = 8'd9; a_mant1 = 8'd250; a_mant2 = 8'd98; a_mant3 = 8'd70;
b_mant0 = 8'd70; b_mant1 = 8'd150; b_mant2 = 8'd43; b_mant3 = 8'd222;
a_exp0 = 10'd355; a_exp1 = 10'd261; a_exp2 = 10'd56; a_exp3 = 10'd355;
b_exp0 = 10'd696; b_exp1 = 10'd821; b_exp2 = 10'd284; b_exp3 = 10'd996;
a_sign0 = 4'd13; a_sign1 = 4'd14; a_sign2 = 4'd10; a_sign3 = 4'd16;
b_sign0 = 4'd13; b_sign1 = 4'd0; b_sign2 = 4'd16; b_sign3 = 4'd13;
@(posedge clk_i);
a_mant0 = 8'd176; a_mant1 = 8'd107; a_mant2 = 8'd64; a_mant3 = 8'd62;
b_mant0 = 8'd169; b_mant1 = 8'd7; b_mant2 = 8'd6; b_mant3 = 8'd241;
a_exp0 = 10'd270; a_exp1 = 10'd544; a_exp2 = 10'd413; a_exp3 = 10'd752;
b_exp0 = 10'd755; b_exp1 = 10'd8; b_exp2 = 10'd546; b_exp3 = 10'd265;
a_sign0 = 4'd12; a_sign1 = 4'd1; a_sign2 = 4'd9; a_sign3 = 4'd16;
b_sign0 = 4'd5; b_sign1 = 4'd11; b_sign2 = 4'd4; b_sign3 = 4'd12;
@(posedge clk_i);
a_mant0 = 8'd10; a_mant1 = 8'd148; a_mant2 = 8'd197; a_mant3 = 8'd55;
b_mant0 = 8'd162; b_mant1 = 8'd63; b_mant2 = 8'd102; b_mant3 = 8'd166;
a_exp0 = 10'd886; a_exp1 = 10'd158; a_exp2 = 10'd707; a_exp3 = 10'd91;
b_exp0 = 10'd992; b_exp1 = 10'd563; b_exp2 = 10'd16; b_exp3 = 10'd8;
a_sign0 = 4'd14; a_sign1 = 4'd1; a_sign2 = 4'd16; a_sign3 = 4'd8;
b_sign0 = 4'd7; b_sign1 = 4'd4; b_sign2 = 4'd1; b_sign3 = 4'd9;
@(posedge clk_i);
a_mant0 = 8'd215; a_mant1 = 8'd173; a_mant2 = 8'd24; a_mant3 = 8'd78;
b_mant0 = 8'd22; b_mant1 = 8'd126; b_mant2 = 8'd134; b_mant3 = 8'd215;
a_exp0 = 10'd447; a_exp1 = 10'd569; a_exp2 = 10'd209; a_exp3 = 10'd153;
b_exp0 = 10'd650; b_exp1 = 10'd796; b_exp2 = 10'd495; b_exp3 = 10'd358;
a_sign0 = 4'd8; a_sign1 = 4'd4; a_sign2 = 4'd15; a_sign3 = 4'd13;
b_sign0 = 4'd9; b_sign1 = 4'd16; b_sign2 = 4'd9; b_sign3 = 4'd1;
@(posedge clk_i);
a_mant0 = 8'd32; a_mant1 = 8'd250; a_mant2 = 8'd138; a_mant3 = 8'd199;
b_mant0 = 8'd63; b_mant1 = 8'd237; b_mant2 = 8'd222; b_mant3 = 8'd195;
a_exp0 = 10'd759; a_exp1 = 10'd672; a_exp2 = 10'd550; a_exp3 = 10'd585;
b_exp0 = 10'd531; b_exp1 = 10'd1006; b_exp2 = 10'd647; b_exp3 = 10'd237;
a_sign0 = 4'd1; a_sign1 = 4'd4; a_sign2 = 4'd14; a_sign3 = 4'd12;
b_sign0 = 4'd7; b_sign1 = 4'd7; b_sign2 = 4'd11; b_sign3 = 4'd4;
@(posedge clk_i);
a_mant0 = 8'd212; a_mant1 = 8'd126; a_mant2 = 8'd96; a_mant3 = 8'd207;
b_mant0 = 8'd151; b_mant1 = 8'd78; b_mant2 = 8'd35; b_mant3 = 8'd120;
a_exp0 = 10'd75; a_exp1 = 10'd367; a_exp2 = 10'd182; a_exp3 = 10'd230;
b_exp0 = 10'd950; b_exp1 = 10'd622; b_exp2 = 10'd548; b_exp3 = 10'd225;
a_sign0 = 4'd6; a_sign1 = 4'd14; a_sign2 = 4'd2; a_sign3 = 4'd8;
b_sign0 = 4'd0; b_sign1 = 4'd12; b_sign2 = 4'd16; b_sign3 = 4'd8;
@(posedge clk_i);
a_mant0 = 8'd225; a_mant1 = 8'd180; a_mant2 = 8'd199; a_mant3 = 8'd230;
b_mant0 = 8'd69; b_mant1 = 8'd55; b_mant2 = 8'd116; b_mant3 = 8'd162;
a_exp0 = 10'd994; a_exp1 = 10'd493; a_exp2 = 10'd94; a_exp3 = 10'd173;
b_exp0 = 10'd58; b_exp1 = 10'd629; b_exp2 = 10'd286; b_exp3 = 10'd222;
a_sign0 = 4'd2; a_sign1 = 4'd10; a_sign2 = 4'd15; a_sign3 = 4'd11;
b_sign0 = 4'd14; b_sign1 = 4'd11; b_sign2 = 4'd1; b_sign3 = 4'd0;
@(posedge clk_i);
shared_exps0 = 8'd150;
shared_exps1 = 8'd107;
rstn = 0;
@(posedge clk_i);
rstn = 1;
a_mant0 = 8'd218; a_mant1 = 8'd136; a_mant2 = 8'd161; a_mant3 = 8'd3;
b_mant0 = 8'd243; b_mant1 = 8'd153; b_mant2 = 8'd219; b_mant3 = 8'd14;
a_exp0 = 10'd495; a_exp1 = 10'd512; a_exp2 = 10'd206; a_exp3 = 10'd348;
b_exp0 = 10'd554; b_exp1 = 10'd94; b_exp2 = 10'd571; b_exp3 = 10'd755;
a_sign0 = 4'd13; a_sign1 = 4'd1; a_sign2 = 4'd3; a_sign3 = 4'd5;
b_sign0 = 4'd1; b_sign1 = 4'd4; b_sign2 = 4'd3; b_sign3 = 4'd8;
@(posedge clk_i);
a_mant0 = 8'd209; a_mant1 = 8'd32; a_mant2 = 8'd240; a_mant3 = 8'd181;
b_mant0 = 8'd5; b_mant1 = 8'd223; b_mant2 = 8'd138; b_mant3 = 8'd43;
a_exp0 = 10'd54; a_exp1 = 10'd349; a_exp2 = 10'd82; a_exp3 = 10'd252;
b_exp0 = 10'd634; b_exp1 = 10'd841; b_exp2 = 10'd895; b_exp3 = 10'd782;
a_sign0 = 4'd2; a_sign1 = 4'd0; a_sign2 = 4'd4; a_sign3 = 4'd9;
b_sign0 = 4'd2; b_sign1 = 4'd15; b_sign2 = 4'd9; b_sign3 = 4'd7;
@(posedge clk_i);
a_mant0 = 8'd124; a_mant1 = 8'd113; a_mant2 = 8'd60; a_mant3 = 8'd91;
b_mant0 = 8'd18; b_mant1 = 8'd110; b_mant2 = 8'd107; b_mant3 = 8'd194;
a_exp0 = 10'd868; a_exp1 = 10'd591; a_exp2 = 10'd523; a_exp3 = 10'd143;
b_exp0 = 10'd228; b_exp1 = 10'd962; b_exp2 = 10'd796; b_exp3 = 10'd52;
a_sign0 = 4'd11; a_sign1 = 4'd12; a_sign2 = 4'd0; a_sign3 = 4'd16;
b_sign0 = 4'd12; b_sign1 = 4'd5; b_sign2 = 4'd3; b_sign3 = 4'd3;
@(posedge clk_i);
a_mant0 = 8'd45; a_mant1 = 8'd73; a_mant2 = 8'd145; a_mant3 = 8'd201;
b_mant0 = 8'd97; b_mant1 = 8'd8; b_mant2 = 8'd129; b_mant3 = 8'd1;
a_exp0 = 10'd770; a_exp1 = 10'd355; a_exp2 = 10'd792; a_exp3 = 10'd414;
b_exp0 = 10'd38; b_exp1 = 10'd134; b_exp2 = 10'd343; b_exp3 = 10'd349;
a_sign0 = 4'd13; a_sign1 = 4'd6; a_sign2 = 4'd8; a_sign3 = 4'd9;
b_sign0 = 4'd11; b_sign1 = 4'd9; b_sign2 = 4'd1; b_sign3 = 4'd12;
@(posedge clk_i);
a_mant0 = 8'd197; a_mant1 = 8'd237; a_mant2 = 8'd168; a_mant3 = 8'd12;
b_mant0 = 8'd36; b_mant1 = 8'd49; b_mant2 = 8'd166; b_mant3 = 8'd166;
a_exp0 = 10'd267; a_exp1 = 10'd169; a_exp2 = 10'd706; a_exp3 = 10'd930;
b_exp0 = 10'd297; b_exp1 = 10'd736; b_exp2 = 10'd971; b_exp3 = 10'd187;
a_sign0 = 4'd1; a_sign1 = 4'd7; a_sign2 = 4'd16; a_sign3 = 4'd10;
b_sign0 = 4'd13; b_sign1 = 4'd7; b_sign2 = 4'd10; b_sign3 = 4'd12;
@(posedge clk_i);
a_mant0 = 8'd141; a_mant1 = 8'd131; a_mant2 = 8'd233; a_mant3 = 8'd187;
b_mant0 = 8'd36; b_mant1 = 8'd44; b_mant2 = 8'd150; b_mant3 = 8'd99;
a_exp0 = 10'd209; a_exp1 = 10'd683; a_exp2 = 10'd87; a_exp3 = 10'd9;
b_exp0 = 10'd96; b_exp1 = 10'd572; b_exp2 = 10'd113; b_exp3 = 10'd904;
a_sign0 = 4'd15; a_sign1 = 4'd5; a_sign2 = 4'd9; a_sign3 = 4'd7;
b_sign0 = 4'd6; b_sign1 = 4'd16; b_sign2 = 4'd13; b_sign3 = 4'd2;
@(posedge clk_i);
a_mant0 = 8'd172; a_mant1 = 8'd57; a_mant2 = 8'd123; a_mant3 = 8'd253;
b_mant0 = 8'd224; b_mant1 = 8'd6; b_mant2 = 8'd74; b_mant3 = 8'd181;
a_exp0 = 10'd890; a_exp1 = 10'd672; a_exp2 = 10'd909; a_exp3 = 10'd267;
b_exp0 = 10'd982; b_exp1 = 10'd411; b_exp2 = 10'd902; b_exp3 = 10'd613;
a_sign0 = 4'd0; a_sign1 = 4'd6; a_sign2 = 4'd0; a_sign3 = 4'd10;
b_sign0 = 4'd15; b_sign1 = 4'd9; b_sign2 = 4'd6; b_sign3 = 4'd14;
@(posedge clk_i);
shared_exps0 = 8'd125;
shared_exps1 = 8'd129;
a_mant0 = 8'd117; a_mant1 = 8'd122; a_mant2 = 8'd25; a_mant3 = 8'd250;
b_mant0 = 8'd33; b_mant1 = 8'd53; b_mant2 = 8'd129; b_mant3 = 8'd47;
a_exp0 = 10'd92; a_exp1 = 10'd948; a_exp2 = 10'd477; a_exp3 = 10'd441;
b_exp0 = 10'd648; b_exp1 = 10'd818; b_exp2 = 10'd455; b_exp3 = 10'd122;
a_sign0 = 4'd15; a_sign1 = 4'd13; a_sign2 = 4'd10; a_sign3 = 4'd9;
b_sign0 = 4'd11; b_sign1 = 4'd10; b_sign2 = 4'd16; b_sign3 = 4'd11;
@(posedge clk_i);
a_mant0 = 8'd106; a_mant1 = 8'd238; a_mant2 = 8'd91; a_mant3 = 8'd177;
b_mant0 = 8'd242; b_mant1 = 8'd103; b_mant2 = 8'd169; b_mant3 = 8'd215;
a_exp0 = 10'd274; a_exp1 = 10'd342; a_exp2 = 10'd888; a_exp3 = 10'd287;
b_exp0 = 10'd325; b_exp1 = 10'd265; b_exp2 = 10'd524; b_exp3 = 10'd768;
a_sign0 = 4'd5; a_sign1 = 4'd11; a_sign2 = 4'd0; a_sign3 = 4'd1;
b_sign0 = 4'd1; b_sign1 = 4'd5; b_sign2 = 4'd3; b_sign3 = 4'd8;
@(posedge clk_i);
a_mant0 = 8'd145; a_mant1 = 8'd115; a_mant2 = 8'd102; a_mant3 = 8'd36;
b_mant0 = 8'd250; b_mant1 = 8'd36; b_mant2 = 8'd172; b_mant3 = 8'd95;
a_exp0 = 10'd908; a_exp1 = 10'd647; a_exp2 = 10'd632; a_exp3 = 10'd211;
b_exp0 = 10'd496; b_exp1 = 10'd625; b_exp2 = 10'd700; b_exp3 = 10'd238;
a_sign0 = 4'd11; a_sign1 = 4'd6; a_sign2 = 4'd7; a_sign3 = 4'd6;
b_sign0 = 4'd11; b_sign1 = 4'd14; b_sign2 = 4'd6; b_sign3 = 4'd13;
@(posedge clk_i);
a_mant0 = 8'd215; a_mant1 = 8'd60; a_mant2 = 8'd10; a_mant3 = 8'd193;
b_mant0 = 8'd241; b_mant1 = 8'd240; b_mant2 = 8'd84; b_mant3 = 8'd172;
a_exp0 = 10'd669; a_exp1 = 10'd787; a_exp2 = 10'd366; a_exp3 = 10'd708;
b_exp0 = 10'd96; b_exp1 = 10'd661; b_exp2 = 10'd38; b_exp3 = 10'd535;
a_sign0 = 4'd7; a_sign1 = 4'd15; a_sign2 = 4'd5; a_sign3 = 4'd11;
b_sign0 = 4'd7; b_sign1 = 4'd7; b_sign2 = 4'd16; b_sign3 = 4'd3;
@(posedge clk_i);
a_mant0 = 8'd239; a_mant1 = 8'd50; a_mant2 = 8'd55; a_mant3 = 8'd14;
b_mant0 = 8'd68; b_mant1 = 8'd81; b_mant2 = 8'd55; b_mant3 = 8'd124;
a_exp0 = 10'd953; a_exp1 = 10'd940; a_exp2 = 10'd107; a_exp3 = 10'd179;
b_exp0 = 10'd161; b_exp1 = 10'd635; b_exp2 = 10'd826; b_exp3 = 10'd849;
a_sign0 = 4'd1; a_sign1 = 4'd14; a_sign2 = 4'd12; a_sign3 = 4'd12;
b_sign0 = 4'd3; b_sign1 = 4'd10; b_sign2 = 4'd0; b_sign3 = 4'd9;
@(posedge clk_i);
a_mant0 = 8'd94; a_mant1 = 8'd196; a_mant2 = 8'd190; a_mant3 = 8'd45;
b_mant0 = 8'd240; b_mant1 = 8'd20; b_mant2 = 8'd169; b_mant3 = 8'd115;
a_exp0 = 10'd359; a_exp1 = 10'd428; a_exp2 = 10'd472; a_exp3 = 10'd859;
b_exp0 = 10'd475; b_exp1 = 10'd678; b_exp2 = 10'd812; b_exp3 = 10'd60;
a_sign0 = 4'd16; a_sign1 = 4'd13; a_sign2 = 4'd5; a_sign3 = 4'd16;
b_sign0 = 4'd5; b_sign1 = 4'd5; b_sign2 = 4'd5; b_sign3 = 4'd1;
@(posedge clk_i);
a_mant0 = 8'd118; a_mant1 = 8'd162; a_mant2 = 8'd245; a_mant3 = 8'd223;
b_mant0 = 8'd176; b_mant1 = 8'd198; b_mant2 = 8'd97; b_mant3 = 8'd133;
a_exp0 = 10'd386; a_exp1 = 10'd486; a_exp2 = 10'd573; a_exp3 = 10'd1006;
b_exp0 = 10'd750; b_exp1 = 10'd618; b_exp2 = 10'd53; b_exp3 = 10'd957;
a_sign0 = 4'd3; a_sign1 = 4'd9; a_sign2 = 4'd3; a_sign3 = 4'd10;
b_sign0 = 4'd8; b_sign1 = 4'd8; b_sign2 = 4'd12; b_sign3 = 4'd1;
@(posedge clk_i);
a_mant0 = 8'd96; a_mant1 = 8'd131; a_mant2 = 8'd148; a_mant3 = 8'd125;
b_mant0 = 8'd56; b_mant1 = 8'd136; b_mant2 = 8'd240; b_mant3 = 8'd145;
a_exp0 = 10'd789; a_exp1 = 10'd760; a_exp2 = 10'd888; a_exp3 = 10'd414;
b_exp0 = 10'd76; b_exp1 = 10'd435; b_exp2 = 10'd782; b_exp3 = 10'd219;
a_sign0 = 4'd5; a_sign1 = 4'd13; a_sign2 = 4'd9; a_sign3 = 4'd9;
b_sign0 = 4'd8; b_sign1 = 4'd10; b_sign2 = 4'd16; b_sign3 = 4'd3;
@(posedge clk_i);
shared_exps0 = 8'd131;
shared_exps1 = 8'd116;
a_mant0 = 8'd215; a_mant1 = 8'd58; a_mant2 = 8'd175; a_mant3 = 8'd26;
b_mant0 = 8'd39; b_mant1 = 8'd202; b_mant2 = 8'd3; b_mant3 = 8'd21;
a_exp0 = 10'd110; a_exp1 = 10'd609; a_exp2 = 10'd822; a_exp3 = 10'd345;
b_exp0 = 10'd303; b_exp1 = 10'd522; b_exp2 = 10'd147; b_exp3 = 10'd494;
a_sign0 = 4'd3; a_sign1 = 4'd2; a_sign2 = 4'd16; a_sign3 = 4'd9;
b_sign0 = 4'd14; b_sign1 = 4'd12; b_sign2 = 4'd9; b_sign3 = 4'd3;
@(posedge clk_i);
a_mant0 = 8'd130; a_mant1 = 8'd20; a_mant2 = 8'd209; a_mant3 = 8'd3;
b_mant0 = 8'd31; b_mant1 = 8'd178; b_mant2 = 8'd93; b_mant3 = 8'd43;
a_exp0 = 10'd655; a_exp1 = 10'd397; a_exp2 = 10'd495; a_exp3 = 10'd665;
b_exp0 = 10'd403; b_exp1 = 10'd97; b_exp2 = 10'd846; b_exp3 = 10'd67;
a_sign0 = 4'd8; a_sign1 = 4'd5; a_sign2 = 4'd2; a_sign3 = 4'd8;
b_sign0 = 4'd2; b_sign1 = 4'd7; b_sign2 = 4'd4; b_sign3 = 4'd7;
@(posedge clk_i);
a_mant0 = 8'd108; a_mant1 = 8'd181; a_mant2 = 8'd2; a_mant3 = 8'd56;
b_mant0 = 8'd45; b_mant1 = 8'd60; b_mant2 = 8'd214; b_mant3 = 8'd234;
a_exp0 = 10'd429; a_exp1 = 10'd402; a_exp2 = 10'd898; a_exp3 = 10'd600;
b_exp0 = 10'd880; b_exp1 = 10'd644; b_exp2 = 10'd687; b_exp3 = 10'd742;
a_sign0 = 4'd16; a_sign1 = 4'd1; a_sign2 = 4'd12; a_sign3 = 4'd14;
b_sign0 = 4'd16; b_sign1 = 4'd11; b_sign2 = 4'd4; b_sign3 = 4'd11;
@(posedge clk_i);
a_mant0 = 8'd172; a_mant1 = 8'd94; a_mant2 = 8'd61; a_mant3 = 8'd72;
b_mant0 = 8'd82; b_mant1 = 8'd203; b_mant2 = 8'd220; b_mant3 = 8'd148;
a_exp0 = 10'd365; a_exp1 = 10'd708; a_exp2 = 10'd206; a_exp3 = 10'd629;
b_exp0 = 10'd982; b_exp1 = 10'd259; b_exp2 = 10'd11; b_exp3 = 10'd281;
a_sign0 = 4'd3; a_sign1 = 4'd11; a_sign2 = 4'd0; a_sign3 = 4'd6;
b_sign0 = 4'd16; b_sign1 = 4'd2; b_sign2 = 4'd12; b_sign3 = 4'd15;
@(posedge clk_i);
a_mant0 = 8'd92; a_mant1 = 8'd231; a_mant2 = 8'd92; a_mant3 = 8'd37;
b_mant0 = 8'd172; b_mant1 = 8'd16; b_mant2 = 8'd81; b_mant3 = 8'd198;
a_exp0 = 10'd678; a_exp1 = 10'd71; a_exp2 = 10'd326; a_exp3 = 10'd652;
b_exp0 = 10'd732; b_exp1 = 10'd214; b_exp2 = 10'd338; b_exp3 = 10'd555;
a_sign0 = 4'd4; a_sign1 = 4'd3; a_sign2 = 4'd1; a_sign3 = 4'd1;
b_sign0 = 4'd16; b_sign1 = 4'd1; b_sign2 = 4'd15; b_sign3 = 4'd4;
@(posedge clk_i);
a_mant0 = 8'd153; a_mant1 = 8'd175; a_mant2 = 8'd78; a_mant3 = 8'd196;
b_mant0 = 8'd37; b_mant1 = 8'd236; b_mant2 = 8'd173; b_mant3 = 8'd21;
a_exp0 = 10'd956; a_exp1 = 10'd674; a_exp2 = 10'd197; a_exp3 = 10'd276;
b_exp0 = 10'd397; b_exp1 = 10'd575; b_exp2 = 10'd736; b_exp3 = 10'd149;
a_sign0 = 4'd6; a_sign1 = 4'd16; a_sign2 = 4'd14; a_sign3 = 4'd7;
b_sign0 = 4'd4; b_sign1 = 4'd13; b_sign2 = 4'd1; b_sign3 = 4'd4;
@(posedge clk_i);
a_mant0 = 8'd110; a_mant1 = 8'd224; a_mant2 = 8'd222; a_mant3 = 8'd250;
b_mant0 = 8'd134; b_mant1 = 8'd62; b_mant2 = 8'd190; b_mant3 = 8'd152;
a_exp0 = 10'd135; a_exp1 = 10'd775; a_exp2 = 10'd592; a_exp3 = 10'd450;
b_exp0 = 10'd263; b_exp1 = 10'd223; b_exp2 = 10'd616; b_exp3 = 10'd728;
a_sign0 = 4'd12; a_sign1 = 4'd15; a_sign2 = 4'd14; a_sign3 = 4'd14;
b_sign0 = 4'd3; b_sign1 = 4'd14; b_sign2 = 4'd4; b_sign3 = 4'd3;
@(posedge clk_i);
a_mant0 = 8'd145; a_mant1 = 8'd35; a_mant2 = 8'd219; a_mant3 = 8'd10;
b_mant0 = 8'd85; b_mant1 = 8'd196; b_mant2 = 8'd255; b_mant3 = 8'd252;
a_exp0 = 10'd350; a_exp1 = 10'd690; a_exp2 = 10'd524; a_exp3 = 10'd431;
b_exp0 = 10'd571; b_exp1 = 10'd145; b_exp2 = 10'd46; b_exp3 = 10'd19;
a_sign0 = 4'd2; a_sign1 = 4'd12; a_sign2 = 4'd4; a_sign3 = 4'd9;
b_sign0 = 4'd11; b_sign1 = 4'd1; b_sign2 = 4'd4; b_sign3 = 4'd0;
@(posedge clk_i);
shared_exps0 = 8'd131;
shared_exps1 = 8'd121;
a_mant0 = 8'd250; a_mant1 = 8'd0; a_mant2 = 8'd89; a_mant3 = 8'd106;
b_mant0 = 8'd91; b_mant1 = 8'd154; b_mant2 = 8'd170; b_mant3 = 8'd217;
a_exp0 = 10'd614; a_exp1 = 10'd315; a_exp2 = 10'd131; a_exp3 = 10'd25;
b_exp0 = 10'd903; b_exp1 = 10'd859; b_exp2 = 10'd410; b_exp3 = 10'd517;
a_sign0 = 4'd1; a_sign1 = 4'd9; a_sign2 = 4'd0; a_sign3 = 4'd0;
b_sign0 = 4'd15; b_sign1 = 4'd12; b_sign2 = 4'd7; b_sign3 = 4'd6;
@(posedge clk_i);
a_mant0 = 8'd108; a_mant1 = 8'd205; a_mant2 = 8'd47; a_mant3 = 8'd93;
b_mant0 = 8'd162; b_mant1 = 8'd248; b_mant2 = 8'd149; b_mant3 = 8'd183;
a_exp0 = 10'd962; a_exp1 = 10'd889; a_exp2 = 10'd985; a_exp3 = 10'd93;
b_exp0 = 10'd556; b_exp1 = 10'd655; b_exp2 = 10'd981; b_exp3 = 10'd530;
a_sign0 = 4'd8; a_sign1 = 4'd13; a_sign2 = 4'd11; a_sign3 = 4'd1;
b_sign0 = 4'd15; b_sign1 = 4'd15; b_sign2 = 4'd16; b_sign3 = 4'd3;
@(posedge clk_i);
a_mant0 = 8'd244; a_mant1 = 8'd207; a_mant2 = 8'd227; a_mant3 = 8'd162;
b_mant0 = 8'd183; b_mant1 = 8'd228; b_mant2 = 8'd199; b_mant3 = 8'd41;
a_exp0 = 10'd732; a_exp1 = 10'd359; a_exp2 = 10'd932; a_exp3 = 10'd168;
b_exp0 = 10'd552; b_exp1 = 10'd273; b_exp2 = 10'd862; b_exp3 = 10'd993;
a_sign0 = 4'd6; a_sign1 = 4'd0; a_sign2 = 4'd9; a_sign3 = 4'd12;
b_sign0 = 4'd12; b_sign1 = 4'd5; b_sign2 = 4'd16; b_sign3 = 4'd3;
@(posedge clk_i);
a_mant0 = 8'd231; a_mant1 = 8'd52; a_mant2 = 8'd6; a_mant3 = 8'd50;
b_mant0 = 8'd246; b_mant1 = 8'd167; b_mant2 = 8'd178; b_mant3 = 8'd130;
a_exp0 = 10'd399; a_exp1 = 10'd864; a_exp2 = 10'd105; a_exp3 = 10'd438;
b_exp0 = 10'd198; b_exp1 = 10'd377; b_exp2 = 10'd210; b_exp3 = 10'd784;
a_sign0 = 4'd3; a_sign1 = 4'd6; a_sign2 = 4'd3; a_sign3 = 4'd12;
b_sign0 = 4'd4; b_sign1 = 4'd11; b_sign2 = 4'd4; b_sign3 = 4'd1;
@(posedge clk_i);
a_mant0 = 8'd170; a_mant1 = 8'd187; a_mant2 = 8'd186; a_mant3 = 8'd254;
b_mant0 = 8'd175; b_mant1 = 8'd26; b_mant2 = 8'd92; b_mant3 = 8'd238;
a_exp0 = 10'd102; a_exp1 = 10'd774; a_exp2 = 10'd991; a_exp3 = 10'd408;
b_exp0 = 10'd477; b_exp1 = 10'd735; b_exp2 = 10'd731; b_exp3 = 10'd178;
a_sign0 = 4'd5; a_sign1 = 4'd6; a_sign2 = 4'd11; a_sign3 = 4'd4;
b_sign0 = 4'd5; b_sign1 = 4'd13; b_sign2 = 4'd6; b_sign3 = 4'd2;
@(posedge clk_i);
a_mant0 = 8'd100; a_mant1 = 8'd38; a_mant2 = 8'd165; a_mant3 = 8'd156;
b_mant0 = 8'd41; b_mant1 = 8'd24; b_mant2 = 8'd114; b_mant3 = 8'd131;
a_exp0 = 10'd340; a_exp1 = 10'd806; a_exp2 = 10'd552; a_exp3 = 10'd108;
b_exp0 = 10'd118; b_exp1 = 10'd672; b_exp2 = 10'd776; b_exp3 = 10'd691;
a_sign0 = 4'd9; a_sign1 = 4'd16; a_sign2 = 4'd16; a_sign3 = 4'd6;
b_sign0 = 4'd14; b_sign1 = 4'd0; b_sign2 = 4'd14; b_sign3 = 4'd15;
@(posedge clk_i);
a_mant0 = 8'd178; a_mant1 = 8'd239; a_mant2 = 8'd202; a_mant3 = 8'd2;
b_mant0 = 8'd60; b_mant1 = 8'd23; b_mant2 = 8'd134; b_mant3 = 8'd123;
a_exp0 = 10'd701; a_exp1 = 10'd759; a_exp2 = 10'd899; a_exp3 = 10'd611;
b_exp0 = 10'd227; b_exp1 = 10'd714; b_exp2 = 10'd468; b_exp3 = 10'd149;
a_sign0 = 4'd11; a_sign1 = 4'd12; a_sign2 = 4'd14; a_sign3 = 4'd2;
b_sign0 = 4'd1; b_sign1 = 4'd10; b_sign2 = 4'd10; b_sign3 = 4'd13;
@(posedge clk_i);
a_mant0 = 8'd209; a_mant1 = 8'd23; a_mant2 = 8'd4; a_mant3 = 8'd101;
b_mant0 = 8'd184; b_mant1 = 8'd167; b_mant2 = 8'd209; b_mant3 = 8'd82;
a_exp0 = 10'd167; a_exp1 = 10'd228; a_exp2 = 10'd103; a_exp3 = 10'd541;
b_exp0 = 10'd575; b_exp1 = 10'd177; b_exp2 = 10'd746; b_exp3 = 10'd161;
a_sign0 = 4'd10; a_sign1 = 4'd6; a_sign2 = 4'd0; a_sign3 = 4'd3;
b_sign0 = 4'd6; b_sign1 = 4'd7; b_sign2 = 4'd7; b_sign3 = 4'd16;
@(posedge clk_i);
shared_exps0 = 8'd139;
shared_exps1 = 8'd149;
rstn = 0;
@(posedge clk_i);
rstn = 1;
a_mant0 = 8'd165; a_mant1 = 8'd72; a_mant2 = 8'd197; a_mant3 = 8'd111;
b_mant0 = 8'd151; b_mant1 = 8'd207; b_mant2 = 8'd58; b_mant3 = 8'd101;
a_exp0 = 10'd992; a_exp1 = 10'd742; a_exp2 = 10'd549; a_exp3 = 10'd354;
b_exp0 = 10'd784; b_exp1 = 10'd871; b_exp2 = 10'd528; b_exp3 = 10'd162;
a_sign0 = 4'd11; a_sign1 = 4'd9; a_sign2 = 4'd15; a_sign3 = 4'd4;
b_sign0 = 4'd7; b_sign1 = 4'd1; b_sign2 = 4'd9; b_sign3 = 4'd13;
@(posedge clk_i);
a_mant0 = 8'd189; a_mant1 = 8'd12; a_mant2 = 8'd61; a_mant3 = 8'd70;
b_mant0 = 8'd214; b_mant1 = 8'd245; b_mant2 = 8'd117; b_mant3 = 8'd78;
a_exp0 = 10'd467; a_exp1 = 10'd102; a_exp2 = 10'd501; a_exp3 = 10'd783;
b_exp0 = 10'd340; b_exp1 = 10'd918; b_exp2 = 10'd887; b_exp3 = 10'd610;
a_sign0 = 4'd3; a_sign1 = 4'd13; a_sign2 = 4'd7; a_sign3 = 4'd8;
b_sign0 = 4'd15; b_sign1 = 4'd4; b_sign2 = 4'd0; b_sign3 = 4'd9;
@(posedge clk_i);
a_mant0 = 8'd8; a_mant1 = 8'd110; a_mant2 = 8'd207; a_mant3 = 8'd78;
b_mant0 = 8'd155; b_mant1 = 8'd14; b_mant2 = 8'd7; b_mant3 = 8'd188;
a_exp0 = 10'd188; a_exp1 = 10'd323; a_exp2 = 10'd906; a_exp3 = 10'd683;
b_exp0 = 10'd510; b_exp1 = 10'd476; b_exp2 = 10'd386; b_exp3 = 10'd580;
a_sign0 = 4'd10; a_sign1 = 4'd15; a_sign2 = 4'd1; a_sign3 = 4'd3;
b_sign0 = 4'd7; b_sign1 = 4'd12; b_sign2 = 4'd0; b_sign3 = 4'd13;
@(posedge clk_i);
a_mant0 = 8'd207; a_mant1 = 8'd190; a_mant2 = 8'd36; a_mant3 = 8'd239;
b_mant0 = 8'd124; b_mant1 = 8'd120; b_mant2 = 8'd89; b_mant3 = 8'd59;
a_exp0 = 10'd705; a_exp1 = 10'd110; a_exp2 = 10'd171; a_exp3 = 10'd759;
b_exp0 = 10'd318; b_exp1 = 10'd810; b_exp2 = 10'd835; b_exp3 = 10'd16;
a_sign0 = 4'd16; a_sign1 = 4'd16; a_sign2 = 4'd2; a_sign3 = 4'd9;
b_sign0 = 4'd6; b_sign1 = 4'd15; b_sign2 = 4'd1; b_sign3 = 4'd7;
@(posedge clk_i);
a_mant0 = 8'd177; a_mant1 = 8'd130; a_mant2 = 8'd137; a_mant3 = 8'd176;
b_mant0 = 8'd55; b_mant1 = 8'd30; b_mant2 = 8'd34; b_mant3 = 8'd193;
a_exp0 = 10'd219; a_exp1 = 10'd205; a_exp2 = 10'd924; a_exp3 = 10'd76;
b_exp0 = 10'd678; b_exp1 = 10'd533; b_exp2 = 10'd271; b_exp3 = 10'd529;
a_sign0 = 4'd3; a_sign1 = 4'd16; a_sign2 = 4'd14; a_sign3 = 4'd2;
b_sign0 = 4'd2; b_sign1 = 4'd11; b_sign2 = 4'd7; b_sign3 = 4'd7;
@(posedge clk_i);
a_mant0 = 8'd218; a_mant1 = 8'd254; a_mant2 = 8'd27; a_mant3 = 8'd6;
b_mant0 = 8'd19; b_mant1 = 8'd87; b_mant2 = 8'd55; b_mant3 = 8'd54;
a_exp0 = 10'd644; a_exp1 = 10'd924; a_exp2 = 10'd811; a_exp3 = 10'd962;
b_exp0 = 10'd29; b_exp1 = 10'd744; b_exp2 = 10'd199; b_exp3 = 10'd214;
a_sign0 = 4'd13; a_sign1 = 4'd16; a_sign2 = 4'd10; a_sign3 = 4'd2;
b_sign0 = 4'd9; b_sign1 = 4'd15; b_sign2 = 4'd6; b_sign3 = 4'd5;
@(posedge clk_i);
a_mant0 = 8'd32; a_mant1 = 8'd148; a_mant2 = 8'd116; a_mant3 = 8'd19;
b_mant0 = 8'd104; b_mant1 = 8'd225; b_mant2 = 8'd237; b_mant3 = 8'd81;
a_exp0 = 10'd648; a_exp1 = 10'd851; a_exp2 = 10'd912; a_exp3 = 10'd4;
b_exp0 = 10'd61; b_exp1 = 10'd14; b_exp2 = 10'd208; b_exp3 = 10'd177;
a_sign0 = 4'd7; a_sign1 = 4'd9; a_sign2 = 4'd6; a_sign3 = 4'd3;
b_sign0 = 4'd9; b_sign1 = 4'd6; b_sign2 = 4'd1; b_sign3 = 4'd15;
@(posedge clk_i);
shared_exps0 = 8'd116;
shared_exps1 = 8'd126;
a_mant0 = 8'd140; a_mant1 = 8'd223; a_mant2 = 8'd79; a_mant3 = 8'd238;
b_mant0 = 8'd221; b_mant1 = 8'd128; b_mant2 = 8'd166; b_mant3 = 8'd141;
a_exp0 = 10'd40; a_exp1 = 10'd438; a_exp2 = 10'd950; a_exp3 = 10'd753;
b_exp0 = 10'd325; b_exp1 = 10'd410; b_exp2 = 10'd997; b_exp3 = 10'd790;
a_sign0 = 4'd15; a_sign1 = 4'd12; a_sign2 = 4'd6; a_sign3 = 4'd6;
b_sign0 = 4'd5; b_sign1 = 4'd3; b_sign2 = 4'd16; b_sign3 = 4'd1;
@(posedge clk_i);
a_mant0 = 8'd85; a_mant1 = 8'd76; a_mant2 = 8'd218; a_mant3 = 8'd157;
b_mant0 = 8'd66; b_mant1 = 8'd178; b_mant2 = 8'd118; b_mant3 = 8'd217;
a_exp0 = 10'd160; a_exp1 = 10'd76; a_exp2 = 10'd89; a_exp3 = 10'd408;
b_exp0 = 10'd369; b_exp1 = 10'd140; b_exp2 = 10'd852; b_exp3 = 10'd640;
a_sign0 = 4'd4; a_sign1 = 4'd3; a_sign2 = 4'd3; a_sign3 = 4'd15;
b_sign0 = 4'd6; b_sign1 = 4'd12; b_sign2 = 4'd4; b_sign3 = 4'd12;
@(posedge clk_i);
a_mant0 = 8'd239; a_mant1 = 8'd55; a_mant2 = 8'd37; a_mant3 = 8'd102;
b_mant0 = 8'd171; b_mant1 = 8'd1; b_mant2 = 8'd185; b_mant3 = 8'd247;
a_exp0 = 10'd607; a_exp1 = 10'd102; a_exp2 = 10'd836; a_exp3 = 10'd592;
b_exp0 = 10'd691; b_exp1 = 10'd658; b_exp2 = 10'd983; b_exp3 = 10'd177;
a_sign0 = 4'd4; a_sign1 = 4'd9; a_sign2 = 4'd9; a_sign3 = 4'd15;
b_sign0 = 4'd11; b_sign1 = 4'd9; b_sign2 = 4'd11; b_sign3 = 4'd7;
@(posedge clk_i);
a_mant0 = 8'd101; a_mant1 = 8'd40; a_mant2 = 8'd62; a_mant3 = 8'd142;
b_mant0 = 8'd107; b_mant1 = 8'd149; b_mant2 = 8'd54; b_mant3 = 8'd161;
a_exp0 = 10'd565; a_exp1 = 10'd712; a_exp2 = 10'd686; a_exp3 = 10'd148;
b_exp0 = 10'd415; b_exp1 = 10'd916; b_exp2 = 10'd402; b_exp3 = 10'd1005;
a_sign0 = 4'd16; a_sign1 = 4'd8; a_sign2 = 4'd3; a_sign3 = 4'd7;
b_sign0 = 4'd13; b_sign1 = 4'd11; b_sign2 = 4'd13; b_sign3 = 4'd16;
@(posedge clk_i);
a_mant0 = 8'd183; a_mant1 = 8'd63; a_mant2 = 8'd146; a_mant3 = 8'd138;
b_mant0 = 8'd194; b_mant1 = 8'd7; b_mant2 = 8'd5; b_mant3 = 8'd207;
a_exp0 = 10'd779; a_exp1 = 10'd11; a_exp2 = 10'd738; a_exp3 = 10'd668;
b_exp0 = 10'd423; b_exp1 = 10'd730; b_exp2 = 10'd247; b_exp3 = 10'd962;
a_sign0 = 4'd13; a_sign1 = 4'd3; a_sign2 = 4'd8; a_sign3 = 4'd11;
b_sign0 = 4'd0; b_sign1 = 4'd1; b_sign2 = 4'd9; b_sign3 = 4'd11;
@(posedge clk_i);
a_mant0 = 8'd218; a_mant1 = 8'd160; a_mant2 = 8'd112; a_mant3 = 8'd252;
b_mant0 = 8'd27; b_mant1 = 8'd187; b_mant2 = 8'd241; b_mant3 = 8'd26;
a_exp0 = 10'd360; a_exp1 = 10'd742; a_exp2 = 10'd975; a_exp3 = 10'd327;
b_exp0 = 10'd368; b_exp1 = 10'd570; b_exp2 = 10'd355; b_exp3 = 10'd259;
a_sign0 = 4'd2; a_sign1 = 4'd5; a_sign2 = 4'd16; a_sign3 = 4'd7;
b_sign0 = 4'd5; b_sign1 = 4'd3; b_sign2 = 4'd5; b_sign3 = 4'd14;
@(posedge clk_i);
a_mant0 = 8'd129; a_mant1 = 8'd136; a_mant2 = 8'd65; a_mant3 = 8'd201;
b_mant0 = 8'd174; b_mant1 = 8'd35; b_mant2 = 8'd74; b_mant3 = 8'd71;
a_exp0 = 10'd362; a_exp1 = 10'd116; a_exp2 = 10'd260; a_exp3 = 10'd41;
b_exp0 = 10'd97; b_exp1 = 10'd582; b_exp2 = 10'd195; b_exp3 = 10'd568;
a_sign0 = 4'd14; a_sign1 = 4'd14; a_sign2 = 4'd6; a_sign3 = 4'd11;
b_sign0 = 4'd12; b_sign1 = 4'd12; b_sign2 = 4'd1; b_sign3 = 4'd0;
@(posedge clk_i);
a_mant0 = 8'd169; a_mant1 = 8'd47; a_mant2 = 8'd153; a_mant3 = 8'd183;
b_mant0 = 8'd134; b_mant1 = 8'd153; b_mant2 = 8'd51; b_mant3 = 8'd123;
a_exp0 = 10'd552; a_exp1 = 10'd387; a_exp2 = 10'd709; a_exp3 = 10'd931;
b_exp0 = 10'd467; b_exp1 = 10'd593; b_exp2 = 10'd411; b_exp3 = 10'd605;
a_sign0 = 4'd11; a_sign1 = 4'd10; a_sign2 = 4'd11; a_sign3 = 4'd3;
b_sign0 = 4'd12; b_sign1 = 4'd1; b_sign2 = 4'd16; b_sign3 = 4'd7;
@(posedge clk_i);
shared_exps0 = 8'd111;
shared_exps1 = 8'd124;
a_mant0 = 8'd93; a_mant1 = 8'd220; a_mant2 = 8'd108; a_mant3 = 8'd4;
b_mant0 = 8'd12; b_mant1 = 8'd247; b_mant2 = 8'd28; b_mant3 = 8'd63;
a_exp0 = 10'd758; a_exp1 = 10'd91; a_exp2 = 10'd708; a_exp3 = 10'd918;
b_exp0 = 10'd610; b_exp1 = 10'd574; b_exp2 = 10'd122; b_exp3 = 10'd486;
a_sign0 = 4'd13; a_sign1 = 4'd6; a_sign2 = 4'd15; a_sign3 = 4'd3;
b_sign0 = 4'd3; b_sign1 = 4'd0; b_sign2 = 4'd9; b_sign3 = 4'd6;
@(posedge clk_i);
a_mant0 = 8'd65; a_mant1 = 8'd110; a_mant2 = 8'd181; a_mant3 = 8'd31;
b_mant0 = 8'd205; b_mant1 = 8'd195; b_mant2 = 8'd7; b_mant3 = 8'd113;
a_exp0 = 10'd290; a_exp1 = 10'd281; a_exp2 = 10'd732; a_exp3 = 10'd666;
b_exp0 = 10'd803; b_exp1 = 10'd514; b_exp2 = 10'd462; b_exp3 = 10'd765;
a_sign0 = 4'd8; a_sign1 = 4'd3; a_sign2 = 4'd11; a_sign3 = 4'd16;
b_sign0 = 4'd13; b_sign1 = 4'd11; b_sign2 = 4'd10; b_sign3 = 4'd14;
@(posedge clk_i);
a_mant0 = 8'd254; a_mant1 = 8'd42; a_mant2 = 8'd226; a_mant3 = 8'd244;
b_mant0 = 8'd160; b_mant1 = 8'd152; b_mant2 = 8'd226; b_mant3 = 8'd120;
a_exp0 = 10'd352; a_exp1 = 10'd579; a_exp2 = 10'd515; a_exp3 = 10'd701;
b_exp0 = 10'd220; b_exp1 = 10'd875; b_exp2 = 10'd366; b_exp3 = 10'd324;
a_sign0 = 4'd7; a_sign1 = 4'd5; a_sign2 = 4'd0; a_sign3 = 4'd12;
b_sign0 = 4'd1; b_sign1 = 4'd15; b_sign2 = 4'd13; b_sign3 = 4'd6;
@(posedge clk_i);
a_mant0 = 8'd65; a_mant1 = 8'd165; a_mant2 = 8'd166; a_mant3 = 8'd29;
b_mant0 = 8'd238; b_mant1 = 8'd58; b_mant2 = 8'd202; b_mant3 = 8'd5;
a_exp0 = 10'd697; a_exp1 = 10'd650; a_exp2 = 10'd967; a_exp3 = 10'd95;
b_exp0 = 10'd417; b_exp1 = 10'd282; b_exp2 = 10'd780; b_exp3 = 10'd219;
a_sign0 = 4'd16; a_sign1 = 4'd11; a_sign2 = 4'd5; a_sign3 = 4'd3;
b_sign0 = 4'd8; b_sign1 = 4'd1; b_sign2 = 4'd12; b_sign3 = 4'd12;
@(posedge clk_i);
a_mant0 = 8'd243; a_mant1 = 8'd139; a_mant2 = 8'd137; a_mant3 = 8'd6;
b_mant0 = 8'd222; b_mant1 = 8'd242; b_mant2 = 8'd101; b_mant3 = 8'd6;
a_exp0 = 10'd295; a_exp1 = 10'd690; a_exp2 = 10'd519; a_exp3 = 10'd601;
b_exp0 = 10'd488; b_exp1 = 10'd312; b_exp2 = 10'd96; b_exp3 = 10'd129;
a_sign0 = 4'd12; a_sign1 = 4'd16; a_sign2 = 4'd13; a_sign3 = 4'd9;
b_sign0 = 4'd0; b_sign1 = 4'd15; b_sign2 = 4'd4; b_sign3 = 4'd9;
@(posedge clk_i);
a_mant0 = 8'd54; a_mant1 = 8'd10; a_mant2 = 8'd171; a_mant3 = 8'd109;
b_mant0 = 8'd73; b_mant1 = 8'd216; b_mant2 = 8'd128; b_mant3 = 8'd137;
a_exp0 = 10'd290; a_exp1 = 10'd917; a_exp2 = 10'd166; a_exp3 = 10'd612;
b_exp0 = 10'd261; b_exp1 = 10'd897; b_exp2 = 10'd239; b_exp3 = 10'd811;
a_sign0 = 4'd11; a_sign1 = 4'd8; a_sign2 = 4'd6; a_sign3 = 4'd6;
b_sign0 = 4'd16; b_sign1 = 4'd15; b_sign2 = 4'd15; b_sign3 = 4'd15;
@(posedge clk_i);
a_mant0 = 8'd97; a_mant1 = 8'd248; a_mant2 = 8'd175; a_mant3 = 8'd111;
b_mant0 = 8'd206; b_mant1 = 8'd19; b_mant2 = 8'd38; b_mant3 = 8'd0;
a_exp0 = 10'd396; a_exp1 = 10'd570; a_exp2 = 10'd158; a_exp3 = 10'd975;
b_exp0 = 10'd303; b_exp1 = 10'd230; b_exp2 = 10'd870; b_exp3 = 10'd379;
a_sign0 = 4'd13; a_sign1 = 4'd4; a_sign2 = 4'd5; a_sign3 = 4'd0;
b_sign0 = 4'd16; b_sign1 = 4'd5; b_sign2 = 4'd1; b_sign3 = 4'd1;
@(posedge clk_i);
a_mant0 = 8'd75; a_mant1 = 8'd25; a_mant2 = 8'd54; a_mant3 = 8'd255;
b_mant0 = 8'd221; b_mant1 = 8'd35; b_mant2 = 8'd46; b_mant3 = 8'd109;
a_exp0 = 10'd515; a_exp1 = 10'd278; a_exp2 = 10'd856; a_exp3 = 10'd939;
b_exp0 = 10'd81; b_exp1 = 10'd134; b_exp2 = 10'd466; b_exp3 = 10'd355;
a_sign0 = 4'd4; a_sign1 = 4'd1; a_sign2 = 4'd12; a_sign3 = 4'd5;
b_sign0 = 4'd3; b_sign1 = 4'd10; b_sign2 = 4'd3; b_sign3 = 4'd9;
@(posedge clk_i);
shared_exps0 = 8'd118;
shared_exps1 = 8'd109;
a_mant0 = 8'd197; a_mant1 = 8'd237; a_mant2 = 8'd91; a_mant3 = 8'd12;
b_mant0 = 8'd208; b_mant1 = 8'd160; b_mant2 = 8'd164; b_mant3 = 8'd30;
a_exp0 = 10'd518; a_exp1 = 10'd62; a_exp2 = 10'd831; a_exp3 = 10'd165;
b_exp0 = 10'd405; b_exp1 = 10'd178; b_exp2 = 10'd54; b_exp3 = 10'd1020;
a_sign0 = 4'd1; a_sign1 = 4'd10; a_sign2 = 4'd14; a_sign3 = 4'd6;
b_sign0 = 4'd9; b_sign1 = 4'd2; b_sign2 = 4'd11; b_sign3 = 4'd13;
@(posedge clk_i);
a_mant0 = 8'd39; a_mant1 = 8'd196; a_mant2 = 8'd81; a_mant3 = 8'd76;
b_mant0 = 8'd38; b_mant1 = 8'd49; b_mant2 = 8'd247; b_mant3 = 8'd98;
a_exp0 = 10'd1003; a_exp1 = 10'd134; a_exp2 = 10'd516; a_exp3 = 10'd616;
b_exp0 = 10'd399; b_exp1 = 10'd447; b_exp2 = 10'd107; b_exp3 = 10'd885;
a_sign0 = 4'd12; a_sign1 = 4'd6; a_sign2 = 4'd13; a_sign3 = 4'd5;
b_sign0 = 4'd0; b_sign1 = 4'd11; b_sign2 = 4'd8; b_sign3 = 4'd12;
@(posedge clk_i);
a_mant0 = 8'd85; a_mant1 = 8'd179; a_mant2 = 8'd5; a_mant3 = 8'd8;
b_mant0 = 8'd7; b_mant1 = 8'd50; b_mant2 = 8'd236; b_mant3 = 8'd70;
a_exp0 = 10'd93; a_exp1 = 10'd409; a_exp2 = 10'd383; a_exp3 = 10'd126;
b_exp0 = 10'd978; b_exp1 = 10'd754; b_exp2 = 10'd690; b_exp3 = 10'd847;
a_sign0 = 4'd8; a_sign1 = 4'd6; a_sign2 = 4'd15; a_sign3 = 4'd2;
b_sign0 = 4'd8; b_sign1 = 4'd2; b_sign2 = 4'd9; b_sign3 = 4'd5;
@(posedge clk_i);
a_mant0 = 8'd214; a_mant1 = 8'd2; a_mant2 = 8'd51; a_mant3 = 8'd219;
b_mant0 = 8'd253; b_mant1 = 8'd145; b_mant2 = 8'd91; b_mant3 = 8'd172;
a_exp0 = 10'd889; a_exp1 = 10'd122; a_exp2 = 10'd859; a_exp3 = 10'd704;
b_exp0 = 10'd854; b_exp1 = 10'd670; b_exp2 = 10'd254; b_exp3 = 10'd641;
a_sign0 = 4'd7; a_sign1 = 4'd3; a_sign2 = 4'd0; a_sign3 = 4'd5;
b_sign0 = 4'd6; b_sign1 = 4'd1; b_sign2 = 4'd12; b_sign3 = 4'd14;
@(posedge clk_i);
a_mant0 = 8'd101; a_mant1 = 8'd40; a_mant2 = 8'd48; a_mant3 = 8'd12;
b_mant0 = 8'd172; b_mant1 = 8'd247; b_mant2 = 8'd156; b_mant3 = 8'd217;
a_exp0 = 10'd619; a_exp1 = 10'd389; a_exp2 = 10'd735; a_exp3 = 10'd907;
b_exp0 = 10'd797; b_exp1 = 10'd52; b_exp2 = 10'd445; b_exp3 = 10'd612;
a_sign0 = 4'd2; a_sign1 = 4'd0; a_sign2 = 4'd4; a_sign3 = 4'd1;
b_sign0 = 4'd12; b_sign1 = 4'd11; b_sign2 = 4'd3; b_sign3 = 4'd1;
@(posedge clk_i);
a_mant0 = 8'd131; a_mant1 = 8'd53; a_mant2 = 8'd76; a_mant3 = 8'd174;
b_mant0 = 8'd144; b_mant1 = 8'd56; b_mant2 = 8'd147; b_mant3 = 8'd211;
a_exp0 = 10'd878; a_exp1 = 10'd561; a_exp2 = 10'd898; a_exp3 = 10'd375;
b_exp0 = 10'd258; b_exp1 = 10'd100; b_exp2 = 10'd23; b_exp3 = 10'd899;
a_sign0 = 4'd11; a_sign1 = 4'd4; a_sign2 = 4'd12; a_sign3 = 4'd3;
b_sign0 = 4'd15; b_sign1 = 4'd2; b_sign2 = 4'd8; b_sign3 = 4'd2;
@(posedge clk_i);
a_mant0 = 8'd155; a_mant1 = 8'd113; a_mant2 = 8'd2; a_mant3 = 8'd171;
b_mant0 = 8'd251; b_mant1 = 8'd223; b_mant2 = 8'd203; b_mant3 = 8'd107;
a_exp0 = 10'd382; a_exp1 = 10'd684; a_exp2 = 10'd961; a_exp3 = 10'd417;
b_exp0 = 10'd898; b_exp1 = 10'd957; b_exp2 = 10'd527; b_exp3 = 10'd25;
a_sign0 = 4'd6; a_sign1 = 4'd10; a_sign2 = 4'd8; a_sign3 = 4'd2;
b_sign0 = 4'd8; b_sign1 = 4'd7; b_sign2 = 4'd5; b_sign3 = 4'd9;
@(posedge clk_i);
a_mant0 = 8'd180; a_mant1 = 8'd245; a_mant2 = 8'd158; a_mant3 = 8'd22;
b_mant0 = 8'd198; b_mant1 = 8'd14; b_mant2 = 8'd19; b_mant3 = 8'd203;
a_exp0 = 10'd9; a_exp1 = 10'd816; a_exp2 = 10'd26; a_exp3 = 10'd851;
b_exp0 = 10'd141; b_exp1 = 10'd295; b_exp2 = 10'd798; b_exp3 = 10'd280;
a_sign0 = 4'd2; a_sign1 = 4'd12; a_sign2 = 4'd14; a_sign3 = 4'd13;
b_sign0 = 4'd8; b_sign1 = 4'd3; b_sign2 = 4'd9; b_sign3 = 4'd2;
@(posedge clk_i);
shared_exps0 = 8'd132;
shared_exps1 = 8'd116;
rstn = 0;
@(posedge clk_i);
rstn = 1;
a_mant0 = 8'd200; a_mant1 = 8'd95; a_mant2 = 8'd62; a_mant3 = 8'd197;
b_mant0 = 8'd137; b_mant1 = 8'd105; b_mant2 = 8'd125; b_mant3 = 8'd62;
a_exp0 = 10'd423; a_exp1 = 10'd963; a_exp2 = 10'd532; a_exp3 = 10'd420;
b_exp0 = 10'd625; b_exp1 = 10'd226; b_exp2 = 10'd615; b_exp3 = 10'd28;
a_sign0 = 4'd11; a_sign1 = 4'd9; a_sign2 = 4'd13; a_sign3 = 4'd8;
b_sign0 = 4'd15; b_sign1 = 4'd8; b_sign2 = 4'd6; b_sign3 = 4'd15;
@(posedge clk_i);
a_mant0 = 8'd22; a_mant1 = 8'd34; a_mant2 = 8'd238; a_mant3 = 8'd75;
b_mant0 = 8'd212; b_mant1 = 8'd219; b_mant2 = 8'd91; b_mant3 = 8'd236;
a_exp0 = 10'd335; a_exp1 = 10'd419; a_exp2 = 10'd428; a_exp3 = 10'd723;
b_exp0 = 10'd63; b_exp1 = 10'd565; b_exp2 = 10'd102; b_exp3 = 10'd274;
a_sign0 = 4'd2; a_sign1 = 4'd14; a_sign2 = 4'd11; a_sign3 = 4'd4;
b_sign0 = 4'd1; b_sign1 = 4'd10; b_sign2 = 4'd16; b_sign3 = 4'd9;
@(posedge clk_i);
a_mant0 = 8'd165; a_mant1 = 8'd225; a_mant2 = 8'd75; a_mant3 = 8'd67;
b_mant0 = 8'd156; b_mant1 = 8'd128; b_mant2 = 8'd46; b_mant3 = 8'd170;
a_exp0 = 10'd652; a_exp1 = 10'd668; a_exp2 = 10'd889; a_exp3 = 10'd688;
b_exp0 = 10'd739; b_exp1 = 10'd566; b_exp2 = 10'd226; b_exp3 = 10'd512;
a_sign0 = 4'd8; a_sign1 = 4'd6; a_sign2 = 4'd14; a_sign3 = 4'd6;
b_sign0 = 4'd6; b_sign1 = 4'd14; b_sign2 = 4'd15; b_sign3 = 4'd2;
@(posedge clk_i);
a_mant0 = 8'd7; a_mant1 = 8'd131; a_mant2 = 8'd207; a_mant3 = 8'd199;
b_mant0 = 8'd199; b_mant1 = 8'd0; b_mant2 = 8'd52; b_mant3 = 8'd42;
a_exp0 = 10'd19; a_exp1 = 10'd641; a_exp2 = 10'd416; a_exp3 = 10'd871;
b_exp0 = 10'd661; b_exp1 = 10'd179; b_exp2 = 10'd740; b_exp3 = 10'd103;
a_sign0 = 4'd16; a_sign1 = 4'd13; a_sign2 = 4'd4; a_sign3 = 4'd9;
b_sign0 = 4'd6; b_sign1 = 4'd14; b_sign2 = 4'd10; b_sign3 = 4'd10;
@(posedge clk_i);
a_mant0 = 8'd105; a_mant1 = 8'd80; a_mant2 = 8'd17; a_mant3 = 8'd223;
b_mant0 = 8'd49; b_mant1 = 8'd157; b_mant2 = 8'd222; b_mant3 = 8'd228;
a_exp0 = 10'd88; a_exp1 = 10'd533; a_exp2 = 10'd556; a_exp3 = 10'd532;
b_exp0 = 10'd596; b_exp1 = 10'd739; b_exp2 = 10'd350; b_exp3 = 10'd264;
a_sign0 = 4'd7; a_sign1 = 4'd16; a_sign2 = 4'd12; a_sign3 = 4'd12;
b_sign0 = 4'd11; b_sign1 = 4'd11; b_sign2 = 4'd16; b_sign3 = 4'd10;
@(posedge clk_i);
a_mant0 = 8'd221; a_mant1 = 8'd129; a_mant2 = 8'd111; a_mant3 = 8'd211;
b_mant0 = 8'd43; b_mant1 = 8'd146; b_mant2 = 8'd227; b_mant3 = 8'd160;
a_exp0 = 10'd367; a_exp1 = 10'd428; a_exp2 = 10'd389; a_exp3 = 10'd775;
b_exp0 = 10'd480; b_exp1 = 10'd511; b_exp2 = 10'd998; b_exp3 = 10'd742;
a_sign0 = 4'd4; a_sign1 = 4'd15; a_sign2 = 4'd16; a_sign3 = 4'd7;
b_sign0 = 4'd5; b_sign1 = 4'd5; b_sign2 = 4'd15; b_sign3 = 4'd15;
@(posedge clk_i);
a_mant0 = 8'd160; a_mant1 = 8'd60; a_mant2 = 8'd75; a_mant3 = 8'd100;
b_mant0 = 8'd12; b_mant1 = 8'd123; b_mant2 = 8'd41; b_mant3 = 8'd183;
a_exp0 = 10'd995; a_exp1 = 10'd582; a_exp2 = 10'd583; a_exp3 = 10'd791;
b_exp0 = 10'd1004; b_exp1 = 10'd754; b_exp2 = 10'd929; b_exp3 = 10'd510;
a_sign0 = 4'd12; a_sign1 = 4'd5; a_sign2 = 4'd8; a_sign3 = 4'd1;
b_sign0 = 4'd10; b_sign1 = 4'd16; b_sign2 = 4'd12; b_sign3 = 4'd9;
@(posedge clk_i);
shared_exps0 = 8'd114;
shared_exps1 = 8'd143;
a_mant0 = 8'd182; a_mant1 = 8'd67; a_mant2 = 8'd221; a_mant3 = 8'd4;
b_mant0 = 8'd162; b_mant1 = 8'd5; b_mant2 = 8'd144; b_mant3 = 8'd195;
a_exp0 = 10'd851; a_exp1 = 10'd98; a_exp2 = 10'd222; a_exp3 = 10'd133;
b_exp0 = 10'd613; b_exp1 = 10'd573; b_exp2 = 10'd887; b_exp3 = 10'd87;
a_sign0 = 4'd7; a_sign1 = 4'd9; a_sign2 = 4'd3; a_sign3 = 4'd15;
b_sign0 = 4'd3; b_sign1 = 4'd16; b_sign2 = 4'd12; b_sign3 = 4'd8;
@(posedge clk_i);
a_mant0 = 8'd205; a_mant1 = 8'd71; a_mant2 = 8'd26; a_mant3 = 8'd101;
b_mant0 = 8'd135; b_mant1 = 8'd10; b_mant2 = 8'd6; b_mant3 = 8'd162;
a_exp0 = 10'd640; a_exp1 = 10'd121; a_exp2 = 10'd217; a_exp3 = 10'd951;
b_exp0 = 10'd186; b_exp1 = 10'd533; b_exp2 = 10'd356; b_exp3 = 10'd653;
a_sign0 = 4'd15; a_sign1 = 4'd5; a_sign2 = 4'd2; a_sign3 = 4'd9;
b_sign0 = 4'd5; b_sign1 = 4'd16; b_sign2 = 4'd16; b_sign3 = 4'd12;
@(posedge clk_i);
a_mant0 = 8'd47; a_mant1 = 8'd75; a_mant2 = 8'd237; a_mant3 = 8'd244;
b_mant0 = 8'd45; b_mant1 = 8'd106; b_mant2 = 8'd157; b_mant3 = 8'd67;
a_exp0 = 10'd155; a_exp1 = 10'd418; a_exp2 = 10'd27; a_exp3 = 10'd668;
b_exp0 = 10'd368; b_exp1 = 10'd367; b_exp2 = 10'd216; b_exp3 = 10'd758;
a_sign0 = 4'd12; a_sign1 = 4'd5; a_sign2 = 4'd7; a_sign3 = 4'd12;
b_sign0 = 4'd7; b_sign1 = 4'd3; b_sign2 = 4'd6; b_sign3 = 4'd8;
@(posedge clk_i);
a_mant0 = 8'd111; a_mant1 = 8'd201; a_mant2 = 8'd20; a_mant3 = 8'd205;
b_mant0 = 8'd60; b_mant1 = 8'd37; b_mant2 = 8'd101; b_mant3 = 8'd186;
a_exp0 = 10'd790; a_exp1 = 10'd779; a_exp2 = 10'd935; a_exp3 = 10'd510;
b_exp0 = 10'd640; b_exp1 = 10'd615; b_exp2 = 10'd632; b_exp3 = 10'd471;
a_sign0 = 4'd2; a_sign1 = 4'd0; a_sign2 = 4'd1; a_sign3 = 4'd12;
b_sign0 = 4'd8; b_sign1 = 4'd8; b_sign2 = 4'd16; b_sign3 = 4'd3;
@(posedge clk_i);
a_mant0 = 8'd229; a_mant1 = 8'd154; a_mant2 = 8'd37; a_mant3 = 8'd34;
b_mant0 = 8'd227; b_mant1 = 8'd113; b_mant2 = 8'd96; b_mant3 = 8'd70;
a_exp0 = 10'd598; a_exp1 = 10'd1017; a_exp2 = 10'd496; a_exp3 = 10'd803;
b_exp0 = 10'd209; b_exp1 = 10'd199; b_exp2 = 10'd152; b_exp3 = 10'd1010;
a_sign0 = 4'd11; a_sign1 = 4'd16; a_sign2 = 4'd16; a_sign3 = 4'd12;
b_sign0 = 4'd1; b_sign1 = 4'd14; b_sign2 = 4'd7; b_sign3 = 4'd7;
@(posedge clk_i);
a_mant0 = 8'd172; a_mant1 = 8'd2; a_mant2 = 8'd130; a_mant3 = 8'd88;
b_mant0 = 8'd201; b_mant1 = 8'd114; b_mant2 = 8'd144; b_mant3 = 8'd10;
a_exp0 = 10'd849; a_exp1 = 10'd402; a_exp2 = 10'd76; a_exp3 = 10'd127;
b_exp0 = 10'd1; b_exp1 = 10'd216; b_exp2 = 10'd304; b_exp3 = 10'd35;
a_sign0 = 4'd8; a_sign1 = 4'd5; a_sign2 = 4'd11; a_sign3 = 4'd4;
b_sign0 = 4'd16; b_sign1 = 4'd14; b_sign2 = 4'd6; b_sign3 = 4'd0;
@(posedge clk_i);
a_mant0 = 8'd44; a_mant1 = 8'd202; a_mant2 = 8'd92; a_mant3 = 8'd190;
b_mant0 = 8'd197; b_mant1 = 8'd196; b_mant2 = 8'd73; b_mant3 = 8'd109;
a_exp0 = 10'd916; a_exp1 = 10'd812; a_exp2 = 10'd431; a_exp3 = 10'd883;
b_exp0 = 10'd880; b_exp1 = 10'd15; b_exp2 = 10'd293; b_exp3 = 10'd547;
a_sign0 = 4'd5; a_sign1 = 4'd3; a_sign2 = 4'd13; a_sign3 = 4'd16;
b_sign0 = 4'd10; b_sign1 = 4'd14; b_sign2 = 4'd16; b_sign3 = 4'd7;
@(posedge clk_i);
a_mant0 = 8'd237; a_mant1 = 8'd75; a_mant2 = 8'd48; a_mant3 = 8'd85;
b_mant0 = 8'd176; b_mant1 = 8'd247; b_mant2 = 8'd15; b_mant3 = 8'd81;
a_exp0 = 10'd454; a_exp1 = 10'd213; a_exp2 = 10'd988; a_exp3 = 10'd739;
b_exp0 = 10'd258; b_exp1 = 10'd790; b_exp2 = 10'd977; b_exp3 = 10'd973;
a_sign0 = 4'd16; a_sign1 = 4'd7; a_sign2 = 4'd6; a_sign3 = 4'd16;
b_sign0 = 4'd4; b_sign1 = 4'd8; b_sign2 = 4'd14; b_sign3 = 4'd12;
@(posedge clk_i);
shared_exps0 = 8'd109;
shared_exps1 = 8'd120;
a_mant0 = 8'd101; a_mant1 = 8'd8; a_mant2 = 8'd5; a_mant3 = 8'd65;
b_mant0 = 8'd95; b_mant1 = 8'd234; b_mant2 = 8'd49; b_mant3 = 8'd16;
a_exp0 = 10'd289; a_exp1 = 10'd822; a_exp2 = 10'd279; a_exp3 = 10'd90;
b_exp0 = 10'd720; b_exp1 = 10'd654; b_exp2 = 10'd746; b_exp3 = 10'd549;
a_sign0 = 4'd2; a_sign1 = 4'd3; a_sign2 = 4'd5; a_sign3 = 4'd6;
b_sign0 = 4'd4; b_sign1 = 4'd8; b_sign2 = 4'd9; b_sign3 = 4'd0;
@(posedge clk_i);
a_mant0 = 8'd117; a_mant1 = 8'd77; a_mant2 = 8'd138; a_mant3 = 8'd142;
b_mant0 = 8'd26; b_mant1 = 8'd59; b_mant2 = 8'd3; b_mant3 = 8'd164;
a_exp0 = 10'd528; a_exp1 = 10'd7; a_exp2 = 10'd134; a_exp3 = 10'd392;
b_exp0 = 10'd502; b_exp1 = 10'd712; b_exp2 = 10'd890; b_exp3 = 10'd110;
a_sign0 = 4'd9; a_sign1 = 4'd12; a_sign2 = 4'd13; a_sign3 = 4'd1;
b_sign0 = 4'd9; b_sign1 = 4'd8; b_sign2 = 4'd13; b_sign3 = 4'd2;
@(posedge clk_i);
a_mant0 = 8'd208; a_mant1 = 8'd131; a_mant2 = 8'd51; a_mant3 = 8'd225;
b_mant0 = 8'd226; b_mant1 = 8'd111; b_mant2 = 8'd217; b_mant3 = 8'd44;
a_exp0 = 10'd1012; a_exp1 = 10'd368; a_exp2 = 10'd370; a_exp3 = 10'd428;
b_exp0 = 10'd911; b_exp1 = 10'd296; b_exp2 = 10'd395; b_exp3 = 10'd121;
a_sign0 = 4'd10; a_sign1 = 4'd7; a_sign2 = 4'd10; a_sign3 = 4'd10;
b_sign0 = 4'd13; b_sign1 = 4'd12; b_sign2 = 4'd4; b_sign3 = 4'd0;
@(posedge clk_i);
a_mant0 = 8'd178; a_mant1 = 8'd115; a_mant2 = 8'd194; a_mant3 = 8'd116;
b_mant0 = 8'd26; b_mant1 = 8'd63; b_mant2 = 8'd186; b_mant3 = 8'd205;
a_exp0 = 10'd658; a_exp1 = 10'd254; a_exp2 = 10'd533; a_exp3 = 10'd20;
b_exp0 = 10'd486; b_exp1 = 10'd604; b_exp2 = 10'd247; b_exp3 = 10'd469;
a_sign0 = 4'd5; a_sign1 = 4'd6; a_sign2 = 4'd10; a_sign3 = 4'd6;
b_sign0 = 4'd11; b_sign1 = 4'd0; b_sign2 = 4'd2; b_sign3 = 4'd9;
@(posedge clk_i);
a_mant0 = 8'd152; a_mant1 = 8'd152; a_mant2 = 8'd210; a_mant3 = 8'd177;
b_mant0 = 8'd207; b_mant1 = 8'd112; b_mant2 = 8'd155; b_mant3 = 8'd191;
a_exp0 = 10'd568; a_exp1 = 10'd436; a_exp2 = 10'd957; a_exp3 = 10'd349;
b_exp0 = 10'd223; b_exp1 = 10'd184; b_exp2 = 10'd10; b_exp3 = 10'd327;
a_sign0 = 4'd10; a_sign1 = 4'd2; a_sign2 = 4'd7; a_sign3 = 4'd8;
b_sign0 = 4'd1; b_sign1 = 4'd4; b_sign2 = 4'd1; b_sign3 = 4'd9;
@(posedge clk_i);
a_mant0 = 8'd30; a_mant1 = 8'd199; a_mant2 = 8'd207; a_mant3 = 8'd64;
b_mant0 = 8'd30; b_mant1 = 8'd217; b_mant2 = 8'd252; b_mant3 = 8'd83;
a_exp0 = 10'd420; a_exp1 = 10'd570; a_exp2 = 10'd742; a_exp3 = 10'd467;
b_exp0 = 10'd418; b_exp1 = 10'd914; b_exp2 = 10'd957; b_exp3 = 10'd381;
a_sign0 = 4'd4; a_sign1 = 4'd0; a_sign2 = 4'd4; a_sign3 = 4'd12;
b_sign0 = 4'd0; b_sign1 = 4'd5; b_sign2 = 4'd14; b_sign3 = 4'd6;
@(posedge clk_i);
a_mant0 = 8'd1; a_mant1 = 8'd70; a_mant2 = 8'd82; a_mant3 = 8'd247;
b_mant0 = 8'd61; b_mant1 = 8'd110; b_mant2 = 8'd119; b_mant3 = 8'd142;
a_exp0 = 10'd456; a_exp1 = 10'd832; a_exp2 = 10'd29; a_exp3 = 10'd319;
b_exp0 = 10'd289; b_exp1 = 10'd189; b_exp2 = 10'd163; b_exp3 = 10'd545;
a_sign0 = 4'd0; a_sign1 = 4'd6; a_sign2 = 4'd5; a_sign3 = 4'd6;
b_sign0 = 4'd6; b_sign1 = 4'd11; b_sign2 = 4'd4; b_sign3 = 4'd13;
@(posedge clk_i);
a_mant0 = 8'd213; a_mant1 = 8'd28; a_mant2 = 8'd37; a_mant3 = 8'd89;
b_mant0 = 8'd82; b_mant1 = 8'd244; b_mant2 = 8'd234; b_mant3 = 8'd100;
a_exp0 = 10'd121; a_exp1 = 10'd102; a_exp2 = 10'd681; a_exp3 = 10'd856;
b_exp0 = 10'd988; b_exp1 = 10'd205; b_exp2 = 10'd777; b_exp3 = 10'd492;
a_sign0 = 4'd16; a_sign1 = 4'd13; a_sign2 = 4'd16; a_sign3 = 4'd1;
b_sign0 = 4'd7; b_sign1 = 4'd11; b_sign2 = 4'd16; b_sign3 = 4'd0;
@(posedge clk_i);
shared_exps0 = 8'd129;
shared_exps1 = 8'd128;
a_mant0 = 8'd14; a_mant1 = 8'd147; a_mant2 = 8'd84; a_mant3 = 8'd93;
b_mant0 = 8'd239; b_mant1 = 8'd135; b_mant2 = 8'd40; b_mant3 = 8'd43;
a_exp0 = 10'd952; a_exp1 = 10'd605; a_exp2 = 10'd129; a_exp3 = 10'd223;
b_exp0 = 10'd757; b_exp1 = 10'd499; b_exp2 = 10'd375; b_exp3 = 10'd523;
a_sign0 = 4'd16; a_sign1 = 4'd0; a_sign2 = 4'd16; a_sign3 = 4'd12;
b_sign0 = 4'd10; b_sign1 = 4'd16; b_sign2 = 4'd6; b_sign3 = 4'd12;
@(posedge clk_i);
a_mant0 = 8'd221; a_mant1 = 8'd181; a_mant2 = 8'd60; a_mant3 = 8'd119;
b_mant0 = 8'd48; b_mant1 = 8'd105; b_mant2 = 8'd100; b_mant3 = 8'd150;
a_exp0 = 10'd36; a_exp1 = 10'd865; a_exp2 = 10'd825; a_exp3 = 10'd30;
b_exp0 = 10'd988; b_exp1 = 10'd406; b_exp2 = 10'd640; b_exp3 = 10'd80;
a_sign0 = 4'd2; a_sign1 = 4'd1; a_sign2 = 4'd13; a_sign3 = 4'd6;
b_sign0 = 4'd7; b_sign1 = 4'd5; b_sign2 = 4'd9; b_sign3 = 4'd10;
@(posedge clk_i);
a_mant0 = 8'd52; a_mant1 = 8'd6; a_mant2 = 8'd35; a_mant3 = 8'd126;
b_mant0 = 8'd151; b_mant1 = 8'd40; b_mant2 = 8'd147; b_mant3 = 8'd211;
a_exp0 = 10'd939; a_exp1 = 10'd632; a_exp2 = 10'd540; a_exp3 = 10'd717;
b_exp0 = 10'd228; b_exp1 = 10'd849; b_exp2 = 10'd466; b_exp3 = 10'd337;
a_sign0 = 4'd14; a_sign1 = 4'd13; a_sign2 = 4'd11; a_sign3 = 4'd0;
b_sign0 = 4'd3; b_sign1 = 4'd14; b_sign2 = 4'd5; b_sign3 = 4'd6;
@(posedge clk_i);
a_mant0 = 8'd203; a_mant1 = 8'd81; a_mant2 = 8'd72; a_mant3 = 8'd154;
b_mant0 = 8'd243; b_mant1 = 8'd129; b_mant2 = 8'd204; b_mant3 = 8'd121;
a_exp0 = 10'd599; a_exp1 = 10'd173; a_exp2 = 10'd563; a_exp3 = 10'd485;
b_exp0 = 10'd935; b_exp1 = 10'd395; b_exp2 = 10'd157; b_exp3 = 10'd714;
a_sign0 = 4'd10; a_sign1 = 4'd6; a_sign2 = 4'd10; a_sign3 = 4'd14;
b_sign0 = 4'd14; b_sign1 = 4'd14; b_sign2 = 4'd7; b_sign3 = 4'd2;
@(posedge clk_i);
a_mant0 = 8'd34; a_mant1 = 8'd9; a_mant2 = 8'd101; a_mant3 = 8'd47;
b_mant0 = 8'd189; b_mant1 = 8'd180; b_mant2 = 8'd106; b_mant3 = 8'd213;
a_exp0 = 10'd451; a_exp1 = 10'd366; a_exp2 = 10'd382; a_exp3 = 10'd337;
b_exp0 = 10'd711; b_exp1 = 10'd955; b_exp2 = 10'd416; b_exp3 = 10'd181;
a_sign0 = 4'd0; a_sign1 = 4'd10; a_sign2 = 4'd10; a_sign3 = 4'd2;
b_sign0 = 4'd7; b_sign1 = 4'd9; b_sign2 = 4'd0; b_sign3 = 4'd15;
@(posedge clk_i);
a_mant0 = 8'd77; a_mant1 = 8'd138; a_mant2 = 8'd212; a_mant3 = 8'd69;
b_mant0 = 8'd243; b_mant1 = 8'd124; b_mant2 = 8'd230; b_mant3 = 8'd182;
a_exp0 = 10'd769; a_exp1 = 10'd462; a_exp2 = 10'd194; a_exp3 = 10'd523;
b_exp0 = 10'd229; b_exp1 = 10'd984; b_exp2 = 10'd348; b_exp3 = 10'd297;
a_sign0 = 4'd11; a_sign1 = 4'd15; a_sign2 = 4'd1; a_sign3 = 4'd7;
b_sign0 = 4'd16; b_sign1 = 4'd12; b_sign2 = 4'd7; b_sign3 = 4'd10;
@(posedge clk_i);
a_mant0 = 8'd130; a_mant1 = 8'd247; a_mant2 = 8'd48; a_mant3 = 8'd224;
b_mant0 = 8'd172; b_mant1 = 8'd99; b_mant2 = 8'd168; b_mant3 = 8'd34;
a_exp0 = 10'd674; a_exp1 = 10'd702; a_exp2 = 10'd119; a_exp3 = 10'd141;
b_exp0 = 10'd817; b_exp1 = 10'd830; b_exp2 = 10'd557; b_exp3 = 10'd981;
a_sign0 = 4'd1; a_sign1 = 4'd3; a_sign2 = 4'd8; a_sign3 = 4'd9;
b_sign0 = 4'd1; b_sign1 = 4'd16; b_sign2 = 4'd13; b_sign3 = 4'd9;
@(posedge clk_i);
a_mant0 = 8'd66; a_mant1 = 8'd178; a_mant2 = 8'd122; a_mant3 = 8'd91;
b_mant0 = 8'd1; b_mant1 = 8'd19; b_mant2 = 8'd25; b_mant3 = 8'd150;
a_exp0 = 10'd860; a_exp1 = 10'd228; a_exp2 = 10'd203; a_exp3 = 10'd480;
b_exp0 = 10'd672; b_exp1 = 10'd277; b_exp2 = 10'd25; b_exp3 = 10'd139;
a_sign0 = 4'd3; a_sign1 = 4'd15; a_sign2 = 4'd6; a_sign3 = 4'd9;
b_sign0 = 4'd10; b_sign1 = 4'd4; b_sign2 = 4'd2; b_sign3 = 4'd1;
@(posedge clk_i);
shared_exps0 = 8'd135;
shared_exps1 = 8'd139;
rstn = 0;
@(posedge clk_i);
rstn = 1;
a_mant0 = 8'd110; a_mant1 = 8'd172; a_mant2 = 8'd185; a_mant3 = 8'd93;
b_mant0 = 8'd32; b_mant1 = 8'd116; b_mant2 = 8'd183; b_mant3 = 8'd148;
a_exp0 = 10'd514; a_exp1 = 10'd868; a_exp2 = 10'd889; a_exp3 = 10'd550;
b_exp0 = 10'd585; b_exp1 = 10'd342; b_exp2 = 10'd975; b_exp3 = 10'd276;
a_sign0 = 4'd2; a_sign1 = 4'd8; a_sign2 = 4'd7; a_sign3 = 4'd3;
b_sign0 = 4'd7; b_sign1 = 4'd1; b_sign2 = 4'd16; b_sign3 = 4'd14;
@(posedge clk_i);
a_mant0 = 8'd69; a_mant1 = 8'd184; a_mant2 = 8'd161; a_mant3 = 8'd124;
b_mant0 = 8'd207; b_mant1 = 8'd28; b_mant2 = 8'd201; b_mant3 = 8'd160;
a_exp0 = 10'd63; a_exp1 = 10'd250; a_exp2 = 10'd595; a_exp3 = 10'd262;
b_exp0 = 10'd650; b_exp1 = 10'd311; b_exp2 = 10'd957; b_exp3 = 10'd898;
a_sign0 = 4'd5; a_sign1 = 4'd13; a_sign2 = 4'd4; a_sign3 = 4'd4;
b_sign0 = 4'd7; b_sign1 = 4'd7; b_sign2 = 4'd4; b_sign3 = 4'd4;
@(posedge clk_i);
a_mant0 = 8'd219; a_mant1 = 8'd229; a_mant2 = 8'd252; a_mant3 = 8'd79;
b_mant0 = 8'd225; b_mant1 = 8'd240; b_mant2 = 8'd99; b_mant3 = 8'd220;
a_exp0 = 10'd936; a_exp1 = 10'd635; a_exp2 = 10'd117; a_exp3 = 10'd138;
b_exp0 = 10'd737; b_exp1 = 10'd140; b_exp2 = 10'd681; b_exp3 = 10'd81;
a_sign0 = 4'd16; a_sign1 = 4'd4; a_sign2 = 4'd13; a_sign3 = 4'd0;
b_sign0 = 4'd15; b_sign1 = 4'd14; b_sign2 = 4'd3; b_sign3 = 4'd6;
@(posedge clk_i);
a_mant0 = 8'd99; a_mant1 = 8'd30; a_mant2 = 8'd215; a_mant3 = 8'd109;
b_mant0 = 8'd52; b_mant1 = 8'd194; b_mant2 = 8'd93; b_mant3 = 8'd58;
a_exp0 = 10'd936; a_exp1 = 10'd926; a_exp2 = 10'd816; a_exp3 = 10'd563;
b_exp0 = 10'd414; b_exp1 = 10'd110; b_exp2 = 10'd448; b_exp3 = 10'd789;
a_sign0 = 4'd7; a_sign1 = 4'd15; a_sign2 = 4'd5; a_sign3 = 4'd7;
b_sign0 = 4'd14; b_sign1 = 4'd2; b_sign2 = 4'd15; b_sign3 = 4'd8;
@(posedge clk_i);
a_mant0 = 8'd181; a_mant1 = 8'd217; a_mant2 = 8'd146; a_mant3 = 8'd252;
b_mant0 = 8'd123; b_mant1 = 8'd135; b_mant2 = 8'd31; b_mant3 = 8'd39;
a_exp0 = 10'd790; a_exp1 = 10'd562; a_exp2 = 10'd510; a_exp3 = 10'd274;
b_exp0 = 10'd623; b_exp1 = 10'd412; b_exp2 = 10'd147; b_exp3 = 10'd984;
a_sign0 = 4'd13; a_sign1 = 4'd0; a_sign2 = 4'd2; a_sign3 = 4'd4;
b_sign0 = 4'd2; b_sign1 = 4'd5; b_sign2 = 4'd3; b_sign3 = 4'd16;
@(posedge clk_i);
a_mant0 = 8'd228; a_mant1 = 8'd25; a_mant2 = 8'd59; a_mant3 = 8'd26;
b_mant0 = 8'd112; b_mant1 = 8'd129; b_mant2 = 8'd62; b_mant3 = 8'd37;
a_exp0 = 10'd127; a_exp1 = 10'd536; a_exp2 = 10'd475; a_exp3 = 10'd885;
b_exp0 = 10'd8; b_exp1 = 10'd951; b_exp2 = 10'd239; b_exp3 = 10'd409;
a_sign0 = 4'd4; a_sign1 = 4'd8; a_sign2 = 4'd7; a_sign3 = 4'd6;
b_sign0 = 4'd12; b_sign1 = 4'd8; b_sign2 = 4'd5; b_sign3 = 4'd14;
@(posedge clk_i);
a_mant0 = 8'd56; a_mant1 = 8'd205; a_mant2 = 8'd216; a_mant3 = 8'd104;
b_mant0 = 8'd125; b_mant1 = 8'd43; b_mant2 = 8'd120; b_mant3 = 8'd14;
a_exp0 = 10'd458; a_exp1 = 10'd156; a_exp2 = 10'd622; a_exp3 = 10'd886;
b_exp0 = 10'd615; b_exp1 = 10'd806; b_exp2 = 10'd49; b_exp3 = 10'd726;
a_sign0 = 4'd15; a_sign1 = 4'd5; a_sign2 = 4'd9; a_sign3 = 4'd3;
b_sign0 = 4'd1; b_sign1 = 4'd12; b_sign2 = 4'd10; b_sign3 = 4'd8;
@(posedge clk_i);
shared_exps0 = 8'd127;
shared_exps1 = 8'd145;
a_mant0 = 8'd252; a_mant1 = 8'd243; a_mant2 = 8'd22; a_mant3 = 8'd151;
b_mant0 = 8'd205; b_mant1 = 8'd178; b_mant2 = 8'd156; b_mant3 = 8'd59;
a_exp0 = 10'd285; a_exp1 = 10'd660; a_exp2 = 10'd538; a_exp3 = 10'd968;
b_exp0 = 10'd104; b_exp1 = 10'd780; b_exp2 = 10'd327; b_exp3 = 10'd726;
a_sign0 = 4'd16; a_sign1 = 4'd2; a_sign2 = 4'd4; a_sign3 = 4'd15;
b_sign0 = 4'd12; b_sign1 = 4'd4; b_sign2 = 4'd15; b_sign3 = 4'd14;
@(posedge clk_i);
a_mant0 = 8'd229; a_mant1 = 8'd43; a_mant2 = 8'd31; a_mant3 = 8'd195;
b_mant0 = 8'd113; b_mant1 = 8'd7; b_mant2 = 8'd75; b_mant3 = 8'd193;
a_exp0 = 10'd553; a_exp1 = 10'd566; a_exp2 = 10'd32; a_exp3 = 10'd425;
b_exp0 = 10'd53; b_exp1 = 10'd427; b_exp2 = 10'd454; b_exp3 = 10'd177;
a_sign0 = 4'd5; a_sign1 = 4'd9; a_sign2 = 4'd10; a_sign3 = 4'd1;
b_sign0 = 4'd2; b_sign1 = 4'd4; b_sign2 = 4'd14; b_sign3 = 4'd7;
@(posedge clk_i);
a_mant0 = 8'd178; a_mant1 = 8'd3; a_mant2 = 8'd112; a_mant3 = 8'd230;
b_mant0 = 8'd212; b_mant1 = 8'd138; b_mant2 = 8'd54; b_mant3 = 8'd40;
a_exp0 = 10'd744; a_exp1 = 10'd608; a_exp2 = 10'd883; a_exp3 = 10'd975;
b_exp0 = 10'd324; b_exp1 = 10'd956; b_exp2 = 10'd805; b_exp3 = 10'd410;
a_sign0 = 4'd9; a_sign1 = 4'd3; a_sign2 = 4'd3; a_sign3 = 4'd0;
b_sign0 = 4'd4; b_sign1 = 4'd10; b_sign2 = 4'd3; b_sign3 = 4'd11;
@(posedge clk_i);
a_mant0 = 8'd107; a_mant1 = 8'd205; a_mant2 = 8'd187; a_mant3 = 8'd224;
b_mant0 = 8'd164; b_mant1 = 8'd153; b_mant2 = 8'd115; b_mant3 = 8'd60;
a_exp0 = 10'd209; a_exp1 = 10'd579; a_exp2 = 10'd99; a_exp3 = 10'd773;
b_exp0 = 10'd472; b_exp1 = 10'd153; b_exp2 = 10'd725; b_exp3 = 10'd640;
a_sign0 = 4'd8; a_sign1 = 4'd6; a_sign2 = 4'd5; a_sign3 = 4'd9;
b_sign0 = 4'd5; b_sign1 = 4'd7; b_sign2 = 4'd5; b_sign3 = 4'd14;
@(posedge clk_i);
a_mant0 = 8'd152; a_mant1 = 8'd218; a_mant2 = 8'd211; a_mant3 = 8'd180;
b_mant0 = 8'd160; b_mant1 = 8'd255; b_mant2 = 8'd174; b_mant3 = 8'd27;
a_exp0 = 10'd370; a_exp1 = 10'd548; a_exp2 = 10'd852; a_exp3 = 10'd112;
b_exp0 = 10'd813; b_exp1 = 10'd689; b_exp2 = 10'd155; b_exp3 = 10'd934;
a_sign0 = 4'd11; a_sign1 = 4'd10; a_sign2 = 4'd1; a_sign3 = 4'd3;
b_sign0 = 4'd14; b_sign1 = 4'd4; b_sign2 = 4'd7; b_sign3 = 4'd12;
@(posedge clk_i);
a_mant0 = 8'd19; a_mant1 = 8'd207; a_mant2 = 8'd114; a_mant3 = 8'd251;
b_mant0 = 8'd85; b_mant1 = 8'd1; b_mant2 = 8'd99; b_mant3 = 8'd255;
a_exp0 = 10'd474; a_exp1 = 10'd271; a_exp2 = 10'd406; a_exp3 = 10'd971;
b_exp0 = 10'd349; b_exp1 = 10'd110; b_exp2 = 10'd518; b_exp3 = 10'd769;
a_sign0 = 4'd16; a_sign1 = 4'd11; a_sign2 = 4'd8; a_sign3 = 4'd2;
b_sign0 = 4'd4; b_sign1 = 4'd11; b_sign2 = 4'd16; b_sign3 = 4'd4;
@(posedge clk_i);
a_mant0 = 8'd174; a_mant1 = 8'd233; a_mant2 = 8'd159; a_mant3 = 8'd130;
b_mant0 = 8'd70; b_mant1 = 8'd5; b_mant2 = 8'd138; b_mant3 = 8'd58;
a_exp0 = 10'd366; a_exp1 = 10'd272; a_exp2 = 10'd325; a_exp3 = 10'd13;
b_exp0 = 10'd799; b_exp1 = 10'd913; b_exp2 = 10'd215; b_exp3 = 10'd264;
a_sign0 = 4'd3; a_sign1 = 4'd15; a_sign2 = 4'd5; a_sign3 = 4'd2;
b_sign0 = 4'd7; b_sign1 = 4'd7; b_sign2 = 4'd15; b_sign3 = 4'd13;
@(posedge clk_i);
a_mant0 = 8'd52; a_mant1 = 8'd229; a_mant2 = 8'd69; a_mant3 = 8'd137;
b_mant0 = 8'd68; b_mant1 = 8'd217; b_mant2 = 8'd179; b_mant3 = 8'd118;
a_exp0 = 10'd149; a_exp1 = 10'd555; a_exp2 = 10'd538; a_exp3 = 10'd950;
b_exp0 = 10'd739; b_exp1 = 10'd927; b_exp2 = 10'd116; b_exp3 = 10'd703;
a_sign0 = 4'd9; a_sign1 = 4'd11; a_sign2 = 4'd3; a_sign3 = 4'd10;
b_sign0 = 4'd4; b_sign1 = 4'd5; b_sign2 = 4'd7; b_sign3 = 4'd6;
@(posedge clk_i);
shared_exps0 = 8'd110;
shared_exps1 = 8'd105;
a_mant0 = 8'd59; a_mant1 = 8'd236; a_mant2 = 8'd230; a_mant3 = 8'd175;
b_mant0 = 8'd77; b_mant1 = 8'd111; b_mant2 = 8'd251; b_mant3 = 8'd114;
a_exp0 = 10'd886; a_exp1 = 10'd78; a_exp2 = 10'd194; a_exp3 = 10'd804;
b_exp0 = 10'd727; b_exp1 = 10'd366; b_exp2 = 10'd412; b_exp3 = 10'd528;
a_sign0 = 4'd7; a_sign1 = 4'd4; a_sign2 = 4'd12; a_sign3 = 4'd3;
b_sign0 = 4'd0; b_sign1 = 4'd8; b_sign2 = 4'd0; b_sign3 = 4'd5;
@(posedge clk_i);
a_mant0 = 8'd26; a_mant1 = 8'd252; a_mant2 = 8'd232; a_mant3 = 8'd60;
b_mant0 = 8'd10; b_mant1 = 8'd61; b_mant2 = 8'd115; b_mant3 = 8'd137;
a_exp0 = 10'd512; a_exp1 = 10'd829; a_exp2 = 10'd818; a_exp3 = 10'd493;
b_exp0 = 10'd541; b_exp1 = 10'd940; b_exp2 = 10'd967; b_exp3 = 10'd60;
a_sign0 = 4'd15; a_sign1 = 4'd13; a_sign2 = 4'd2; a_sign3 = 4'd13;
b_sign0 = 4'd3; b_sign1 = 4'd13; b_sign2 = 4'd11; b_sign3 = 4'd13;
@(posedge clk_i);
a_mant0 = 8'd134; a_mant1 = 8'd41; a_mant2 = 8'd45; a_mant3 = 8'd197;
b_mant0 = 8'd78; b_mant1 = 8'd148; b_mant2 = 8'd213; b_mant3 = 8'd98;
a_exp0 = 10'd170; a_exp1 = 10'd208; a_exp2 = 10'd469; a_exp3 = 10'd637;
b_exp0 = 10'd943; b_exp1 = 10'd483; b_exp2 = 10'd493; b_exp3 = 10'd316;
a_sign0 = 4'd9; a_sign1 = 4'd3; a_sign2 = 4'd3; a_sign3 = 4'd16;
b_sign0 = 4'd11; b_sign1 = 4'd16; b_sign2 = 4'd16; b_sign3 = 4'd10;
@(posedge clk_i);
a_mant0 = 8'd27; a_mant1 = 8'd123; a_mant2 = 8'd134; a_mant3 = 8'd225;
b_mant0 = 8'd58; b_mant1 = 8'd181; b_mant2 = 8'd3; b_mant3 = 8'd122;
a_exp0 = 10'd795; a_exp1 = 10'd445; a_exp2 = 10'd814; a_exp3 = 10'd743;
b_exp0 = 10'd882; b_exp1 = 10'd541; b_exp2 = 10'd657; b_exp3 = 10'd343;
a_sign0 = 4'd15; a_sign1 = 4'd13; a_sign2 = 4'd5; a_sign3 = 4'd9;
b_sign0 = 4'd16; b_sign1 = 4'd10; b_sign2 = 4'd13; b_sign3 = 4'd8;
@(posedge clk_i);
a_mant0 = 8'd41; a_mant1 = 8'd96; a_mant2 = 8'd174; a_mant3 = 8'd254;
b_mant0 = 8'd241; b_mant1 = 8'd249; b_mant2 = 8'd158; b_mant3 = 8'd121;
a_exp0 = 10'd291; a_exp1 = 10'd757; a_exp2 = 10'd836; a_exp3 = 10'd534;
b_exp0 = 10'd134; b_exp1 = 10'd498; b_exp2 = 10'd760; b_exp3 = 10'd738;
a_sign0 = 4'd1; a_sign1 = 4'd7; a_sign2 = 4'd9; a_sign3 = 4'd9;
b_sign0 = 4'd16; b_sign1 = 4'd10; b_sign2 = 4'd1; b_sign3 = 4'd5;
@(posedge clk_i);
a_mant0 = 8'd173; a_mant1 = 8'd78; a_mant2 = 8'd244; a_mant3 = 8'd221;
b_mant0 = 8'd114; b_mant1 = 8'd85; b_mant2 = 8'd95; b_mant3 = 8'd248;
a_exp0 = 10'd860; a_exp1 = 10'd351; a_exp2 = 10'd350; a_exp3 = 10'd915;
b_exp0 = 10'd193; b_exp1 = 10'd672; b_exp2 = 10'd883; b_exp3 = 10'd700;
a_sign0 = 4'd12; a_sign1 = 4'd7; a_sign2 = 4'd11; a_sign3 = 4'd9;
b_sign0 = 4'd5; b_sign1 = 4'd11; b_sign2 = 4'd5; b_sign3 = 4'd6;
@(posedge clk_i);
a_mant0 = 8'd83; a_mant1 = 8'd25; a_mant2 = 8'd252; a_mant3 = 8'd24;
b_mant0 = 8'd75; b_mant1 = 8'd122; b_mant2 = 8'd81; b_mant3 = 8'd148;
a_exp0 = 10'd817; a_exp1 = 10'd750; a_exp2 = 10'd375; a_exp3 = 10'd492;
b_exp0 = 10'd97; b_exp1 = 10'd993; b_exp2 = 10'd631; b_exp3 = 10'd584;
a_sign0 = 4'd2; a_sign1 = 4'd10; a_sign2 = 4'd7; a_sign3 = 4'd13;
b_sign0 = 4'd11; b_sign1 = 4'd1; b_sign2 = 4'd1; b_sign3 = 4'd2;
@(posedge clk_i);
a_mant0 = 8'd41; a_mant1 = 8'd227; a_mant2 = 8'd251; a_mant3 = 8'd253;
b_mant0 = 8'd61; b_mant1 = 8'd194; b_mant2 = 8'd138; b_mant3 = 8'd127;
a_exp0 = 10'd517; a_exp1 = 10'd720; a_exp2 = 10'd966; a_exp3 = 10'd38;
b_exp0 = 10'd441; b_exp1 = 10'd747; b_exp2 = 10'd565; b_exp3 = 10'd924;
a_sign0 = 4'd12; a_sign1 = 4'd7; a_sign2 = 4'd7; a_sign3 = 4'd3;
b_sign0 = 4'd16; b_sign1 = 4'd4; b_sign2 = 4'd9; b_sign3 = 4'd12;
@(posedge clk_i);
shared_exps0 = 8'd131;
shared_exps1 = 8'd119;
a_mant0 = 8'd80; a_mant1 = 8'd86; a_mant2 = 8'd99; a_mant3 = 8'd62;
b_mant0 = 8'd81; b_mant1 = 8'd22; b_mant2 = 8'd178; b_mant3 = 8'd187;
a_exp0 = 10'd226; a_exp1 = 10'd276; a_exp2 = 10'd345; a_exp3 = 10'd507;
b_exp0 = 10'd764; b_exp1 = 10'd758; b_exp2 = 10'd855; b_exp3 = 10'd602;
a_sign0 = 4'd9; a_sign1 = 4'd0; a_sign2 = 4'd13; a_sign3 = 4'd10;
b_sign0 = 4'd15; b_sign1 = 4'd3; b_sign2 = 4'd15; b_sign3 = 4'd16;
@(posedge clk_i);
a_mant0 = 8'd199; a_mant1 = 8'd80; a_mant2 = 8'd170; a_mant3 = 8'd65;
b_mant0 = 8'd209; b_mant1 = 8'd51; b_mant2 = 8'd243; b_mant3 = 8'd88;
a_exp0 = 10'd259; a_exp1 = 10'd598; a_exp2 = 10'd442; a_exp3 = 10'd511;
b_exp0 = 10'd686; b_exp1 = 10'd626; b_exp2 = 10'd753; b_exp3 = 10'd534;
a_sign0 = 4'd16; a_sign1 = 4'd13; a_sign2 = 4'd16; a_sign3 = 4'd6;
b_sign0 = 4'd10; b_sign1 = 4'd12; b_sign2 = 4'd5; b_sign3 = 4'd5;
@(posedge clk_i);
a_mant0 = 8'd139; a_mant1 = 8'd186; a_mant2 = 8'd47; a_mant3 = 8'd36;
b_mant0 = 8'd250; b_mant1 = 8'd204; b_mant2 = 8'd79; b_mant3 = 8'd229;
a_exp0 = 10'd949; a_exp1 = 10'd94; a_exp2 = 10'd107; a_exp3 = 10'd285;
b_exp0 = 10'd910; b_exp1 = 10'd919; b_exp2 = 10'd454; b_exp3 = 10'd411;
a_sign0 = 4'd8; a_sign1 = 4'd14; a_sign2 = 4'd7; a_sign3 = 4'd2;
b_sign0 = 4'd15; b_sign1 = 4'd6; b_sign2 = 4'd10; b_sign3 = 4'd1;
@(posedge clk_i);
a_mant0 = 8'd24; a_mant1 = 8'd163; a_mant2 = 8'd222; a_mant3 = 8'd124;
b_mant0 = 8'd156; b_mant1 = 8'd116; b_mant2 = 8'd100; b_mant3 = 8'd26;
a_exp0 = 10'd818; a_exp1 = 10'd503; a_exp2 = 10'd492; a_exp3 = 10'd983;
b_exp0 = 10'd650; b_exp1 = 10'd6; b_exp2 = 10'd330; b_exp3 = 10'd849;
a_sign0 = 4'd2; a_sign1 = 4'd5; a_sign2 = 4'd3; a_sign3 = 4'd16;
b_sign0 = 4'd12; b_sign1 = 4'd5; b_sign2 = 4'd9; b_sign3 = 4'd6;
@(posedge clk_i);
a_mant0 = 8'd220; a_mant1 = 8'd181; a_mant2 = 8'd123; a_mant3 = 8'd208;
b_mant0 = 8'd162; b_mant1 = 8'd148; b_mant2 = 8'd106; b_mant3 = 8'd238;
a_exp0 = 10'd421; a_exp1 = 10'd1003; a_exp2 = 10'd987; a_exp3 = 10'd351;
b_exp0 = 10'd590; b_exp1 = 10'd407; b_exp2 = 10'd703; b_exp3 = 10'd219;
a_sign0 = 4'd8; a_sign1 = 4'd11; a_sign2 = 4'd6; a_sign3 = 4'd0;
b_sign0 = 4'd8; b_sign1 = 4'd7; b_sign2 = 4'd13; b_sign3 = 4'd5;
@(posedge clk_i);
a_mant0 = 8'd157; a_mant1 = 8'd181; a_mant2 = 8'd134; a_mant3 = 8'd152;
b_mant0 = 8'd61; b_mant1 = 8'd90; b_mant2 = 8'd134; b_mant3 = 8'd58;
a_exp0 = 10'd213; a_exp1 = 10'd519; a_exp2 = 10'd375; a_exp3 = 10'd566;
b_exp0 = 10'd674; b_exp1 = 10'd806; b_exp2 = 10'd838; b_exp3 = 10'd430;
a_sign0 = 4'd10; a_sign1 = 4'd15; a_sign2 = 4'd12; a_sign3 = 4'd7;
b_sign0 = 4'd11; b_sign1 = 4'd15; b_sign2 = 4'd2; b_sign3 = 4'd11;
@(posedge clk_i);
a_mant0 = 8'd212; a_mant1 = 8'd241; a_mant2 = 8'd52; a_mant3 = 8'd6;
b_mant0 = 8'd99; b_mant1 = 8'd99; b_mant2 = 8'd194; b_mant3 = 8'd197;
a_exp0 = 10'd590; a_exp1 = 10'd406; a_exp2 = 10'd914; a_exp3 = 10'd54;
b_exp0 = 10'd261; b_exp1 = 10'd574; b_exp2 = 10'd534; b_exp3 = 10'd370;
a_sign0 = 4'd11; a_sign1 = 4'd1; a_sign2 = 4'd16; a_sign3 = 4'd16;
b_sign0 = 4'd15; b_sign1 = 4'd12; b_sign2 = 4'd0; b_sign3 = 4'd4;
@(posedge clk_i);
a_mant0 = 8'd56; a_mant1 = 8'd31; a_mant2 = 8'd101; a_mant3 = 8'd43;
b_mant0 = 8'd153; b_mant1 = 8'd31; b_mant2 = 8'd129; b_mant3 = 8'd48;
a_exp0 = 10'd323; a_exp1 = 10'd463; a_exp2 = 10'd584; a_exp3 = 10'd380;
b_exp0 = 10'd989; b_exp1 = 10'd924; b_exp2 = 10'd969; b_exp3 = 10'd943;
a_sign0 = 4'd2; a_sign1 = 4'd16; a_sign2 = 4'd4; a_sign3 = 4'd0;
b_sign0 = 4'd8; b_sign1 = 4'd15; b_sign2 = 4'd12; b_sign3 = 4'd0;
@(posedge clk_i);
shared_exps0 = 8'd135;
shared_exps1 = 8'd127;
rstn = 0;
@(posedge clk_i);
rstn = 1;
a_mant0 = 8'd17; a_mant1 = 8'd172; a_mant2 = 8'd48; a_mant3 = 8'd1;
b_mant0 = 8'd97; b_mant1 = 8'd72; b_mant2 = 8'd181; b_mant3 = 8'd251;
a_exp0 = 10'd306; a_exp1 = 10'd233; a_exp2 = 10'd463; a_exp3 = 10'd551;
b_exp0 = 10'd608; b_exp1 = 10'd636; b_exp2 = 10'd433; b_exp3 = 10'd178;
a_sign0 = 4'd8; a_sign1 = 4'd0; a_sign2 = 4'd3; a_sign3 = 4'd7;
b_sign0 = 4'd10; b_sign1 = 4'd4; b_sign2 = 4'd2; b_sign3 = 4'd0;
@(posedge clk_i);
a_mant0 = 8'd18; a_mant1 = 8'd78; a_mant2 = 8'd117; a_mant3 = 8'd170;
b_mant0 = 8'd52; b_mant1 = 8'd137; b_mant2 = 8'd83; b_mant3 = 8'd199;
a_exp0 = 10'd497; a_exp1 = 10'd307; a_exp2 = 10'd961; a_exp3 = 10'd165;
b_exp0 = 10'd381; b_exp1 = 10'd692; b_exp2 = 10'd62; b_exp3 = 10'd315;
a_sign0 = 4'd15; a_sign1 = 4'd10; a_sign2 = 4'd11; a_sign3 = 4'd13;
b_sign0 = 4'd10; b_sign1 = 4'd2; b_sign2 = 4'd16; b_sign3 = 4'd13;
@(posedge clk_i);
a_mant0 = 8'd230; a_mant1 = 8'd0; a_mant2 = 8'd19; a_mant3 = 8'd147;
b_mant0 = 8'd71; b_mant1 = 8'd64; b_mant2 = 8'd50; b_mant3 = 8'd116;
a_exp0 = 10'd810; a_exp1 = 10'd629; a_exp2 = 10'd386; a_exp3 = 10'd149;
b_exp0 = 10'd909; b_exp1 = 10'd804; b_exp2 = 10'd925; b_exp3 = 10'd373;
a_sign0 = 4'd10; a_sign1 = 4'd10; a_sign2 = 4'd7; a_sign3 = 4'd11;
b_sign0 = 4'd4; b_sign1 = 4'd11; b_sign2 = 4'd16; b_sign3 = 4'd3;
@(posedge clk_i);
a_mant0 = 8'd125; a_mant1 = 8'd122; a_mant2 = 8'd208; a_mant3 = 8'd26;
b_mant0 = 8'd172; b_mant1 = 8'd83; b_mant2 = 8'd79; b_mant3 = 8'd46;
a_exp0 = 10'd140; a_exp1 = 10'd196; a_exp2 = 10'd387; a_exp3 = 10'd810;
b_exp0 = 10'd752; b_exp1 = 10'd496; b_exp2 = 10'd867; b_exp3 = 10'd737;
a_sign0 = 4'd8; a_sign1 = 4'd13; a_sign2 = 4'd5; a_sign3 = 4'd2;
b_sign0 = 4'd16; b_sign1 = 4'd16; b_sign2 = 4'd13; b_sign3 = 4'd12;
@(posedge clk_i);
a_mant0 = 8'd205; a_mant1 = 8'd254; a_mant2 = 8'd242; a_mant3 = 8'd128;
b_mant0 = 8'd161; b_mant1 = 8'd99; b_mant2 = 8'd97; b_mant3 = 8'd7;
a_exp0 = 10'd676; a_exp1 = 10'd835; a_exp2 = 10'd805; a_exp3 = 10'd496;
b_exp0 = 10'd689; b_exp1 = 10'd623; b_exp2 = 10'd885; b_exp3 = 10'd128;
a_sign0 = 4'd6; a_sign1 = 4'd7; a_sign2 = 4'd2; a_sign3 = 4'd12;
b_sign0 = 4'd2; b_sign1 = 4'd5; b_sign2 = 4'd4; b_sign3 = 4'd0;
@(posedge clk_i);
a_mant0 = 8'd32; a_mant1 = 8'd89; a_mant2 = 8'd232; a_mant3 = 8'd97;
b_mant0 = 8'd138; b_mant1 = 8'd55; b_mant2 = 8'd212; b_mant3 = 8'd228;
a_exp0 = 10'd9; a_exp1 = 10'd25; a_exp2 = 10'd848; a_exp3 = 10'd94;
b_exp0 = 10'd985; b_exp1 = 10'd1014; b_exp2 = 10'd984; b_exp3 = 10'd256;
a_sign0 = 4'd5; a_sign1 = 4'd1; a_sign2 = 4'd8; a_sign3 = 4'd15;
b_sign0 = 4'd2; b_sign1 = 4'd6; b_sign2 = 4'd6; b_sign3 = 4'd13;
@(posedge clk_i);
a_mant0 = 8'd32; a_mant1 = 8'd183; a_mant2 = 8'd97; a_mant3 = 8'd78;
b_mant0 = 8'd166; b_mant1 = 8'd231; b_mant2 = 8'd75; b_mant3 = 8'd199;
a_exp0 = 10'd51; a_exp1 = 10'd967; a_exp2 = 10'd115; a_exp3 = 10'd444;
b_exp0 = 10'd446; b_exp1 = 10'd352; b_exp2 = 10'd81; b_exp3 = 10'd559;
a_sign0 = 4'd1; a_sign1 = 4'd7; a_sign2 = 4'd4; a_sign3 = 4'd0;
b_sign0 = 4'd8; b_sign1 = 4'd10; b_sign2 = 4'd12; b_sign3 = 4'd6;
@(posedge clk_i);
shared_exps0 = 8'd132;
shared_exps1 = 8'd104;
a_mant0 = 8'd117; a_mant1 = 8'd208; a_mant2 = 8'd168; a_mant3 = 8'd163;
b_mant0 = 8'd172; b_mant1 = 8'd255; b_mant2 = 8'd203; b_mant3 = 8'd144;
a_exp0 = 10'd107; a_exp1 = 10'd352; a_exp2 = 10'd122; a_exp3 = 10'd733;
b_exp0 = 10'd698; b_exp1 = 10'd310; b_exp2 = 10'd255; b_exp3 = 10'd326;
a_sign0 = 4'd4; a_sign1 = 4'd5; a_sign2 = 4'd4; a_sign3 = 4'd14;
b_sign0 = 4'd5; b_sign1 = 4'd12; b_sign2 = 4'd12; b_sign3 = 4'd7;
@(posedge clk_i);
a_mant0 = 8'd151; a_mant1 = 8'd19; a_mant2 = 8'd52; a_mant3 = 8'd92;
b_mant0 = 8'd31; b_mant1 = 8'd176; b_mant2 = 8'd123; b_mant3 = 8'd163;
a_exp0 = 10'd672; a_exp1 = 10'd988; a_exp2 = 10'd949; a_exp3 = 10'd204;
b_exp0 = 10'd984; b_exp1 = 10'd922; b_exp2 = 10'd533; b_exp3 = 10'd186;
a_sign0 = 4'd11; a_sign1 = 4'd15; a_sign2 = 4'd3; a_sign3 = 4'd0;
b_sign0 = 4'd11; b_sign1 = 4'd6; b_sign2 = 4'd8; b_sign3 = 4'd16;
@(posedge clk_i);
a_mant0 = 8'd163; a_mant1 = 8'd220; a_mant2 = 8'd209; a_mant3 = 8'd30;
b_mant0 = 8'd55; b_mant1 = 8'd119; b_mant2 = 8'd203; b_mant3 = 8'd243;
a_exp0 = 10'd75; a_exp1 = 10'd45; a_exp2 = 10'd336; a_exp3 = 10'd822;
b_exp0 = 10'd127; b_exp1 = 10'd498; b_exp2 = 10'd671; b_exp3 = 10'd906;
a_sign0 = 4'd15; a_sign1 = 4'd5; a_sign2 = 4'd6; a_sign3 = 4'd7;
b_sign0 = 4'd2; b_sign1 = 4'd12; b_sign2 = 4'd1; b_sign3 = 4'd8;
@(posedge clk_i);
a_mant0 = 8'd155; a_mant1 = 8'd73; a_mant2 = 8'd95; a_mant3 = 8'd87;
b_mant0 = 8'd203; b_mant1 = 8'd7; b_mant2 = 8'd136; b_mant3 = 8'd76;
a_exp0 = 10'd362; a_exp1 = 10'd315; a_exp2 = 10'd729; a_exp3 = 10'd821;
b_exp0 = 10'd455; b_exp1 = 10'd577; b_exp2 = 10'd602; b_exp3 = 10'd860;
a_sign0 = 4'd3; a_sign1 = 4'd6; a_sign2 = 4'd8; a_sign3 = 4'd10;
b_sign0 = 4'd13; b_sign1 = 4'd0; b_sign2 = 4'd9; b_sign3 = 4'd5;
@(posedge clk_i);
a_mant0 = 8'd117; a_mant1 = 8'd63; a_mant2 = 8'd118; a_mant3 = 8'd66;
b_mant0 = 8'd70; b_mant1 = 8'd89; b_mant2 = 8'd159; b_mant3 = 8'd207;
a_exp0 = 10'd800; a_exp1 = 10'd167; a_exp2 = 10'd224; a_exp3 = 10'd486;
b_exp0 = 10'd680; b_exp1 = 10'd287; b_exp2 = 10'd444; b_exp3 = 10'd633;
a_sign0 = 4'd10; a_sign1 = 4'd8; a_sign2 = 4'd10; a_sign3 = 4'd1;
b_sign0 = 4'd10; b_sign1 = 4'd11; b_sign2 = 4'd0; b_sign3 = 4'd9;
@(posedge clk_i);
a_mant0 = 8'd12; a_mant1 = 8'd205; a_mant2 = 8'd154; a_mant3 = 8'd171;
b_mant0 = 8'd163; b_mant1 = 8'd116; b_mant2 = 8'd123; b_mant3 = 8'd75;
a_exp0 = 10'd667; a_exp1 = 10'd194; a_exp2 = 10'd553; a_exp3 = 10'd383;
b_exp0 = 10'd578; b_exp1 = 10'd17; b_exp2 = 10'd549; b_exp3 = 10'd800;
a_sign0 = 4'd0; a_sign1 = 4'd3; a_sign2 = 4'd15; a_sign3 = 4'd8;
b_sign0 = 4'd13; b_sign1 = 4'd2; b_sign2 = 4'd14; b_sign3 = 4'd5;
@(posedge clk_i);
a_mant0 = 8'd62; a_mant1 = 8'd79; a_mant2 = 8'd9; a_mant3 = 8'd145;
b_mant0 = 8'd47; b_mant1 = 8'd250; b_mant2 = 8'd62; b_mant3 = 8'd197;
a_exp0 = 10'd282; a_exp1 = 10'd605; a_exp2 = 10'd216; a_exp3 = 10'd854;
b_exp0 = 10'd98; b_exp1 = 10'd890; b_exp2 = 10'd156; b_exp3 = 10'd320;
a_sign0 = 4'd11; a_sign1 = 4'd14; a_sign2 = 4'd6; a_sign3 = 4'd16;
b_sign0 = 4'd10; b_sign1 = 4'd3; b_sign2 = 4'd16; b_sign3 = 4'd1;
@(posedge clk_i);
a_mant0 = 8'd92; a_mant1 = 8'd90; a_mant2 = 8'd173; a_mant3 = 8'd32;
b_mant0 = 8'd80; b_mant1 = 8'd210; b_mant2 = 8'd130; b_mant3 = 8'd185;
a_exp0 = 10'd717; a_exp1 = 10'd1013; a_exp2 = 10'd967; a_exp3 = 10'd382;
b_exp0 = 10'd620; b_exp1 = 10'd405; b_exp2 = 10'd445; b_exp3 = 10'd933;
a_sign0 = 4'd12; a_sign1 = 4'd12; a_sign2 = 4'd11; a_sign3 = 4'd4;
b_sign0 = 4'd5; b_sign1 = 4'd2; b_sign2 = 4'd3; b_sign3 = 4'd1;
@(posedge clk_i);
shared_exps0 = 8'd129;
shared_exps1 = 8'd110;
a_mant0 = 8'd148; a_mant1 = 8'd37; a_mant2 = 8'd123; a_mant3 = 8'd167;
b_mant0 = 8'd92; b_mant1 = 8'd64; b_mant2 = 8'd67; b_mant3 = 8'd28;
a_exp0 = 10'd428; a_exp1 = 10'd996; a_exp2 = 10'd259; a_exp3 = 10'd164;
b_exp0 = 10'd808; b_exp1 = 10'd29; b_exp2 = 10'd977; b_exp3 = 10'd33;
a_sign0 = 4'd6; a_sign1 = 4'd12; a_sign2 = 4'd6; a_sign3 = 4'd10;
b_sign0 = 4'd14; b_sign1 = 4'd13; b_sign2 = 4'd13; b_sign3 = 4'd13;
@(posedge clk_i);
a_mant0 = 8'd85; a_mant1 = 8'd55; a_mant2 = 8'd206; a_mant3 = 8'd24;
b_mant0 = 8'd153; b_mant1 = 8'd145; b_mant2 = 8'd120; b_mant3 = 8'd158;
a_exp0 = 10'd6; a_exp1 = 10'd571; a_exp2 = 10'd537; a_exp3 = 10'd233;
b_exp0 = 10'd856; b_exp1 = 10'd229; b_exp2 = 10'd742; b_exp3 = 10'd753;
a_sign0 = 4'd10; a_sign1 = 4'd16; a_sign2 = 4'd9; a_sign3 = 4'd6;
b_sign0 = 4'd10; b_sign1 = 4'd9; b_sign2 = 4'd11; b_sign3 = 4'd1;
@(posedge clk_i);
a_mant0 = 8'd119; a_mant1 = 8'd105; a_mant2 = 8'd61; a_mant3 = 8'd124;
b_mant0 = 8'd246; b_mant1 = 8'd188; b_mant2 = 8'd91; b_mant3 = 8'd55;
a_exp0 = 10'd511; a_exp1 = 10'd569; a_exp2 = 10'd1003; a_exp3 = 10'd620;
b_exp0 = 10'd540; b_exp1 = 10'd707; b_exp2 = 10'd171; b_exp3 = 10'd762;
a_sign0 = 4'd3; a_sign1 = 4'd15; a_sign2 = 4'd14; a_sign3 = 4'd16;
b_sign0 = 4'd13; b_sign1 = 4'd7; b_sign2 = 4'd14; b_sign3 = 4'd0;
@(posedge clk_i);
a_mant0 = 8'd119; a_mant1 = 8'd33; a_mant2 = 8'd233; a_mant3 = 8'd205;
b_mant0 = 8'd114; b_mant1 = 8'd222; b_mant2 = 8'd51; b_mant3 = 8'd90;
a_exp0 = 10'd831; a_exp1 = 10'd815; a_exp2 = 10'd152; a_exp3 = 10'd657;
b_exp0 = 10'd904; b_exp1 = 10'd653; b_exp2 = 10'd175; b_exp3 = 10'd477;
a_sign0 = 4'd13; a_sign1 = 4'd14; a_sign2 = 4'd14; a_sign3 = 4'd0;
b_sign0 = 4'd8; b_sign1 = 4'd6; b_sign2 = 4'd15; b_sign3 = 4'd4;
@(posedge clk_i);
a_mant0 = 8'd16; a_mant1 = 8'd214; a_mant2 = 8'd116; a_mant3 = 8'd25;
b_mant0 = 8'd24; b_mant1 = 8'd202; b_mant2 = 8'd43; b_mant3 = 8'd221;
a_exp0 = 10'd165; a_exp1 = 10'd1015; a_exp2 = 10'd226; a_exp3 = 10'd586;
b_exp0 = 10'd254; b_exp1 = 10'd900; b_exp2 = 10'd223; b_exp3 = 10'd789;
a_sign0 = 4'd6; a_sign1 = 4'd4; a_sign2 = 4'd5; a_sign3 = 4'd0;
b_sign0 = 4'd1; b_sign1 = 4'd8; b_sign2 = 4'd3; b_sign3 = 4'd12;
@(posedge clk_i);
a_mant0 = 8'd175; a_mant1 = 8'd225; a_mant2 = 8'd119; a_mant3 = 8'd221;
b_mant0 = 8'd111; b_mant1 = 8'd56; b_mant2 = 8'd65; b_mant3 = 8'd206;
a_exp0 = 10'd786; a_exp1 = 10'd218; a_exp2 = 10'd718; a_exp3 = 10'd600;
b_exp0 = 10'd535; b_exp1 = 10'd543; b_exp2 = 10'd622; b_exp3 = 10'd163;
a_sign0 = 4'd10; a_sign1 = 4'd5; a_sign2 = 4'd13; a_sign3 = 4'd7;
b_sign0 = 4'd16; b_sign1 = 4'd6; b_sign2 = 4'd14; b_sign3 = 4'd7;
@(posedge clk_i);
a_mant0 = 8'd137; a_mant1 = 8'd179; a_mant2 = 8'd170; a_mant3 = 8'd246;
b_mant0 = 8'd98; b_mant1 = 8'd170; b_mant2 = 8'd95; b_mant3 = 8'd242;
a_exp0 = 10'd635; a_exp1 = 10'd206; a_exp2 = 10'd294; a_exp3 = 10'd632;
b_exp0 = 10'd285; b_exp1 = 10'd109; b_exp2 = 10'd542; b_exp3 = 10'd190;
a_sign0 = 4'd13; a_sign1 = 4'd4; a_sign2 = 4'd3; a_sign3 = 4'd5;
b_sign0 = 4'd12; b_sign1 = 4'd6; b_sign2 = 4'd4; b_sign3 = 4'd0;
@(posedge clk_i);
a_mant0 = 8'd170; a_mant1 = 8'd192; a_mant2 = 8'd32; a_mant3 = 8'd76;
b_mant0 = 8'd98; b_mant1 = 8'd136; b_mant2 = 8'd108; b_mant3 = 8'd31;
a_exp0 = 10'd543; a_exp1 = 10'd594; a_exp2 = 10'd283; a_exp3 = 10'd794;
b_exp0 = 10'd33; b_exp1 = 10'd508; b_exp2 = 10'd349; b_exp3 = 10'd684;
a_sign0 = 4'd5; a_sign1 = 4'd5; a_sign2 = 4'd5; a_sign3 = 4'd16;
b_sign0 = 4'd3; b_sign1 = 4'd8; b_sign2 = 4'd2; b_sign3 = 4'd11;
@(posedge clk_i);
shared_exps0 = 8'd115;
shared_exps1 = 8'd106;
a_mant0 = 8'd185; a_mant1 = 8'd170; a_mant2 = 8'd80; a_mant3 = 8'd4;
b_mant0 = 8'd43; b_mant1 = 8'd111; b_mant2 = 8'd19; b_mant3 = 8'd180;
a_exp0 = 10'd596; a_exp1 = 10'd328; a_exp2 = 10'd270; a_exp3 = 10'd249;
b_exp0 = 10'd139; b_exp1 = 10'd627; b_exp2 = 10'd388; b_exp3 = 10'd1021;
a_sign0 = 4'd15; a_sign1 = 4'd6; a_sign2 = 4'd12; a_sign3 = 4'd13;
b_sign0 = 4'd6; b_sign1 = 4'd15; b_sign2 = 4'd4; b_sign3 = 4'd12;
@(posedge clk_i);
a_mant0 = 8'd172; a_mant1 = 8'd102; a_mant2 = 8'd119; a_mant3 = 8'd97;
b_mant0 = 8'd242; b_mant1 = 8'd45; b_mant2 = 8'd41; b_mant3 = 8'd178;
a_exp0 = 10'd381; a_exp1 = 10'd210; a_exp2 = 10'd175; a_exp3 = 10'd794;
b_exp0 = 10'd734; b_exp1 = 10'd778; b_exp2 = 10'd868; b_exp3 = 10'd552;
a_sign0 = 4'd0; a_sign1 = 4'd13; a_sign2 = 4'd9; a_sign3 = 4'd4;
b_sign0 = 4'd15; b_sign1 = 4'd14; b_sign2 = 4'd4; b_sign3 = 4'd3;
@(posedge clk_i);
a_mant0 = 8'd18; a_mant1 = 8'd160; a_mant2 = 8'd94; a_mant3 = 8'd121;
b_mant0 = 8'd201; b_mant1 = 8'd123; b_mant2 = 8'd252; b_mant3 = 8'd114;
a_exp0 = 10'd926; a_exp1 = 10'd850; a_exp2 = 10'd717; a_exp3 = 10'd318;
b_exp0 = 10'd689; b_exp1 = 10'd626; b_exp2 = 10'd543; b_exp3 = 10'd518;
a_sign0 = 4'd1; a_sign1 = 4'd4; a_sign2 = 4'd2; a_sign3 = 4'd7;
b_sign0 = 4'd12; b_sign1 = 4'd0; b_sign2 = 4'd4; b_sign3 = 4'd7;
@(posedge clk_i);
a_mant0 = 8'd239; a_mant1 = 8'd71; a_mant2 = 8'd230; a_mant3 = 8'd199;
b_mant0 = 8'd190; b_mant1 = 8'd238; b_mant2 = 8'd62; b_mant3 = 8'd72;
a_exp0 = 10'd820; a_exp1 = 10'd192; a_exp2 = 10'd863; a_exp3 = 10'd356;
b_exp0 = 10'd974; b_exp1 = 10'd889; b_exp2 = 10'd784; b_exp3 = 10'd615;
a_sign0 = 4'd7; a_sign1 = 4'd4; a_sign2 = 4'd2; a_sign3 = 4'd0;
b_sign0 = 4'd6; b_sign1 = 4'd0; b_sign2 = 4'd11; b_sign3 = 4'd14;
@(posedge clk_i);
a_mant0 = 8'd139; a_mant1 = 8'd140; a_mant2 = 8'd125; a_mant3 = 8'd196;
b_mant0 = 8'd44; b_mant1 = 8'd178; b_mant2 = 8'd184; b_mant3 = 8'd191;
a_exp0 = 10'd615; a_exp1 = 10'd733; a_exp2 = 10'd480; a_exp3 = 10'd528;
b_exp0 = 10'd830; b_exp1 = 10'd583; b_exp2 = 10'd662; b_exp3 = 10'd835;
a_sign0 = 4'd2; a_sign1 = 4'd16; a_sign2 = 4'd5; a_sign3 = 4'd16;
b_sign0 = 4'd14; b_sign1 = 4'd16; b_sign2 = 4'd8; b_sign3 = 4'd6;
@(posedge clk_i);
a_mant0 = 8'd189; a_mant1 = 8'd222; a_mant2 = 8'd197; a_mant3 = 8'd99;
b_mant0 = 8'd109; b_mant1 = 8'd154; b_mant2 = 8'd174; b_mant3 = 8'd253;
a_exp0 = 10'd125; a_exp1 = 10'd753; a_exp2 = 10'd969; a_exp3 = 10'd267;
b_exp0 = 10'd841; b_exp1 = 10'd68; b_exp2 = 10'd480; b_exp3 = 10'd926;
a_sign0 = 4'd8; a_sign1 = 4'd12; a_sign2 = 4'd7; a_sign3 = 4'd13;
b_sign0 = 4'd11; b_sign1 = 4'd6; b_sign2 = 4'd6; b_sign3 = 4'd12;
@(posedge clk_i);
a_mant0 = 8'd17; a_mant1 = 8'd247; a_mant2 = 8'd191; a_mant3 = 8'd196;
b_mant0 = 8'd212; b_mant1 = 8'd151; b_mant2 = 8'd235; b_mant3 = 8'd27;
a_exp0 = 10'd970; a_exp1 = 10'd164; a_exp2 = 10'd870; a_exp3 = 10'd593;
b_exp0 = 10'd384; b_exp1 = 10'd208; b_exp2 = 10'd531; b_exp3 = 10'd360;
a_sign0 = 4'd1; a_sign1 = 4'd8; a_sign2 = 4'd12; a_sign3 = 4'd5;
b_sign0 = 4'd5; b_sign1 = 4'd4; b_sign2 = 4'd5; b_sign3 = 4'd8;
@(posedge clk_i);
a_mant0 = 8'd56; a_mant1 = 8'd218; a_mant2 = 8'd251; a_mant3 = 8'd133;
b_mant0 = 8'd181; b_mant1 = 8'd251; b_mant2 = 8'd80; b_mant3 = 8'd243;
a_exp0 = 10'd369; a_exp1 = 10'd158; a_exp2 = 10'd573; a_exp3 = 10'd155;
b_exp0 = 10'd699; b_exp1 = 10'd284; b_exp2 = 10'd530; b_exp3 = 10'd505;
a_sign0 = 4'd1; a_sign1 = 4'd2; a_sign2 = 4'd6; a_sign3 = 4'd5;
b_sign0 = 4'd15; b_sign1 = 4'd7; b_sign2 = 4'd9; b_sign3 = 4'd3;
@(posedge clk_i);
shared_exps0 = 8'd127;
shared_exps1 = 8'd123;
rstn = 0;
@(posedge clk_i);
rstn = 1;
a_mant0 = 8'd97; a_mant1 = 8'd237; a_mant2 = 8'd36; a_mant3 = 8'd235;
b_mant0 = 8'd128; b_mant1 = 8'd218; b_mant2 = 8'd110; b_mant3 = 8'd189;
a_exp0 = 10'd413; a_exp1 = 10'd998; a_exp2 = 10'd407; a_exp3 = 10'd37;
b_exp0 = 10'd77; b_exp1 = 10'd876; b_exp2 = 10'd949; b_exp3 = 10'd902;
a_sign0 = 4'd16; a_sign1 = 4'd1; a_sign2 = 4'd3; a_sign3 = 4'd14;
b_sign0 = 4'd12; b_sign1 = 4'd8; b_sign2 = 4'd9; b_sign3 = 4'd16;
@(posedge clk_i);
a_mant0 = 8'd85; a_mant1 = 8'd253; a_mant2 = 8'd197; a_mant3 = 8'd206;
b_mant0 = 8'd206; b_mant1 = 8'd71; b_mant2 = 8'd40; b_mant3 = 8'd89;
a_exp0 = 10'd631; a_exp1 = 10'd613; a_exp2 = 10'd76; a_exp3 = 10'd540;
b_exp0 = 10'd748; b_exp1 = 10'd756; b_exp2 = 10'd811; b_exp3 = 10'd377;
a_sign0 = 4'd5; a_sign1 = 4'd4; a_sign2 = 4'd10; a_sign3 = 4'd6;
b_sign0 = 4'd11; b_sign1 = 4'd14; b_sign2 = 4'd4; b_sign3 = 4'd2;
@(posedge clk_i);
a_mant0 = 8'd209; a_mant1 = 8'd213; a_mant2 = 8'd126; a_mant3 = 8'd156;
b_mant0 = 8'd63; b_mant1 = 8'd225; b_mant2 = 8'd26; b_mant3 = 8'd31;
a_exp0 = 10'd603; a_exp1 = 10'd626; a_exp2 = 10'd62; a_exp3 = 10'd216;
b_exp0 = 10'd948; b_exp1 = 10'd762; b_exp2 = 10'd954; b_exp3 = 10'd535;
a_sign0 = 4'd6; a_sign1 = 4'd14; a_sign2 = 4'd2; a_sign3 = 4'd2;
b_sign0 = 4'd5; b_sign1 = 4'd5; b_sign2 = 4'd1; b_sign3 = 4'd1;
@(posedge clk_i);
a_mant0 = 8'd137; a_mant1 = 8'd50; a_mant2 = 8'd88; a_mant3 = 8'd113;
b_mant0 = 8'd81; b_mant1 = 8'd104; b_mant2 = 8'd57; b_mant3 = 8'd201;
a_exp0 = 10'd907; a_exp1 = 10'd161; a_exp2 = 10'd720; a_exp3 = 10'd717;
b_exp0 = 10'd912; b_exp1 = 10'd766; b_exp2 = 10'd889; b_exp3 = 10'd306;
a_sign0 = 4'd16; a_sign1 = 4'd13; a_sign2 = 4'd3; a_sign3 = 4'd14;
b_sign0 = 4'd14; b_sign1 = 4'd2; b_sign2 = 4'd7; b_sign3 = 4'd12;
@(posedge clk_i);
a_mant0 = 8'd158; a_mant1 = 8'd142; a_mant2 = 8'd164; a_mant3 = 8'd66;
b_mant0 = 8'd26; b_mant1 = 8'd246; b_mant2 = 8'd220; b_mant3 = 8'd38;
a_exp0 = 10'd916; a_exp1 = 10'd868; a_exp2 = 10'd409; a_exp3 = 10'd392;
b_exp0 = 10'd515; b_exp1 = 10'd952; b_exp2 = 10'd688; b_exp3 = 10'd851;
a_sign0 = 4'd1; a_sign1 = 4'd6; a_sign2 = 4'd0; a_sign3 = 4'd6;
b_sign0 = 4'd0; b_sign1 = 4'd2; b_sign2 = 4'd5; b_sign3 = 4'd15;
@(posedge clk_i);
a_mant0 = 8'd5; a_mant1 = 8'd246; a_mant2 = 8'd87; a_mant3 = 8'd128;
b_mant0 = 8'd34; b_mant1 = 8'd25; b_mant2 = 8'd227; b_mant3 = 8'd224;
a_exp0 = 10'd584; a_exp1 = 10'd488; a_exp2 = 10'd788; a_exp3 = 10'd287;
b_exp0 = 10'd177; b_exp1 = 10'd368; b_exp2 = 10'd275; b_exp3 = 10'd818;
a_sign0 = 4'd3; a_sign1 = 4'd4; a_sign2 = 4'd8; a_sign3 = 4'd16;
b_sign0 = 4'd0; b_sign1 = 4'd11; b_sign2 = 4'd3; b_sign3 = 4'd3;
@(posedge clk_i);
a_mant0 = 8'd57; a_mant1 = 8'd10; a_mant2 = 8'd175; a_mant3 = 8'd241;
b_mant0 = 8'd98; b_mant1 = 8'd165; b_mant2 = 8'd184; b_mant3 = 8'd234;
a_exp0 = 10'd606; a_exp1 = 10'd316; a_exp2 = 10'd362; a_exp3 = 10'd835;
b_exp0 = 10'd426; b_exp1 = 10'd810; b_exp2 = 10'd755; b_exp3 = 10'd337;
a_sign0 = 4'd3; a_sign1 = 4'd15; a_sign2 = 4'd0; a_sign3 = 4'd0;
b_sign0 = 4'd13; b_sign1 = 4'd9; b_sign2 = 4'd11; b_sign3 = 4'd12;
@(posedge clk_i);
shared_exps0 = 8'd124;
shared_exps1 = 8'd113;
a_mant0 = 8'd23; a_mant1 = 8'd65; a_mant2 = 8'd60; a_mant3 = 8'd162;
b_mant0 = 8'd140; b_mant1 = 8'd118; b_mant2 = 8'd53; b_mant3 = 8'd43;
a_exp0 = 10'd840; a_exp1 = 10'd385; a_exp2 = 10'd428; a_exp3 = 10'd162;
b_exp0 = 10'd378; b_exp1 = 10'd847; b_exp2 = 10'd841; b_exp3 = 10'd420;
a_sign0 = 4'd5; a_sign1 = 4'd3; a_sign2 = 4'd4; a_sign3 = 4'd16;
b_sign0 = 4'd0; b_sign1 = 4'd8; b_sign2 = 4'd6; b_sign3 = 4'd4;
@(posedge clk_i);
a_mant0 = 8'd7; a_mant1 = 8'd6; a_mant2 = 8'd221; a_mant3 = 8'd242;
b_mant0 = 8'd148; b_mant1 = 8'd151; b_mant2 = 8'd12; b_mant3 = 8'd220;
a_exp0 = 10'd412; a_exp1 = 10'd438; a_exp2 = 10'd46; a_exp3 = 10'd858;
b_exp0 = 10'd340; b_exp1 = 10'd780; b_exp2 = 10'd766; b_exp3 = 10'd629;
a_sign0 = 4'd13; a_sign1 = 4'd4; a_sign2 = 4'd16; a_sign3 = 4'd8;
b_sign0 = 4'd11; b_sign1 = 4'd9; b_sign2 = 4'd11; b_sign3 = 4'd8;
@(posedge clk_i);
a_mant0 = 8'd138; a_mant1 = 8'd30; a_mant2 = 8'd60; a_mant3 = 8'd16;
b_mant0 = 8'd143; b_mant1 = 8'd14; b_mant2 = 8'd4; b_mant3 = 8'd217;
a_exp0 = 10'd518; a_exp1 = 10'd971; a_exp2 = 10'd721; a_exp3 = 10'd866;
b_exp0 = 10'd932; b_exp1 = 10'd263; b_exp2 = 10'd612; b_exp3 = 10'd299;
a_sign0 = 4'd15; a_sign1 = 4'd3; a_sign2 = 4'd5; a_sign3 = 4'd0;
b_sign0 = 4'd7; b_sign1 = 4'd1; b_sign2 = 4'd5; b_sign3 = 4'd13;
@(posedge clk_i);
a_mant0 = 8'd201; a_mant1 = 8'd156; a_mant2 = 8'd235; a_mant3 = 8'd33;
b_mant0 = 8'd229; b_mant1 = 8'd2; b_mant2 = 8'd3; b_mant3 = 8'd125;
a_exp0 = 10'd959; a_exp1 = 10'd162; a_exp2 = 10'd886; a_exp3 = 10'd580;
b_exp0 = 10'd6; b_exp1 = 10'd848; b_exp2 = 10'd428; b_exp3 = 10'd278;
a_sign0 = 4'd13; a_sign1 = 4'd15; a_sign2 = 4'd2; a_sign3 = 4'd3;
b_sign0 = 4'd7; b_sign1 = 4'd14; b_sign2 = 4'd6; b_sign3 = 4'd13;
@(posedge clk_i);
a_mant0 = 8'd236; a_mant1 = 8'd32; a_mant2 = 8'd109; a_mant3 = 8'd9;
b_mant0 = 8'd105; b_mant1 = 8'd237; b_mant2 = 8'd251; b_mant3 = 8'd192;
a_exp0 = 10'd839; a_exp1 = 10'd806; a_exp2 = 10'd450; a_exp3 = 10'd23;
b_exp0 = 10'd554; b_exp1 = 10'd541; b_exp2 = 10'd194; b_exp3 = 10'd462;
a_sign0 = 4'd7; a_sign1 = 4'd14; a_sign2 = 4'd12; a_sign3 = 4'd10;
b_sign0 = 4'd1; b_sign1 = 4'd0; b_sign2 = 4'd11; b_sign3 = 4'd9;
@(posedge clk_i);
a_mant0 = 8'd172; a_mant1 = 8'd203; a_mant2 = 8'd65; a_mant3 = 8'd154;
b_mant0 = 8'd100; b_mant1 = 8'd144; b_mant2 = 8'd122; b_mant3 = 8'd134;
a_exp0 = 10'd87; a_exp1 = 10'd702; a_exp2 = 10'd220; a_exp3 = 10'd403;
b_exp0 = 10'd618; b_exp1 = 10'd337; b_exp2 = 10'd64; b_exp3 = 10'd936;
a_sign0 = 4'd6; a_sign1 = 4'd12; a_sign2 = 4'd13; a_sign3 = 4'd9;
b_sign0 = 4'd11; b_sign1 = 4'd11; b_sign2 = 4'd9; b_sign3 = 4'd0;
@(posedge clk_i);
a_mant0 = 8'd4; a_mant1 = 8'd47; a_mant2 = 8'd4; a_mant3 = 8'd100;
b_mant0 = 8'd106; b_mant1 = 8'd235; b_mant2 = 8'd162; b_mant3 = 8'd169;
a_exp0 = 10'd713; a_exp1 = 10'd215; a_exp2 = 10'd45; a_exp3 = 10'd509;
b_exp0 = 10'd356; b_exp1 = 10'd295; b_exp2 = 10'd1008; b_exp3 = 10'd573;
a_sign0 = 4'd6; a_sign1 = 4'd14; a_sign2 = 4'd5; a_sign3 = 4'd16;
b_sign0 = 4'd1; b_sign1 = 4'd8; b_sign2 = 4'd2; b_sign3 = 4'd1;
@(posedge clk_i);
a_mant0 = 8'd223; a_mant1 = 8'd85; a_mant2 = 8'd183; a_mant3 = 8'd79;
b_mant0 = 8'd7; b_mant1 = 8'd74; b_mant2 = 8'd130; b_mant3 = 8'd228;
a_exp0 = 10'd411; a_exp1 = 10'd195; a_exp2 = 10'd413; a_exp3 = 10'd964;
b_exp0 = 10'd909; b_exp1 = 10'd641; b_exp2 = 10'd948; b_exp3 = 10'd939;
a_sign0 = 4'd10; a_sign1 = 4'd5; a_sign2 = 4'd12; a_sign3 = 4'd11;
b_sign0 = 4'd10; b_sign1 = 4'd5; b_sign2 = 4'd3; b_sign3 = 4'd11;
@(posedge clk_i);
shared_exps0 = 8'd122;
shared_exps1 = 8'd116;
a_mant0 = 8'd99; a_mant1 = 8'd168; a_mant2 = 8'd40; a_mant3 = 8'd231;
b_mant0 = 8'd47; b_mant1 = 8'd17; b_mant2 = 8'd39; b_mant3 = 8'd72;
a_exp0 = 10'd760; a_exp1 = 10'd218; a_exp2 = 10'd980; a_exp3 = 10'd171;
b_exp0 = 10'd574; b_exp1 = 10'd245; b_exp2 = 10'd145; b_exp3 = 10'd537;
a_sign0 = 4'd7; a_sign1 = 4'd3; a_sign2 = 4'd9; a_sign3 = 4'd8;
b_sign0 = 4'd2; b_sign1 = 4'd2; b_sign2 = 4'd4; b_sign3 = 4'd3;
@(posedge clk_i);
a_mant0 = 8'd46; a_mant1 = 8'd63; a_mant2 = 8'd60; a_mant3 = 8'd172;
b_mant0 = 8'd77; b_mant1 = 8'd11; b_mant2 = 8'd51; b_mant3 = 8'd198;
a_exp0 = 10'd918; a_exp1 = 10'd965; a_exp2 = 10'd569; a_exp3 = 10'd245;
b_exp0 = 10'd726; b_exp1 = 10'd707; b_exp2 = 10'd778; b_exp3 = 10'd628;
a_sign0 = 4'd8; a_sign1 = 4'd3; a_sign2 = 4'd4; a_sign3 = 4'd16;
b_sign0 = 4'd2; b_sign1 = 4'd9; b_sign2 = 4'd0; b_sign3 = 4'd16;
@(posedge clk_i);
a_mant0 = 8'd37; a_mant1 = 8'd44; a_mant2 = 8'd41; a_mant3 = 8'd175;
b_mant0 = 8'd223; b_mant1 = 8'd84; b_mant2 = 8'd170; b_mant3 = 8'd248;
a_exp0 = 10'd367; a_exp1 = 10'd269; a_exp2 = 10'd748; a_exp3 = 10'd442;
b_exp0 = 10'd785; b_exp1 = 10'd859; b_exp2 = 10'd155; b_exp3 = 10'd378;
a_sign0 = 4'd16; a_sign1 = 4'd13; a_sign2 = 4'd8; a_sign3 = 4'd4;
b_sign0 = 4'd4; b_sign1 = 4'd8; b_sign2 = 4'd14; b_sign3 = 4'd16;
@(posedge clk_i);
a_mant0 = 8'd176; a_mant1 = 8'd46; a_mant2 = 8'd209; a_mant3 = 8'd223;
b_mant0 = 8'd54; b_mant1 = 8'd41; b_mant2 = 8'd101; b_mant3 = 8'd46;
a_exp0 = 10'd594; a_exp1 = 10'd336; a_exp2 = 10'd568; a_exp3 = 10'd466;
b_exp0 = 10'd508; b_exp1 = 10'd840; b_exp2 = 10'd942; b_exp3 = 10'd60;
a_sign0 = 4'd16; a_sign1 = 4'd1; a_sign2 = 4'd5; a_sign3 = 4'd2;
b_sign0 = 4'd2; b_sign1 = 4'd4; b_sign2 = 4'd4; b_sign3 = 4'd5;
@(posedge clk_i);
a_mant0 = 8'd54; a_mant1 = 8'd20; a_mant2 = 8'd135; a_mant3 = 8'd208;
b_mant0 = 8'd178; b_mant1 = 8'd24; b_mant2 = 8'd218; b_mant3 = 8'd10;
a_exp0 = 10'd820; a_exp1 = 10'd457; a_exp2 = 10'd564; a_exp3 = 10'd146;
b_exp0 = 10'd84; b_exp1 = 10'd59; b_exp2 = 10'd312; b_exp3 = 10'd549;
a_sign0 = 4'd4; a_sign1 = 4'd9; a_sign2 = 4'd9; a_sign3 = 4'd0;
b_sign0 = 4'd13; b_sign1 = 4'd12; b_sign2 = 4'd7; b_sign3 = 4'd6;
@(posedge clk_i);
a_mant0 = 8'd77; a_mant1 = 8'd166; a_mant2 = 8'd14; a_mant3 = 8'd217;
b_mant0 = 8'd165; b_mant1 = 8'd128; b_mant2 = 8'd196; b_mant3 = 8'd84;
a_exp0 = 10'd419; a_exp1 = 10'd349; a_exp2 = 10'd562; a_exp3 = 10'd516;
b_exp0 = 10'd24; b_exp1 = 10'd310; b_exp2 = 10'd938; b_exp3 = 10'd42;
a_sign0 = 4'd16; a_sign1 = 4'd14; a_sign2 = 4'd9; a_sign3 = 4'd1;
b_sign0 = 4'd10; b_sign1 = 4'd10; b_sign2 = 4'd6; b_sign3 = 4'd1;
@(posedge clk_i);
a_mant0 = 8'd134; a_mant1 = 8'd69; a_mant2 = 8'd110; a_mant3 = 8'd140;
b_mant0 = 8'd17; b_mant1 = 8'd174; b_mant2 = 8'd86; b_mant3 = 8'd32;
a_exp0 = 10'd548; a_exp1 = 10'd652; a_exp2 = 10'd811; a_exp3 = 10'd338;
b_exp0 = 10'd964; b_exp1 = 10'd857; b_exp2 = 10'd91; b_exp3 = 10'd140;
a_sign0 = 4'd14; a_sign1 = 4'd16; a_sign2 = 4'd6; a_sign3 = 4'd13;
b_sign0 = 4'd11; b_sign1 = 4'd11; b_sign2 = 4'd13; b_sign3 = 4'd9;
@(posedge clk_i);
a_mant0 = 8'd21; a_mant1 = 8'd91; a_mant2 = 8'd15; a_mant3 = 8'd119;
b_mant0 = 8'd152; b_mant1 = 8'd145; b_mant2 = 8'd116; b_mant3 = 8'd1;
a_exp0 = 10'd813; a_exp1 = 10'd731; a_exp2 = 10'd353; a_exp3 = 10'd873;
b_exp0 = 10'd621; b_exp1 = 10'd642; b_exp2 = 10'd293; b_exp3 = 10'd142;
a_sign0 = 4'd6; a_sign1 = 4'd7; a_sign2 = 4'd10; a_sign3 = 4'd0;
b_sign0 = 4'd0; b_sign1 = 4'd14; b_sign2 = 4'd15; b_sign3 = 4'd9;
@(posedge clk_i);
shared_exps0 = 8'd128;
shared_exps1 = 8'd114;
a_mant0 = 8'd93; a_mant1 = 8'd179; a_mant2 = 8'd189; a_mant3 = 8'd95;
b_mant0 = 8'd176; b_mant1 = 8'd34; b_mant2 = 8'd118; b_mant3 = 8'd77;
a_exp0 = 10'd936; a_exp1 = 10'd1000; a_exp2 = 10'd595; a_exp3 = 10'd253;
b_exp0 = 10'd4; b_exp1 = 10'd535; b_exp2 = 10'd328; b_exp3 = 10'd73;
a_sign0 = 4'd3; a_sign1 = 4'd12; a_sign2 = 4'd9; a_sign3 = 4'd5;
b_sign0 = 4'd15; b_sign1 = 4'd9; b_sign2 = 4'd14; b_sign3 = 4'd0;
@(posedge clk_i);
a_mant0 = 8'd127; a_mant1 = 8'd223; a_mant2 = 8'd1; a_mant3 = 8'd206;
b_mant0 = 8'd79; b_mant1 = 8'd32; b_mant2 = 8'd238; b_mant3 = 8'd95;
a_exp0 = 10'd738; a_exp1 = 10'd617; a_exp2 = 10'd273; a_exp3 = 10'd253;
b_exp0 = 10'd222; b_exp1 = 10'd79; b_exp2 = 10'd312; b_exp3 = 10'd539;
a_sign0 = 4'd8; a_sign1 = 4'd3; a_sign2 = 4'd13; a_sign3 = 4'd1;
b_sign0 = 4'd0; b_sign1 = 4'd12; b_sign2 = 4'd3; b_sign3 = 4'd10;
@(posedge clk_i);
a_mant0 = 8'd130; a_mant1 = 8'd240; a_mant2 = 8'd173; a_mant3 = 8'd161;
b_mant0 = 8'd254; b_mant1 = 8'd254; b_mant2 = 8'd154; b_mant3 = 8'd252;
a_exp0 = 10'd713; a_exp1 = 10'd809; a_exp2 = 10'd760; a_exp3 = 10'd443;
b_exp0 = 10'd555; b_exp1 = 10'd680; b_exp2 = 10'd438; b_exp3 = 10'd146;
a_sign0 = 4'd9; a_sign1 = 4'd16; a_sign2 = 4'd10; a_sign3 = 4'd0;
b_sign0 = 4'd7; b_sign1 = 4'd11; b_sign2 = 4'd15; b_sign3 = 4'd16;
@(posedge clk_i);
a_mant0 = 8'd141; a_mant1 = 8'd223; a_mant2 = 8'd76; a_mant3 = 8'd131;
b_mant0 = 8'd23; b_mant1 = 8'd70; b_mant2 = 8'd250; b_mant3 = 8'd49;
a_exp0 = 10'd514; a_exp1 = 10'd966; a_exp2 = 10'd159; a_exp3 = 10'd199;
b_exp0 = 10'd459; b_exp1 = 10'd602; b_exp2 = 10'd141; b_exp3 = 10'd525;
a_sign0 = 4'd16; a_sign1 = 4'd5; a_sign2 = 4'd15; a_sign3 = 4'd9;
b_sign0 = 4'd2; b_sign1 = 4'd11; b_sign2 = 4'd7; b_sign3 = 4'd14;
@(posedge clk_i);
a_mant0 = 8'd223; a_mant1 = 8'd12; a_mant2 = 8'd170; a_mant3 = 8'd96;
b_mant0 = 8'd244; b_mant1 = 8'd215; b_mant2 = 8'd81; b_mant3 = 8'd95;
a_exp0 = 10'd177; a_exp1 = 10'd552; a_exp2 = 10'd12; a_exp3 = 10'd699;
b_exp0 = 10'd437; b_exp1 = 10'd416; b_exp2 = 10'd958; b_exp3 = 10'd408;
a_sign0 = 4'd4; a_sign1 = 4'd13; a_sign2 = 4'd16; a_sign3 = 4'd5;
b_sign0 = 4'd16; b_sign1 = 4'd8; b_sign2 = 4'd7; b_sign3 = 4'd8;
@(posedge clk_i);
a_mant0 = 8'd242; a_mant1 = 8'd9; a_mant2 = 8'd206; a_mant3 = 8'd62;
b_mant0 = 8'd102; b_mant1 = 8'd240; b_mant2 = 8'd16; b_mant3 = 8'd60;
a_exp0 = 10'd278; a_exp1 = 10'd195; a_exp2 = 10'd185; a_exp3 = 10'd884;
b_exp0 = 10'd396; b_exp1 = 10'd1008; b_exp2 = 10'd363; b_exp3 = 10'd83;
a_sign0 = 4'd4; a_sign1 = 4'd14; a_sign2 = 4'd5; a_sign3 = 4'd3;
b_sign0 = 4'd9; b_sign1 = 4'd12; b_sign2 = 4'd3; b_sign3 = 4'd14;
@(posedge clk_i);
a_mant0 = 8'd124; a_mant1 = 8'd201; a_mant2 = 8'd185; a_mant3 = 8'd149;
b_mant0 = 8'd194; b_mant1 = 8'd129; b_mant2 = 8'd103; b_mant3 = 8'd19;
a_exp0 = 10'd181; a_exp1 = 10'd939; a_exp2 = 10'd446; a_exp3 = 10'd687;
b_exp0 = 10'd56; b_exp1 = 10'd372; b_exp2 = 10'd961; b_exp3 = 10'd614;
a_sign0 = 4'd8; a_sign1 = 4'd10; a_sign2 = 4'd8; a_sign3 = 4'd5;
b_sign0 = 4'd3; b_sign1 = 4'd12; b_sign2 = 4'd3; b_sign3 = 4'd15;
@(posedge clk_i);
a_mant0 = 8'd218; a_mant1 = 8'd151; a_mant2 = 8'd163; a_mant3 = 8'd30;
b_mant0 = 8'd77; b_mant1 = 8'd151; b_mant2 = 8'd8; b_mant3 = 8'd59;
a_exp0 = 10'd929; a_exp1 = 10'd604; a_exp2 = 10'd98; a_exp3 = 10'd517;
b_exp0 = 10'd335; b_exp1 = 10'd648; b_exp2 = 10'd425; b_exp3 = 10'd705;
a_sign0 = 4'd6; a_sign1 = 4'd10; a_sign2 = 4'd16; a_sign3 = 4'd16;
b_sign0 = 4'd9; b_sign1 = 4'd0; b_sign2 = 4'd14; b_sign3 = 4'd8;
@(posedge clk_i);
shared_exps0 = 8'd162;
shared_exps1 = 8'd97;
rstn = 0;
@(posedge clk_i);
rstn = 1;
a_mant0 = 8'd82; a_mant1 = 8'd202; a_mant2 = 8'd95; a_mant3 = 8'd7;
b_mant0 = 8'd180; b_mant1 = 8'd110; b_mant2 = 8'd78; b_mant3 = 8'd241;
a_exp0 = 10'd506; a_exp1 = 10'd810; a_exp2 = 10'd973; a_exp3 = 10'd852;
b_exp0 = 10'd183; b_exp1 = 10'd335; b_exp2 = 10'd113; b_exp3 = 10'd256;
a_sign0 = 4'd15; a_sign1 = 4'd5; a_sign2 = 4'd5; a_sign3 = 4'd2;
b_sign0 = 4'd16; b_sign1 = 4'd12; b_sign2 = 4'd10; b_sign3 = 4'd7;
@(posedge clk_i);
a_mant0 = 8'd224; a_mant1 = 8'd50; a_mant2 = 8'd206; a_mant3 = 8'd23;
b_mant0 = 8'd89; b_mant1 = 8'd89; b_mant2 = 8'd115; b_mant3 = 8'd196;
a_exp0 = 10'd572; a_exp1 = 10'd89; a_exp2 = 10'd698; a_exp3 = 10'd409;
b_exp0 = 10'd105; b_exp1 = 10'd525; b_exp2 = 10'd1014; b_exp3 = 10'd289;
a_sign0 = 4'd5; a_sign1 = 4'd12; a_sign2 = 4'd16; a_sign3 = 4'd3;
b_sign0 = 4'd14; b_sign1 = 4'd11; b_sign2 = 4'd13; b_sign3 = 4'd14;
@(posedge clk_i);
a_mant0 = 8'd10; a_mant1 = 8'd8; a_mant2 = 8'd105; a_mant3 = 8'd136;
b_mant0 = 8'd87; b_mant1 = 8'd177; b_mant2 = 8'd138; b_mant3 = 8'd102;
a_exp0 = 10'd8; a_exp1 = 10'd639; a_exp2 = 10'd521; a_exp3 = 10'd35;
b_exp0 = 10'd552; b_exp1 = 10'd983; b_exp2 = 10'd420; b_exp3 = 10'd586;
a_sign0 = 4'd3; a_sign1 = 4'd1; a_sign2 = 4'd10; a_sign3 = 4'd11;
b_sign0 = 4'd9; b_sign1 = 4'd10; b_sign2 = 4'd4; b_sign3 = 4'd13;
@(posedge clk_i);
a_mant0 = 8'd86; a_mant1 = 8'd26; a_mant2 = 8'd125; a_mant3 = 8'd87;
b_mant0 = 8'd136; b_mant1 = 8'd191; b_mant2 = 8'd44; b_mant3 = 8'd20;
a_exp0 = 10'd884; a_exp1 = 10'd543; a_exp2 = 10'd267; a_exp3 = 10'd64;
b_exp0 = 10'd644; b_exp1 = 10'd577; b_exp2 = 10'd669; b_exp3 = 10'd667;
a_sign0 = 4'd8; a_sign1 = 4'd11; a_sign2 = 4'd2; a_sign3 = 4'd9;
b_sign0 = 4'd4; b_sign1 = 4'd16; b_sign2 = 4'd6; b_sign3 = 4'd15;
@(posedge clk_i);
a_mant0 = 8'd45; a_mant1 = 8'd116; a_mant2 = 8'd57; a_mant3 = 8'd147;
b_mant0 = 8'd9; b_mant1 = 8'd16; b_mant2 = 8'd241; b_mant3 = 8'd36;
a_exp0 = 10'd923; a_exp1 = 10'd519; a_exp2 = 10'd267; a_exp3 = 10'd186;
b_exp0 = 10'd435; b_exp1 = 10'd267; b_exp2 = 10'd790; b_exp3 = 10'd216;
a_sign0 = 4'd12; a_sign1 = 4'd3; a_sign2 = 4'd2; a_sign3 = 4'd0;
b_sign0 = 4'd4; b_sign1 = 4'd10; b_sign2 = 4'd7; b_sign3 = 4'd0;
@(posedge clk_i);
a_mant0 = 8'd237; a_mant1 = 8'd205; a_mant2 = 8'd172; a_mant3 = 8'd186;
b_mant0 = 8'd57; b_mant1 = 8'd139; b_mant2 = 8'd202; b_mant3 = 8'd75;
a_exp0 = 10'd770; a_exp1 = 10'd760; a_exp2 = 10'd758; a_exp3 = 10'd693;
b_exp0 = 10'd918; b_exp1 = 10'd315; b_exp2 = 10'd313; b_exp3 = 10'd597;
a_sign0 = 4'd5; a_sign1 = 4'd15; a_sign2 = 4'd8; a_sign3 = 4'd6;
b_sign0 = 4'd9; b_sign1 = 4'd4; b_sign2 = 4'd8; b_sign3 = 4'd16;
@(posedge clk_i);
a_mant0 = 8'd212; a_mant1 = 8'd77; a_mant2 = 8'd61; a_mant3 = 8'd70;
b_mant0 = 8'd59; b_mant1 = 8'd0; b_mant2 = 8'd79; b_mant3 = 8'd62;
a_exp0 = 10'd488; a_exp1 = 10'd55; a_exp2 = 10'd981; a_exp3 = 10'd260;
b_exp0 = 10'd484; b_exp1 = 10'd677; b_exp2 = 10'd746; b_exp3 = 10'd561;
a_sign0 = 4'd9; a_sign1 = 4'd5; a_sign2 = 4'd15; a_sign3 = 4'd15;
b_sign0 = 4'd0; b_sign1 = 4'd1; b_sign2 = 4'd0; b_sign3 = 4'd15;
@(posedge clk_i);
shared_exps0 = 8'd132;
shared_exps1 = 8'd119;
a_mant0 = 8'd36; a_mant1 = 8'd131; a_mant2 = 8'd146; a_mant3 = 8'd156;
b_mant0 = 8'd196; b_mant1 = 8'd100; b_mant2 = 8'd173; b_mant3 = 8'd183;
a_exp0 = 10'd972; a_exp1 = 10'd182; a_exp2 = 10'd104; a_exp3 = 10'd685;
b_exp0 = 10'd271; b_exp1 = 10'd17; b_exp2 = 10'd600; b_exp3 = 10'd217;
a_sign0 = 4'd15; a_sign1 = 4'd10; a_sign2 = 4'd11; a_sign3 = 4'd16;
b_sign0 = 4'd11; b_sign1 = 4'd9; b_sign2 = 4'd3; b_sign3 = 4'd2;
@(posedge clk_i);
a_mant0 = 8'd210; a_mant1 = 8'd164; a_mant2 = 8'd202; a_mant3 = 8'd189;
b_mant0 = 8'd49; b_mant1 = 8'd240; b_mant2 = 8'd201; b_mant3 = 8'd67;
a_exp0 = 10'd531; a_exp1 = 10'd109; a_exp2 = 10'd320; a_exp3 = 10'd883;
b_exp0 = 10'd845; b_exp1 = 10'd48; b_exp2 = 10'd248; b_exp3 = 10'd999;
a_sign0 = 4'd1; a_sign1 = 4'd14; a_sign2 = 4'd7; a_sign3 = 4'd16;
b_sign0 = 4'd12; b_sign1 = 4'd2; b_sign2 = 4'd10; b_sign3 = 4'd0;
@(posedge clk_i);
a_mant0 = 8'd98; a_mant1 = 8'd25; a_mant2 = 8'd180; a_mant3 = 8'd133;
b_mant0 = 8'd89; b_mant1 = 8'd241; b_mant2 = 8'd29; b_mant3 = 8'd71;
a_exp0 = 10'd329; a_exp1 = 10'd703; a_exp2 = 10'd37; a_exp3 = 10'd881;
b_exp0 = 10'd1003; b_exp1 = 10'd454; b_exp2 = 10'd115; b_exp3 = 10'd341;
a_sign0 = 4'd4; a_sign1 = 4'd10; a_sign2 = 4'd9; a_sign3 = 4'd2;
b_sign0 = 4'd11; b_sign1 = 4'd13; b_sign2 = 4'd5; b_sign3 = 4'd15;
@(posedge clk_i);
a_mant0 = 8'd85; a_mant1 = 8'd172; a_mant2 = 8'd2; a_mant3 = 8'd15;
b_mant0 = 8'd235; b_mant1 = 8'd221; b_mant2 = 8'd39; b_mant3 = 8'd67;
a_exp0 = 10'd803; a_exp1 = 10'd635; a_exp2 = 10'd800; a_exp3 = 10'd685;
b_exp0 = 10'd811; b_exp1 = 10'd671; b_exp2 = 10'd977; b_exp3 = 10'd447;
a_sign0 = 4'd5; a_sign1 = 4'd2; a_sign2 = 4'd10; a_sign3 = 4'd2;
b_sign0 = 4'd12; b_sign1 = 4'd2; b_sign2 = 4'd8; b_sign3 = 4'd3;
@(posedge clk_i);
a_mant0 = 8'd236; a_mant1 = 8'd197; a_mant2 = 8'd236; a_mant3 = 8'd64;
b_mant0 = 8'd141; b_mant1 = 8'd28; b_mant2 = 8'd157; b_mant3 = 8'd40;
a_exp0 = 10'd1008; a_exp1 = 10'd410; a_exp2 = 10'd287; a_exp3 = 10'd104;
b_exp0 = 10'd251; b_exp1 = 10'd122; b_exp2 = 10'd359; b_exp3 = 10'd762;
a_sign0 = 4'd5; a_sign1 = 4'd11; a_sign2 = 4'd15; a_sign3 = 4'd9;
b_sign0 = 4'd13; b_sign1 = 4'd15; b_sign2 = 4'd4; b_sign3 = 4'd9;
@(posedge clk_i);
a_mant0 = 8'd124; a_mant1 = 8'd244; a_mant2 = 8'd7; a_mant3 = 8'd214;
b_mant0 = 8'd190; b_mant1 = 8'd106; b_mant2 = 8'd28; b_mant3 = 8'd15;
a_exp0 = 10'd687; a_exp1 = 10'd996; a_exp2 = 10'd142; a_exp3 = 10'd500;
b_exp0 = 10'd16; b_exp1 = 10'd377; b_exp2 = 10'd888; b_exp3 = 10'd88;
a_sign0 = 4'd6; a_sign1 = 4'd7; a_sign2 = 4'd0; a_sign3 = 4'd7;
b_sign0 = 4'd13; b_sign1 = 4'd16; b_sign2 = 4'd11; b_sign3 = 4'd13;
@(posedge clk_i);
a_mant0 = 8'd86; a_mant1 = 8'd140; a_mant2 = 8'd61; a_mant3 = 8'd45;
b_mant0 = 8'd175; b_mant1 = 8'd114; b_mant2 = 8'd74; b_mant3 = 8'd27;
a_exp0 = 10'd98; a_exp1 = 10'd919; a_exp2 = 10'd11; a_exp3 = 10'd445;
b_exp0 = 10'd753; b_exp1 = 10'd1021; b_exp2 = 10'd404; b_exp3 = 10'd511;
a_sign0 = 4'd16; a_sign1 = 4'd14; a_sign2 = 4'd15; a_sign3 = 4'd15;
b_sign0 = 4'd10; b_sign1 = 4'd7; b_sign2 = 4'd16; b_sign3 = 4'd11;
@(posedge clk_i);
a_mant0 = 8'd20; a_mant1 = 8'd176; a_mant2 = 8'd173; a_mant3 = 8'd173;
b_mant0 = 8'd21; b_mant1 = 8'd104; b_mant2 = 8'd66; b_mant3 = 8'd236;
a_exp0 = 10'd122; a_exp1 = 10'd120; a_exp2 = 10'd98; a_exp3 = 10'd740;
b_exp0 = 10'd941; b_exp1 = 10'd370; b_exp2 = 10'd413; b_exp3 = 10'd580;
a_sign0 = 4'd15; a_sign1 = 4'd11; a_sign2 = 4'd0; a_sign3 = 4'd14;
b_sign0 = 4'd4; b_sign1 = 4'd4; b_sign2 = 4'd8; b_sign3 = 4'd9;
@(posedge clk_i);
shared_exps0 = 8'd141;
shared_exps1 = 8'd136;
a_mant0 = 8'd35; a_mant1 = 8'd208; a_mant2 = 8'd91; a_mant3 = 8'd149;
b_mant0 = 8'd52; b_mant1 = 8'd75; b_mant2 = 8'd160; b_mant3 = 8'd59;
a_exp0 = 10'd40; a_exp1 = 10'd202; a_exp2 = 10'd501; a_exp3 = 10'd211;
b_exp0 = 10'd263; b_exp1 = 10'd988; b_exp2 = 10'd855; b_exp3 = 10'd693;
a_sign0 = 4'd2; a_sign1 = 4'd0; a_sign2 = 4'd1; a_sign3 = 4'd16;
b_sign0 = 4'd1; b_sign1 = 4'd1; b_sign2 = 4'd6; b_sign3 = 4'd10;
@(posedge clk_i);
a_mant0 = 8'd219; a_mant1 = 8'd65; a_mant2 = 8'd121; a_mant3 = 8'd255;
b_mant0 = 8'd126; b_mant1 = 8'd79; b_mant2 = 8'd184; b_mant3 = 8'd48;
a_exp0 = 10'd641; a_exp1 = 10'd682; a_exp2 = 10'd884; a_exp3 = 10'd273;
b_exp0 = 10'd87; b_exp1 = 10'd714; b_exp2 = 10'd72; b_exp3 = 10'd910;
a_sign0 = 4'd16; a_sign1 = 4'd10; a_sign2 = 4'd15; a_sign3 = 4'd3;
b_sign0 = 4'd0; b_sign1 = 4'd11; b_sign2 = 4'd8; b_sign3 = 4'd5;
@(posedge clk_i);
a_mant0 = 8'd40; a_mant1 = 8'd209; a_mant2 = 8'd14; a_mant3 = 8'd31;
b_mant0 = 8'd103; b_mant1 = 8'd228; b_mant2 = 8'd243; b_mant3 = 8'd253;
a_exp0 = 10'd915; a_exp1 = 10'd491; a_exp2 = 10'd959; a_exp3 = 10'd109;
b_exp0 = 10'd934; b_exp1 = 10'd980; b_exp2 = 10'd412; b_exp3 = 10'd661;
a_sign0 = 4'd7; a_sign1 = 4'd3; a_sign2 = 4'd12; a_sign3 = 4'd0;
b_sign0 = 4'd15; b_sign1 = 4'd10; b_sign2 = 4'd1; b_sign3 = 4'd2;
@(posedge clk_i);
a_mant0 = 8'd217; a_mant1 = 8'd142; a_mant2 = 8'd188; a_mant3 = 8'd239;
b_mant0 = 8'd191; b_mant1 = 8'd134; b_mant2 = 8'd154; b_mant3 = 8'd89;
a_exp0 = 10'd1004; a_exp1 = 10'd363; a_exp2 = 10'd710; a_exp3 = 10'd651;
b_exp0 = 10'd678; b_exp1 = 10'd802; b_exp2 = 10'd200; b_exp3 = 10'd193;
a_sign0 = 4'd14; a_sign1 = 4'd10; a_sign2 = 4'd16; a_sign3 = 4'd6;
b_sign0 = 4'd4; b_sign1 = 4'd1; b_sign2 = 4'd1; b_sign3 = 4'd5;
@(posedge clk_i);
a_mant0 = 8'd103; a_mant1 = 8'd244; a_mant2 = 8'd22; a_mant3 = 8'd166;
b_mant0 = 8'd209; b_mant1 = 8'd222; b_mant2 = 8'd33; b_mant3 = 8'd88;
a_exp0 = 10'd374; a_exp1 = 10'd134; a_exp2 = 10'd190; a_exp3 = 10'd453;
b_exp0 = 10'd375; b_exp1 = 10'd464; b_exp2 = 10'd433; b_exp3 = 10'd536;
a_sign0 = 4'd4; a_sign1 = 4'd13; a_sign2 = 4'd8; a_sign3 = 4'd12;
b_sign0 = 4'd5; b_sign1 = 4'd11; b_sign2 = 4'd11; b_sign3 = 4'd12;
@(posedge clk_i);
a_mant0 = 8'd176; a_mant1 = 8'd149; a_mant2 = 8'd255; a_mant3 = 8'd236;
b_mant0 = 8'd249; b_mant1 = 8'd90; b_mant2 = 8'd16; b_mant3 = 8'd137;
a_exp0 = 10'd49; a_exp1 = 10'd67; a_exp2 = 10'd370; a_exp3 = 10'd392;
b_exp0 = 10'd967; b_exp1 = 10'd472; b_exp2 = 10'd250; b_exp3 = 10'd746;
a_sign0 = 4'd3; a_sign1 = 4'd7; a_sign2 = 4'd2; a_sign3 = 4'd8;
b_sign0 = 4'd6; b_sign1 = 4'd10; b_sign2 = 4'd1; b_sign3 = 4'd16;
@(posedge clk_i);
a_mant0 = 8'd156; a_mant1 = 8'd226; a_mant2 = 8'd85; a_mant3 = 8'd9;
b_mant0 = 8'd46; b_mant1 = 8'd246; b_mant2 = 8'd44; b_mant3 = 8'd152;
a_exp0 = 10'd663; a_exp1 = 10'd288; a_exp2 = 10'd391; a_exp3 = 10'd76;
b_exp0 = 10'd258; b_exp1 = 10'd110; b_exp2 = 10'd848; b_exp3 = 10'd640;
a_sign0 = 4'd6; a_sign1 = 4'd10; a_sign2 = 4'd15; a_sign3 = 4'd3;
b_sign0 = 4'd11; b_sign1 = 4'd11; b_sign2 = 4'd13; b_sign3 = 4'd7;
@(posedge clk_i);
a_mant0 = 8'd39; a_mant1 = 8'd227; a_mant2 = 8'd227; a_mant3 = 8'd18;
b_mant0 = 8'd67; b_mant1 = 8'd95; b_mant2 = 8'd75; b_mant3 = 8'd187;
a_exp0 = 10'd758; a_exp1 = 10'd230; a_exp2 = 10'd959; a_exp3 = 10'd949;
b_exp0 = 10'd325; b_exp1 = 10'd874; b_exp2 = 10'd901; b_exp3 = 10'd1;
a_sign0 = 4'd1; a_sign1 = 4'd2; a_sign2 = 4'd1; a_sign3 = 4'd7;
b_sign0 = 4'd6; b_sign1 = 4'd14; b_sign2 = 4'd4; b_sign3 = 4'd5;
@(posedge clk_i);
shared_exps0 = 8'd146;
shared_exps1 = 8'd102;
a_mant0 = 8'd157; a_mant1 = 8'd226; a_mant2 = 8'd111; a_mant3 = 8'd116;
b_mant0 = 8'd38; b_mant1 = 8'd90; b_mant2 = 8'd198; b_mant3 = 8'd128;
a_exp0 = 10'd416; a_exp1 = 10'd111; a_exp2 = 10'd913; a_exp3 = 10'd409;
b_exp0 = 10'd610; b_exp1 = 10'd505; b_exp2 = 10'd456; b_exp3 = 10'd913;
a_sign0 = 4'd16; a_sign1 = 4'd9; a_sign2 = 4'd0; a_sign3 = 4'd4;
b_sign0 = 4'd7; b_sign1 = 4'd0; b_sign2 = 4'd16; b_sign3 = 4'd9;
@(posedge clk_i);
a_mant0 = 8'd126; a_mant1 = 8'd171; a_mant2 = 8'd226; a_mant3 = 8'd193;
b_mant0 = 8'd228; b_mant1 = 8'd40; b_mant2 = 8'd217; b_mant3 = 8'd80;
a_exp0 = 10'd620; a_exp1 = 10'd653; a_exp2 = 10'd757; a_exp3 = 10'd278;
b_exp0 = 10'd1007; b_exp1 = 10'd377; b_exp2 = 10'd132; b_exp3 = 10'd118;
a_sign0 = 4'd9; a_sign1 = 4'd0; a_sign2 = 4'd15; a_sign3 = 4'd2;
b_sign0 = 4'd2; b_sign1 = 4'd11; b_sign2 = 4'd6; b_sign3 = 4'd4;
@(posedge clk_i);
a_mant0 = 8'd61; a_mant1 = 8'd118; a_mant2 = 8'd37; a_mant3 = 8'd48;
b_mant0 = 8'd34; b_mant1 = 8'd250; b_mant2 = 8'd55; b_mant3 = 8'd182;
a_exp0 = 10'd173; a_exp1 = 10'd196; a_exp2 = 10'd712; a_exp3 = 10'd454;
b_exp0 = 10'd817; b_exp1 = 10'd994; b_exp2 = 10'd166; b_exp3 = 10'd803;
a_sign0 = 4'd16; a_sign1 = 4'd0; a_sign2 = 4'd10; a_sign3 = 4'd8;
b_sign0 = 4'd1; b_sign1 = 4'd9; b_sign2 = 4'd3; b_sign3 = 4'd0;
@(posedge clk_i);
a_mant0 = 8'd105; a_mant1 = 8'd209; a_mant2 = 8'd228; a_mant3 = 8'd144;
b_mant0 = 8'd66; b_mant1 = 8'd112; b_mant2 = 8'd70; b_mant3 = 8'd201;
a_exp0 = 10'd342; a_exp1 = 10'd559; a_exp2 = 10'd72; a_exp3 = 10'd848;
b_exp0 = 10'd451; b_exp1 = 10'd799; b_exp2 = 10'd540; b_exp3 = 10'd97;
a_sign0 = 4'd6; a_sign1 = 4'd5; a_sign2 = 4'd2; a_sign3 = 4'd3;
b_sign0 = 4'd6; b_sign1 = 4'd3; b_sign2 = 4'd15; b_sign3 = 4'd5;
@(posedge clk_i);
a_mant0 = 8'd212; a_mant1 = 8'd184; a_mant2 = 8'd169; a_mant3 = 8'd26;
b_mant0 = 8'd206; b_mant1 = 8'd151; b_mant2 = 8'd252; b_mant3 = 8'd176;
a_exp0 = 10'd860; a_exp1 = 10'd537; a_exp2 = 10'd533; a_exp3 = 10'd775;
b_exp0 = 10'd948; b_exp1 = 10'd952; b_exp2 = 10'd857; b_exp3 = 10'd521;
a_sign0 = 4'd4; a_sign1 = 4'd4; a_sign2 = 4'd11; a_sign3 = 4'd14;
b_sign0 = 4'd10; b_sign1 = 4'd9; b_sign2 = 4'd7; b_sign3 = 4'd12;
@(posedge clk_i);
a_mant0 = 8'd252; a_mant1 = 8'd37; a_mant2 = 8'd98; a_mant3 = 8'd11;
b_mant0 = 8'd126; b_mant1 = 8'd231; b_mant2 = 8'd7; b_mant3 = 8'd82;
a_exp0 = 10'd982; a_exp1 = 10'd431; a_exp2 = 10'd522; a_exp3 = 10'd107;
b_exp0 = 10'd157; b_exp1 = 10'd614; b_exp2 = 10'd487; b_exp3 = 10'd7;
a_sign0 = 4'd13; a_sign1 = 4'd7; a_sign2 = 4'd4; a_sign3 = 4'd7;
b_sign0 = 4'd5; b_sign1 = 4'd16; b_sign2 = 4'd16; b_sign3 = 4'd10;
@(posedge clk_i);
a_mant0 = 8'd248; a_mant1 = 8'd9; a_mant2 = 8'd6; a_mant3 = 8'd70;
b_mant0 = 8'd198; b_mant1 = 8'd153; b_mant2 = 8'd135; b_mant3 = 8'd58;
a_exp0 = 10'd924; a_exp1 = 10'd818; a_exp2 = 10'd830; a_exp3 = 10'd113;
b_exp0 = 10'd745; b_exp1 = 10'd962; b_exp2 = 10'd781; b_exp3 = 10'd809;
a_sign0 = 4'd13; a_sign1 = 4'd9; a_sign2 = 4'd12; a_sign3 = 4'd6;
b_sign0 = 4'd8; b_sign1 = 4'd3; b_sign2 = 4'd1; b_sign3 = 4'd13;
@(posedge clk_i);
a_mant0 = 8'd4; a_mant1 = 8'd90; a_mant2 = 8'd227; a_mant3 = 8'd198;
b_mant0 = 8'd7; b_mant1 = 8'd52; b_mant2 = 8'd216; b_mant3 = 8'd104;
a_exp0 = 10'd815; a_exp1 = 10'd115; a_exp2 = 10'd599; a_exp3 = 10'd721;
b_exp0 = 10'd225; b_exp1 = 10'd982; b_exp2 = 10'd780; b_exp3 = 10'd53;
a_sign0 = 4'd9; a_sign1 = 4'd7; a_sign2 = 4'd0; a_sign3 = 4'd0;
b_sign0 = 4'd14; b_sign1 = 4'd11; b_sign2 = 4'd10; b_sign3 = 4'd4;
@(posedge clk_i);
shared_exps0 = 8'd132;
shared_exps1 = 8'd138;
rstn = 0;
@(posedge clk_i);
rstn = 1;
a_mant0 = 8'd59; a_mant1 = 8'd35; a_mant2 = 8'd230; a_mant3 = 8'd198;
b_mant0 = 8'd255; b_mant1 = 8'd50; b_mant2 = 8'd172; b_mant3 = 8'd154;
a_exp0 = 10'd334; a_exp1 = 10'd71; a_exp2 = 10'd302; a_exp3 = 10'd312;
b_exp0 = 10'd722; b_exp1 = 10'd262; b_exp2 = 10'd164; b_exp3 = 10'd838;
a_sign0 = 4'd7; a_sign1 = 4'd10; a_sign2 = 4'd16; a_sign3 = 4'd8;
b_sign0 = 4'd6; b_sign1 = 4'd10; b_sign2 = 4'd0; b_sign3 = 4'd2;
@(posedge clk_i);
a_mant0 = 8'd99; a_mant1 = 8'd205; a_mant2 = 8'd1; a_mant3 = 8'd178;
b_mant0 = 8'd155; b_mant1 = 8'd147; b_mant2 = 8'd221; b_mant3 = 8'd27;
a_exp0 = 10'd555; a_exp1 = 10'd258; a_exp2 = 10'd901; a_exp3 = 10'd30;
b_exp0 = 10'd986; b_exp1 = 10'd1016; b_exp2 = 10'd548; b_exp3 = 10'd486;
a_sign0 = 4'd9; a_sign1 = 4'd15; a_sign2 = 4'd1; a_sign3 = 4'd16;
b_sign0 = 4'd8; b_sign1 = 4'd10; b_sign2 = 4'd16; b_sign3 = 4'd2;
@(posedge clk_i);
a_mant0 = 8'd3; a_mant1 = 8'd167; a_mant2 = 8'd95; a_mant3 = 8'd35;
b_mant0 = 8'd17; b_mant1 = 8'd25; b_mant2 = 8'd24; b_mant3 = 8'd47;
a_exp0 = 10'd981; a_exp1 = 10'd955; a_exp2 = 10'd786; a_exp3 = 10'd457;
b_exp0 = 10'd837; b_exp1 = 10'd509; b_exp2 = 10'd204; b_exp3 = 10'd548;
a_sign0 = 4'd12; a_sign1 = 4'd7; a_sign2 = 4'd12; a_sign3 = 4'd9;
b_sign0 = 4'd3; b_sign1 = 4'd7; b_sign2 = 4'd11; b_sign3 = 4'd16;
@(posedge clk_i);
a_mant0 = 8'd16; a_mant1 = 8'd209; a_mant2 = 8'd67; a_mant3 = 8'd200;
b_mant0 = 8'd76; b_mant1 = 8'd186; b_mant2 = 8'd143; b_mant3 = 8'd119;
a_exp0 = 10'd145; a_exp1 = 10'd462; a_exp2 = 10'd189; a_exp3 = 10'd55;
b_exp0 = 10'd883; b_exp1 = 10'd966; b_exp2 = 10'd412; b_exp3 = 10'd1022;
a_sign0 = 4'd15; a_sign1 = 4'd8; a_sign2 = 4'd10; a_sign3 = 4'd6;
b_sign0 = 4'd11; b_sign1 = 4'd4; b_sign2 = 4'd12; b_sign3 = 4'd4;
@(posedge clk_i);
a_mant0 = 8'd116; a_mant1 = 8'd135; a_mant2 = 8'd178; a_mant3 = 8'd171;
b_mant0 = 8'd238; b_mant1 = 8'd190; b_mant2 = 8'd248; b_mant3 = 8'd251;
a_exp0 = 10'd341; a_exp1 = 10'd338; a_exp2 = 10'd214; a_exp3 = 10'd377;
b_exp0 = 10'd518; b_exp1 = 10'd249; b_exp2 = 10'd230; b_exp3 = 10'd483;
a_sign0 = 4'd9; a_sign1 = 4'd15; a_sign2 = 4'd0; a_sign3 = 4'd1;
b_sign0 = 4'd8; b_sign1 = 4'd7; b_sign2 = 4'd16; b_sign3 = 4'd13;
@(posedge clk_i);
a_mant0 = 8'd244; a_mant1 = 8'd182; a_mant2 = 8'd17; a_mant3 = 8'd17;
b_mant0 = 8'd244; b_mant1 = 8'd231; b_mant2 = 8'd25; b_mant3 = 8'd37;
a_exp0 = 10'd799; a_exp1 = 10'd174; a_exp2 = 10'd817; a_exp3 = 10'd250;
b_exp0 = 10'd989; b_exp1 = 10'd188; b_exp2 = 10'd679; b_exp3 = 10'd38;
a_sign0 = 4'd9; a_sign1 = 4'd8; a_sign2 = 4'd9; a_sign3 = 4'd6;
b_sign0 = 4'd6; b_sign1 = 4'd2; b_sign2 = 4'd12; b_sign3 = 4'd2;
@(posedge clk_i);
a_mant0 = 8'd249; a_mant1 = 8'd197; a_mant2 = 8'd116; a_mant3 = 8'd98;
b_mant0 = 8'd182; b_mant1 = 8'd3; b_mant2 = 8'd171; b_mant3 = 8'd248;
a_exp0 = 10'd988; a_exp1 = 10'd861; a_exp2 = 10'd459; a_exp3 = 10'd416;
b_exp0 = 10'd361; b_exp1 = 10'd650; b_exp2 = 10'd35; b_exp3 = 10'd217;
a_sign0 = 4'd3; a_sign1 = 4'd9; a_sign2 = 4'd2; a_sign3 = 4'd13;
b_sign0 = 4'd8; b_sign1 = 4'd5; b_sign2 = 4'd11; b_sign3 = 4'd4;
@(posedge clk_i);
shared_exps0 = 8'd99;
shared_exps1 = 8'd128;
a_mant0 = 8'd1; a_mant1 = 8'd18; a_mant2 = 8'd184; a_mant3 = 8'd254;
b_mant0 = 8'd254; b_mant1 = 8'd180; b_mant2 = 8'd34; b_mant3 = 8'd58;
a_exp0 = 10'd647; a_exp1 = 10'd460; a_exp2 = 10'd193; a_exp3 = 10'd525;
b_exp0 = 10'd728; b_exp1 = 10'd320; b_exp2 = 10'd165; b_exp3 = 10'd945;
a_sign0 = 4'd2; a_sign1 = 4'd4; a_sign2 = 4'd13; a_sign3 = 4'd5;
b_sign0 = 4'd2; b_sign1 = 4'd8; b_sign2 = 4'd12; b_sign3 = 4'd11;
@(posedge clk_i);
a_mant0 = 8'd118; a_mant1 = 8'd174; a_mant2 = 8'd111; a_mant3 = 8'd107;
b_mant0 = 8'd85; b_mant1 = 8'd77; b_mant2 = 8'd20; b_mant3 = 8'd107;
a_exp0 = 10'd351; a_exp1 = 10'd388; a_exp2 = 10'd1019; a_exp3 = 10'd426;
b_exp0 = 10'd920; b_exp1 = 10'd818; b_exp2 = 10'd199; b_exp3 = 10'd378;
a_sign0 = 4'd3; a_sign1 = 4'd8; a_sign2 = 4'd0; a_sign3 = 4'd2;
b_sign0 = 4'd11; b_sign1 = 4'd8; b_sign2 = 4'd3; b_sign3 = 4'd11;
@(posedge clk_i);
a_mant0 = 8'd58; a_mant1 = 8'd147; a_mant2 = 8'd45; a_mant3 = 8'd189;
b_mant0 = 8'd89; b_mant1 = 8'd24; b_mant2 = 8'd21; b_mant3 = 8'd231;
a_exp0 = 10'd444; a_exp1 = 10'd25; a_exp2 = 10'd269; a_exp3 = 10'd946;
b_exp0 = 10'd383; b_exp1 = 10'd323; b_exp2 = 10'd906; b_exp3 = 10'd92;
a_sign0 = 4'd5; a_sign1 = 4'd2; a_sign2 = 4'd10; a_sign3 = 4'd2;
b_sign0 = 4'd6; b_sign1 = 4'd8; b_sign2 = 4'd14; b_sign3 = 4'd11;
@(posedge clk_i);
a_mant0 = 8'd31; a_mant1 = 8'd167; a_mant2 = 8'd250; a_mant3 = 8'd200;
b_mant0 = 8'd168; b_mant1 = 8'd158; b_mant2 = 8'd145; b_mant3 = 8'd89;
a_exp0 = 10'd243; a_exp1 = 10'd481; a_exp2 = 10'd908; a_exp3 = 10'd662;
b_exp0 = 10'd146; b_exp1 = 10'd124; b_exp2 = 10'd741; b_exp3 = 10'd990;
a_sign0 = 4'd10; a_sign1 = 4'd2; a_sign2 = 4'd7; a_sign3 = 4'd15;
b_sign0 = 4'd16; b_sign1 = 4'd16; b_sign2 = 4'd5; b_sign3 = 4'd16;
@(posedge clk_i);
a_mant0 = 8'd19; a_mant1 = 8'd216; a_mant2 = 8'd182; a_mant3 = 8'd28;
b_mant0 = 8'd72; b_mant1 = 8'd5; b_mant2 = 8'd218; b_mant3 = 8'd164;
a_exp0 = 10'd158; a_exp1 = 10'd982; a_exp2 = 10'd747; a_exp3 = 10'd890;
b_exp0 = 10'd743; b_exp1 = 10'd199; b_exp2 = 10'd149; b_exp3 = 10'd708;
a_sign0 = 4'd15; a_sign1 = 4'd4; a_sign2 = 4'd7; a_sign3 = 4'd2;
b_sign0 = 4'd11; b_sign1 = 4'd14; b_sign2 = 4'd3; b_sign3 = 4'd3;
@(posedge clk_i);
a_mant0 = 8'd210; a_mant1 = 8'd49; a_mant2 = 8'd245; a_mant3 = 8'd125;
b_mant0 = 8'd130; b_mant1 = 8'd47; b_mant2 = 8'd225; b_mant3 = 8'd114;
a_exp0 = 10'd814; a_exp1 = 10'd920; a_exp2 = 10'd242; a_exp3 = 10'd252;
b_exp0 = 10'd651; b_exp1 = 10'd446; b_exp2 = 10'd202; b_exp3 = 10'd153;
a_sign0 = 4'd6; a_sign1 = 4'd11; a_sign2 = 4'd14; a_sign3 = 4'd3;
b_sign0 = 4'd8; b_sign1 = 4'd1; b_sign2 = 4'd8; b_sign3 = 4'd9;
@(posedge clk_i);
a_mant0 = 8'd69; a_mant1 = 8'd220; a_mant2 = 8'd151; a_mant3 = 8'd131;
b_mant0 = 8'd217; b_mant1 = 8'd255; b_mant2 = 8'd77; b_mant3 = 8'd73;
a_exp0 = 10'd644; a_exp1 = 10'd573; a_exp2 = 10'd979; a_exp3 = 10'd904;
b_exp0 = 10'd725; b_exp1 = 10'd319; b_exp2 = 10'd459; b_exp3 = 10'd937;
a_sign0 = 4'd5; a_sign1 = 4'd7; a_sign2 = 4'd11; a_sign3 = 4'd6;
b_sign0 = 4'd2; b_sign1 = 4'd6; b_sign2 = 4'd16; b_sign3 = 4'd6;
@(posedge clk_i);
a_mant0 = 8'd6; a_mant1 = 8'd184; a_mant2 = 8'd43; a_mant3 = 8'd197;
b_mant0 = 8'd238; b_mant1 = 8'd211; b_mant2 = 8'd254; b_mant3 = 8'd147;
a_exp0 = 10'd891; a_exp1 = 10'd697; a_exp2 = 10'd477; a_exp3 = 10'd151;
b_exp0 = 10'd716; b_exp1 = 10'd794; b_exp2 = 10'd449; b_exp3 = 10'd181;
a_sign0 = 4'd0; a_sign1 = 4'd16; a_sign2 = 4'd0; a_sign3 = 4'd2;
b_sign0 = 4'd0; b_sign1 = 4'd3; b_sign2 = 4'd4; b_sign3 = 4'd3;
@(posedge clk_i);
shared_exps0 = 8'd137;
shared_exps1 = 8'd125;
a_mant0 = 8'd178; a_mant1 = 8'd189; a_mant2 = 8'd186; a_mant3 = 8'd178;
b_mant0 = 8'd91; b_mant1 = 8'd214; b_mant2 = 8'd123; b_mant3 = 8'd137;
a_exp0 = 10'd350; a_exp1 = 10'd285; a_exp2 = 10'd602; a_exp3 = 10'd140;
b_exp0 = 10'd89; b_exp1 = 10'd654; b_exp2 = 10'd461; b_exp3 = 10'd258;
a_sign0 = 4'd0; a_sign1 = 4'd11; a_sign2 = 4'd13; a_sign3 = 4'd3;
b_sign0 = 4'd10; b_sign1 = 4'd8; b_sign2 = 4'd0; b_sign3 = 4'd13;
@(posedge clk_i);
a_mant0 = 8'd65; a_mant1 = 8'd53; a_mant2 = 8'd202; a_mant3 = 8'd156;
b_mant0 = 8'd21; b_mant1 = 8'd106; b_mant2 = 8'd55; b_mant3 = 8'd78;
a_exp0 = 10'd610; a_exp1 = 10'd965; a_exp2 = 10'd1023; a_exp3 = 10'd856;
b_exp0 = 10'd469; b_exp1 = 10'd246; b_exp2 = 10'd751; b_exp3 = 10'd2;
a_sign0 = 4'd6; a_sign1 = 4'd10; a_sign2 = 4'd11; a_sign3 = 4'd6;
b_sign0 = 4'd12; b_sign1 = 4'd13; b_sign2 = 4'd0; b_sign3 = 4'd10;
@(posedge clk_i);
a_mant0 = 8'd241; a_mant1 = 8'd229; a_mant2 = 8'd169; a_mant3 = 8'd179;
b_mant0 = 8'd98; b_mant1 = 8'd174; b_mant2 = 8'd54; b_mant3 = 8'd253;
a_exp0 = 10'd686; a_exp1 = 10'd340; a_exp2 = 10'd1018; a_exp3 = 10'd27;
b_exp0 = 10'd26; b_exp1 = 10'd937; b_exp2 = 10'd349; b_exp3 = 10'd814;
a_sign0 = 4'd10; a_sign1 = 4'd3; a_sign2 = 4'd4; a_sign3 = 4'd5;
b_sign0 = 4'd14; b_sign1 = 4'd14; b_sign2 = 4'd0; b_sign3 = 4'd0;
@(posedge clk_i);
a_mant0 = 8'd19; a_mant1 = 8'd84; a_mant2 = 8'd221; a_mant3 = 8'd217;
b_mant0 = 8'd50; b_mant1 = 8'd127; b_mant2 = 8'd81; b_mant3 = 8'd122;
a_exp0 = 10'd787; a_exp1 = 10'd285; a_exp2 = 10'd573; a_exp3 = 10'd972;
b_exp0 = 10'd18; b_exp1 = 10'd465; b_exp2 = 10'd843; b_exp3 = 10'd925;
a_sign0 = 4'd16; a_sign1 = 4'd4; a_sign2 = 4'd16; a_sign3 = 4'd4;
b_sign0 = 4'd1; b_sign1 = 4'd12; b_sign2 = 4'd11; b_sign3 = 4'd4;
@(posedge clk_i);
a_mant0 = 8'd211; a_mant1 = 8'd211; a_mant2 = 8'd33; a_mant3 = 8'd163;
b_mant0 = 8'd42; b_mant1 = 8'd242; b_mant2 = 8'd163; b_mant3 = 8'd180;
a_exp0 = 10'd208; a_exp1 = 10'd486; a_exp2 = 10'd581; a_exp3 = 10'd989;
b_exp0 = 10'd626; b_exp1 = 10'd975; b_exp2 = 10'd949; b_exp3 = 10'd642;
a_sign0 = 4'd11; a_sign1 = 4'd12; a_sign2 = 4'd1; a_sign3 = 4'd2;
b_sign0 = 4'd2; b_sign1 = 4'd12; b_sign2 = 4'd8; b_sign3 = 4'd0;
@(posedge clk_i);
a_mant0 = 8'd8; a_mant1 = 8'd51; a_mant2 = 8'd148; a_mant3 = 8'd61;
b_mant0 = 8'd58; b_mant1 = 8'd65; b_mant2 = 8'd124; b_mant3 = 8'd39;
a_exp0 = 10'd265; a_exp1 = 10'd173; a_exp2 = 10'd879; a_exp3 = 10'd184;
b_exp0 = 10'd990; b_exp1 = 10'd105; b_exp2 = 10'd899; b_exp3 = 10'd107;
a_sign0 = 4'd5; a_sign1 = 4'd5; a_sign2 = 4'd9; a_sign3 = 4'd1;
b_sign0 = 4'd2; b_sign1 = 4'd1; b_sign2 = 4'd14; b_sign3 = 4'd2;
@(posedge clk_i);
a_mant0 = 8'd231; a_mant1 = 8'd18; a_mant2 = 8'd212; a_mant3 = 8'd91;
b_mant0 = 8'd219; b_mant1 = 8'd126; b_mant2 = 8'd158; b_mant3 = 8'd142;
a_exp0 = 10'd147; a_exp1 = 10'd986; a_exp2 = 10'd1016; a_exp3 = 10'd926;
b_exp0 = 10'd496; b_exp1 = 10'd918; b_exp2 = 10'd958; b_exp3 = 10'd92;
a_sign0 = 4'd3; a_sign1 = 4'd13; a_sign2 = 4'd6; a_sign3 = 4'd4;
b_sign0 = 4'd10; b_sign1 = 4'd14; b_sign2 = 4'd4; b_sign3 = 4'd2;
@(posedge clk_i);
a_mant0 = 8'd74; a_mant1 = 8'd53; a_mant2 = 8'd46; a_mant3 = 8'd94;
b_mant0 = 8'd95; b_mant1 = 8'd132; b_mant2 = 8'd72; b_mant3 = 8'd154;
a_exp0 = 10'd517; a_exp1 = 10'd6; a_exp2 = 10'd148; a_exp3 = 10'd603;
b_exp0 = 10'd835; b_exp1 = 10'd446; b_exp2 = 10'd183; b_exp3 = 10'd266;
a_sign0 = 4'd10; a_sign1 = 4'd6; a_sign2 = 4'd15; a_sign3 = 4'd11;
b_sign0 = 4'd9; b_sign1 = 4'd8; b_sign2 = 4'd7; b_sign3 = 4'd16;
@(posedge clk_i);
shared_exps0 = 8'd120;
shared_exps1 = 8'd143;
a_mant0 = 8'd171; a_mant1 = 8'd201; a_mant2 = 8'd16; a_mant3 = 8'd194;
b_mant0 = 8'd221; b_mant1 = 8'd109; b_mant2 = 8'd245; b_mant3 = 8'd191;
a_exp0 = 10'd424; a_exp1 = 10'd61; a_exp2 = 10'd979; a_exp3 = 10'd28;
b_exp0 = 10'd545; b_exp1 = 10'd95; b_exp2 = 10'd473; b_exp3 = 10'd261;
a_sign0 = 4'd13; a_sign1 = 4'd14; a_sign2 = 4'd3; a_sign3 = 4'd6;
b_sign0 = 4'd13; b_sign1 = 4'd12; b_sign2 = 4'd5; b_sign3 = 4'd7;
@(posedge clk_i);
a_mant0 = 8'd67; a_mant1 = 8'd62; a_mant2 = 8'd138; a_mant3 = 8'd99;
b_mant0 = 8'd155; b_mant1 = 8'd154; b_mant2 = 8'd20; b_mant3 = 8'd190;
a_exp0 = 10'd71; a_exp1 = 10'd143; a_exp2 = 10'd216; a_exp3 = 10'd220;
b_exp0 = 10'd202; b_exp1 = 10'd434; b_exp2 = 10'd493; b_exp3 = 10'd947;
a_sign0 = 4'd1; a_sign1 = 4'd16; a_sign2 = 4'd15; a_sign3 = 4'd15;
b_sign0 = 4'd2; b_sign1 = 4'd10; b_sign2 = 4'd10; b_sign3 = 4'd0;
@(posedge clk_i);
a_mant0 = 8'd36; a_mant1 = 8'd7; a_mant2 = 8'd250; a_mant3 = 8'd113;
b_mant0 = 8'd242; b_mant1 = 8'd116; b_mant2 = 8'd41; b_mant3 = 8'd215;
a_exp0 = 10'd881; a_exp1 = 10'd907; a_exp2 = 10'd218; a_exp3 = 10'd537;
b_exp0 = 10'd46; b_exp1 = 10'd83; b_exp2 = 10'd57; b_exp3 = 10'd918;
a_sign0 = 4'd8; a_sign1 = 4'd16; a_sign2 = 4'd15; a_sign3 = 4'd10;
b_sign0 = 4'd8; b_sign1 = 4'd6; b_sign2 = 4'd1; b_sign3 = 4'd10;
@(posedge clk_i);
a_mant0 = 8'd20; a_mant1 = 8'd168; a_mant2 = 8'd105; a_mant3 = 8'd131;
b_mant0 = 8'd177; b_mant1 = 8'd241; b_mant2 = 8'd182; b_mant3 = 8'd26;
a_exp0 = 10'd288; a_exp1 = 10'd545; a_exp2 = 10'd868; a_exp3 = 10'd720;
b_exp0 = 10'd502; b_exp1 = 10'd976; b_exp2 = 10'd890; b_exp3 = 10'd402;
a_sign0 = 4'd11; a_sign1 = 4'd8; a_sign2 = 4'd6; a_sign3 = 4'd3;
b_sign0 = 4'd16; b_sign1 = 4'd3; b_sign2 = 4'd11; b_sign3 = 4'd0;
@(posedge clk_i);
a_mant0 = 8'd208; a_mant1 = 8'd183; a_mant2 = 8'd200; a_mant3 = 8'd248;
b_mant0 = 8'd172; b_mant1 = 8'd46; b_mant2 = 8'd24; b_mant3 = 8'd43;
a_exp0 = 10'd512; a_exp1 = 10'd537; a_exp2 = 10'd218; a_exp3 = 10'd771;
b_exp0 = 10'd259; b_exp1 = 10'd263; b_exp2 = 10'd290; b_exp3 = 10'd226;
a_sign0 = 4'd11; a_sign1 = 4'd2; a_sign2 = 4'd2; a_sign3 = 4'd2;
b_sign0 = 4'd12; b_sign1 = 4'd7; b_sign2 = 4'd12; b_sign3 = 4'd3;
@(posedge clk_i);
a_mant0 = 8'd136; a_mant1 = 8'd180; a_mant2 = 8'd116; a_mant3 = 8'd136;
b_mant0 = 8'd204; b_mant1 = 8'd121; b_mant2 = 8'd231; b_mant3 = 8'd92;
a_exp0 = 10'd30; a_exp1 = 10'd352; a_exp2 = 10'd610; a_exp3 = 10'd950;
b_exp0 = 10'd445; b_exp1 = 10'd760; b_exp2 = 10'd263; b_exp3 = 10'd507;
a_sign0 = 4'd3; a_sign1 = 4'd15; a_sign2 = 4'd1; a_sign3 = 4'd7;
b_sign0 = 4'd5; b_sign1 = 4'd0; b_sign2 = 4'd10; b_sign3 = 4'd3;
@(posedge clk_i);
a_mant0 = 8'd35; a_mant1 = 8'd149; a_mant2 = 8'd75; a_mant3 = 8'd90;
b_mant0 = 8'd80; b_mant1 = 8'd94; b_mant2 = 8'd177; b_mant3 = 8'd166;
a_exp0 = 10'd312; a_exp1 = 10'd798; a_exp2 = 10'd823; a_exp3 = 10'd667;
b_exp0 = 10'd73; b_exp1 = 10'd639; b_exp2 = 10'd423; b_exp3 = 10'd142;
a_sign0 = 4'd3; a_sign1 = 4'd12; a_sign2 = 4'd13; a_sign3 = 4'd9;
b_sign0 = 4'd5; b_sign1 = 4'd3; b_sign2 = 4'd15; b_sign3 = 4'd3;
@(posedge clk_i);
a_mant0 = 8'd13; a_mant1 = 8'd10; a_mant2 = 8'd214; a_mant3 = 8'd79;
b_mant0 = 8'd190; b_mant1 = 8'd129; b_mant2 = 8'd70; b_mant3 = 8'd89;
a_exp0 = 10'd198; a_exp1 = 10'd364; a_exp2 = 10'd535; a_exp3 = 10'd716;
b_exp0 = 10'd470; b_exp1 = 10'd179; b_exp2 = 10'd99; b_exp3 = 10'd370;
a_sign0 = 4'd11; a_sign1 = 4'd9; a_sign2 = 4'd8; a_sign3 = 4'd10;
b_sign0 = 4'd12; b_sign1 = 4'd4; b_sign2 = 4'd9; b_sign3 = 4'd10;
@(posedge clk_i);
shared_exps0 = 8'd124;
shared_exps1 = 8'd144;
rstn = 0;
@(posedge clk_i);
rstn = 1;
a_mant0 = 8'd249; a_mant1 = 8'd76; a_mant2 = 8'd156; a_mant3 = 8'd224;
b_mant0 = 8'd59; b_mant1 = 8'd235; b_mant2 = 8'd207; b_mant3 = 8'd26;
a_exp0 = 10'd1023; a_exp1 = 10'd871; a_exp2 = 10'd113; a_exp3 = 10'd176;
b_exp0 = 10'd917; b_exp1 = 10'd867; b_exp2 = 10'd893; b_exp3 = 10'd834;
a_sign0 = 4'd12; a_sign1 = 4'd6; a_sign2 = 4'd2; a_sign3 = 4'd1;
b_sign0 = 4'd4; b_sign1 = 4'd5; b_sign2 = 4'd10; b_sign3 = 4'd9;
@(posedge clk_i);
a_mant0 = 8'd35; a_mant1 = 8'd1; a_mant2 = 8'd59; a_mant3 = 8'd180;
b_mant0 = 8'd126; b_mant1 = 8'd28; b_mant2 = 8'd98; b_mant3 = 8'd50;
a_exp0 = 10'd59; a_exp1 = 10'd888; a_exp2 = 10'd751; a_exp3 = 10'd493;
b_exp0 = 10'd998; b_exp1 = 10'd663; b_exp2 = 10'd101; b_exp3 = 10'd778;
a_sign0 = 4'd7; a_sign1 = 4'd7; a_sign2 = 4'd15; a_sign3 = 4'd15;
b_sign0 = 4'd10; b_sign1 = 4'd16; b_sign2 = 4'd8; b_sign3 = 4'd9;
@(posedge clk_i);
a_mant0 = 8'd137; a_mant1 = 8'd39; a_mant2 = 8'd209; a_mant3 = 8'd139;
b_mant0 = 8'd90; b_mant1 = 8'd95; b_mant2 = 8'd198; b_mant3 = 8'd168;
a_exp0 = 10'd478; a_exp1 = 10'd685; a_exp2 = 10'd762; a_exp3 = 10'd851;
b_exp0 = 10'd559; b_exp1 = 10'd775; b_exp2 = 10'd145; b_exp3 = 10'd718;
a_sign0 = 4'd12; a_sign1 = 4'd5; a_sign2 = 4'd16; a_sign3 = 4'd16;
b_sign0 = 4'd10; b_sign1 = 4'd0; b_sign2 = 4'd5; b_sign3 = 4'd3;
@(posedge clk_i);
a_mant0 = 8'd243; a_mant1 = 8'd121; a_mant2 = 8'd109; a_mant3 = 8'd195;
b_mant0 = 8'd248; b_mant1 = 8'd121; b_mant2 = 8'd228; b_mant3 = 8'd88;
a_exp0 = 10'd607; a_exp1 = 10'd172; a_exp2 = 10'd605; a_exp3 = 10'd829;
b_exp0 = 10'd162; b_exp1 = 10'd48; b_exp2 = 10'd540; b_exp3 = 10'd215;
a_sign0 = 4'd0; a_sign1 = 4'd4; a_sign2 = 4'd10; a_sign3 = 4'd6;
b_sign0 = 4'd8; b_sign1 = 4'd14; b_sign2 = 4'd16; b_sign3 = 4'd3;
@(posedge clk_i);
a_mant0 = 8'd207; a_mant1 = 8'd76; a_mant2 = 8'd43; a_mant3 = 8'd154;
b_mant0 = 8'd187; b_mant1 = 8'd108; b_mant2 = 8'd106; b_mant3 = 8'd235;
a_exp0 = 10'd244; a_exp1 = 10'd427; a_exp2 = 10'd195; a_exp3 = 10'd315;
b_exp0 = 10'd66; b_exp1 = 10'd254; b_exp2 = 10'd364; b_exp3 = 10'd919;
a_sign0 = 4'd16; a_sign1 = 4'd14; a_sign2 = 4'd7; a_sign3 = 4'd14;
b_sign0 = 4'd14; b_sign1 = 4'd2; b_sign2 = 4'd7; b_sign3 = 4'd9;
@(posedge clk_i);
a_mant0 = 8'd19; a_mant1 = 8'd203; a_mant2 = 8'd174; a_mant3 = 8'd102;
b_mant0 = 8'd146; b_mant1 = 8'd146; b_mant2 = 8'd141; b_mant3 = 8'd167;
a_exp0 = 10'd514; a_exp1 = 10'd990; a_exp2 = 10'd716; a_exp3 = 10'd498;
b_exp0 = 10'd448; b_exp1 = 10'd846; b_exp2 = 10'd411; b_exp3 = 10'd329;
a_sign0 = 4'd8; a_sign1 = 4'd2; a_sign2 = 4'd6; a_sign3 = 4'd13;
b_sign0 = 4'd5; b_sign1 = 4'd12; b_sign2 = 4'd0; b_sign3 = 4'd16;
@(posedge clk_i);
a_mant0 = 8'd18; a_mant1 = 8'd112; a_mant2 = 8'd183; a_mant3 = 8'd193;
b_mant0 = 8'd46; b_mant1 = 8'd108; b_mant2 = 8'd39; b_mant3 = 8'd164;
a_exp0 = 10'd686; a_exp1 = 10'd249; a_exp2 = 10'd281; a_exp3 = 10'd1018;
b_exp0 = 10'd873; b_exp1 = 10'd562; b_exp2 = 10'd520; b_exp3 = 10'd845;
a_sign0 = 4'd0; a_sign1 = 4'd14; a_sign2 = 4'd1; a_sign3 = 4'd7;
b_sign0 = 4'd14; b_sign1 = 4'd15; b_sign2 = 4'd7; b_sign3 = 4'd11;
@(posedge clk_i);
shared_exps0 = 8'd107;
shared_exps1 = 8'd120;
a_mant0 = 8'd147; a_mant1 = 8'd95; a_mant2 = 8'd14; a_mant3 = 8'd85;
b_mant0 = 8'd150; b_mant1 = 8'd34; b_mant2 = 8'd220; b_mant3 = 8'd219;
a_exp0 = 10'd757; a_exp1 = 10'd377; a_exp2 = 10'd195; a_exp3 = 10'd736;
b_exp0 = 10'd584; b_exp1 = 10'd503; b_exp2 = 10'd797; b_exp3 = 10'd311;
a_sign0 = 4'd5; a_sign1 = 4'd3; a_sign2 = 4'd5; a_sign3 = 4'd7;
b_sign0 = 4'd0; b_sign1 = 4'd4; b_sign2 = 4'd3; b_sign3 = 4'd1;
@(posedge clk_i);
a_mant0 = 8'd79; a_mant1 = 8'd64; a_mant2 = 8'd50; a_mant3 = 8'd71;
b_mant0 = 8'd155; b_mant1 = 8'd190; b_mant2 = 8'd150; b_mant3 = 8'd221;
a_exp0 = 10'd959; a_exp1 = 10'd296; a_exp2 = 10'd864; a_exp3 = 10'd645;
b_exp0 = 10'd880; b_exp1 = 10'd875; b_exp2 = 10'd584; b_exp3 = 10'd467;
a_sign0 = 4'd7; a_sign1 = 4'd2; a_sign2 = 4'd12; a_sign3 = 4'd12;
b_sign0 = 4'd14; b_sign1 = 4'd16; b_sign2 = 4'd8; b_sign3 = 4'd4;
@(posedge clk_i);
a_mant0 = 8'd249; a_mant1 = 8'd56; a_mant2 = 8'd135; a_mant3 = 8'd238;
b_mant0 = 8'd206; b_mant1 = 8'd251; b_mant2 = 8'd87; b_mant3 = 8'd194;
a_exp0 = 10'd566; a_exp1 = 10'd983; a_exp2 = 10'd28; a_exp3 = 10'd300;
b_exp0 = 10'd531; b_exp1 = 10'd239; b_exp2 = 10'd22; b_exp3 = 10'd926;
a_sign0 = 4'd5; a_sign1 = 4'd2; a_sign2 = 4'd16; a_sign3 = 4'd9;
b_sign0 = 4'd15; b_sign1 = 4'd8; b_sign2 = 4'd15; b_sign3 = 4'd12;
@(posedge clk_i);
a_mant0 = 8'd36; a_mant1 = 8'd118; a_mant2 = 8'd155; a_mant3 = 8'd49;
b_mant0 = 8'd84; b_mant1 = 8'd200; b_mant2 = 8'd39; b_mant3 = 8'd241;
a_exp0 = 10'd832; a_exp1 = 10'd140; a_exp2 = 10'd466; a_exp3 = 10'd1023;
b_exp0 = 10'd770; b_exp1 = 10'd736; b_exp2 = 10'd241; b_exp3 = 10'd786;
a_sign0 = 4'd8; a_sign1 = 4'd14; a_sign2 = 4'd10; a_sign3 = 4'd15;
b_sign0 = 4'd9; b_sign1 = 4'd4; b_sign2 = 4'd3; b_sign3 = 4'd16;
@(posedge clk_i);
a_mant0 = 8'd248; a_mant1 = 8'd20; a_mant2 = 8'd247; a_mant3 = 8'd8;
b_mant0 = 8'd120; b_mant1 = 8'd140; b_mant2 = 8'd236; b_mant3 = 8'd78;
a_exp0 = 10'd872; a_exp1 = 10'd788; a_exp2 = 10'd333; a_exp3 = 10'd8;
b_exp0 = 10'd591; b_exp1 = 10'd716; b_exp2 = 10'd664; b_exp3 = 10'd615;
a_sign0 = 4'd8; a_sign1 = 4'd9; a_sign2 = 4'd5; a_sign3 = 4'd13;
b_sign0 = 4'd10; b_sign1 = 4'd11; b_sign2 = 4'd13; b_sign3 = 4'd16;
@(posedge clk_i);
a_mant0 = 8'd49; a_mant1 = 8'd29; a_mant2 = 8'd94; a_mant3 = 8'd173;
b_mant0 = 8'd82; b_mant1 = 8'd38; b_mant2 = 8'd51; b_mant3 = 8'd75;
a_exp0 = 10'd809; a_exp1 = 10'd321; a_exp2 = 10'd224; a_exp3 = 10'd803;
b_exp0 = 10'd749; b_exp1 = 10'd773; b_exp2 = 10'd112; b_exp3 = 10'd908;
a_sign0 = 4'd11; a_sign1 = 4'd2; a_sign2 = 4'd5; a_sign3 = 4'd2;
b_sign0 = 4'd8; b_sign1 = 4'd16; b_sign2 = 4'd5; b_sign3 = 4'd14;
@(posedge clk_i);
a_mant0 = 8'd148; a_mant1 = 8'd79; a_mant2 = 8'd100; a_mant3 = 8'd127;
b_mant0 = 8'd54; b_mant1 = 8'd78; b_mant2 = 8'd198; b_mant3 = 8'd60;
a_exp0 = 10'd270; a_exp1 = 10'd1023; a_exp2 = 10'd724; a_exp3 = 10'd489;
b_exp0 = 10'd25; b_exp1 = 10'd429; b_exp2 = 10'd620; b_exp3 = 10'd1014;
a_sign0 = 4'd16; a_sign1 = 4'd12; a_sign2 = 4'd9; a_sign3 = 4'd5;
b_sign0 = 4'd12; b_sign1 = 4'd9; b_sign2 = 4'd0; b_sign3 = 4'd0;
@(posedge clk_i);
a_mant0 = 8'd78; a_mant1 = 8'd150; a_mant2 = 8'd125; a_mant3 = 8'd128;
b_mant0 = 8'd122; b_mant1 = 8'd228; b_mant2 = 8'd186; b_mant3 = 8'd176;
a_exp0 = 10'd597; a_exp1 = 10'd545; a_exp2 = 10'd431; a_exp3 = 10'd57;
b_exp0 = 10'd58; b_exp1 = 10'd778; b_exp2 = 10'd50; b_exp3 = 10'd928;
a_sign0 = 4'd6; a_sign1 = 4'd5; a_sign2 = 4'd7; a_sign3 = 4'd14;
b_sign0 = 4'd3; b_sign1 = 4'd1; b_sign2 = 4'd15; b_sign3 = 4'd10;
@(posedge clk_i);
shared_exps0 = 8'd116;
shared_exps1 = 8'd150;
a_mant0 = 8'd216; a_mant1 = 8'd221; a_mant2 = 8'd85; a_mant3 = 8'd146;
b_mant0 = 8'd76; b_mant1 = 8'd123; b_mant2 = 8'd223; b_mant3 = 8'd186;
a_exp0 = 10'd710; a_exp1 = 10'd539; a_exp2 = 10'd626; a_exp3 = 10'd916;
b_exp0 = 10'd671; b_exp1 = 10'd176; b_exp2 = 10'd932; b_exp3 = 10'd845;
a_sign0 = 4'd12; a_sign1 = 4'd13; a_sign2 = 4'd11; a_sign3 = 4'd5;
b_sign0 = 4'd16; b_sign1 = 4'd15; b_sign2 = 4'd13; b_sign3 = 4'd14;
@(posedge clk_i);
a_mant0 = 8'd21; a_mant1 = 8'd146; a_mant2 = 8'd72; a_mant3 = 8'd174;
b_mant0 = 8'd113; b_mant1 = 8'd224; b_mant2 = 8'd215; b_mant3 = 8'd228;
a_exp0 = 10'd505; a_exp1 = 10'd672; a_exp2 = 10'd758; a_exp3 = 10'd928;
b_exp0 = 10'd879; b_exp1 = 10'd502; b_exp2 = 10'd57; b_exp3 = 10'd872;
a_sign0 = 4'd3; a_sign1 = 4'd0; a_sign2 = 4'd11; a_sign3 = 4'd15;
b_sign0 = 4'd13; b_sign1 = 4'd9; b_sign2 = 4'd12; b_sign3 = 4'd11;
@(posedge clk_i);
a_mant0 = 8'd84; a_mant1 = 8'd174; a_mant2 = 8'd71; a_mant3 = 8'd93;
b_mant0 = 8'd92; b_mant1 = 8'd18; b_mant2 = 8'd235; b_mant3 = 8'd126;
a_exp0 = 10'd379; a_exp1 = 10'd762; a_exp2 = 10'd1004; a_exp3 = 10'd449;
b_exp0 = 10'd746; b_exp1 = 10'd505; b_exp2 = 10'd286; b_exp3 = 10'd147;
a_sign0 = 4'd14; a_sign1 = 4'd15; a_sign2 = 4'd13; a_sign3 = 4'd8;
b_sign0 = 4'd11; b_sign1 = 4'd13; b_sign2 = 4'd16; b_sign3 = 4'd1;
@(posedge clk_i);
a_mant0 = 8'd78; a_mant1 = 8'd234; a_mant2 = 8'd244; a_mant3 = 8'd227;
b_mant0 = 8'd236; b_mant1 = 8'd146; b_mant2 = 8'd27; b_mant3 = 8'd242;
a_exp0 = 10'd707; a_exp1 = 10'd995; a_exp2 = 10'd57; a_exp3 = 10'd244;
b_exp0 = 10'd773; b_exp1 = 10'd376; b_exp2 = 10'd48; b_exp3 = 10'd886;
a_sign0 = 4'd5; a_sign1 = 4'd0; a_sign2 = 4'd15; a_sign3 = 4'd6;
b_sign0 = 4'd5; b_sign1 = 4'd11; b_sign2 = 4'd5; b_sign3 = 4'd2;
@(posedge clk_i);
a_mant0 = 8'd211; a_mant1 = 8'd60; a_mant2 = 8'd46; a_mant3 = 8'd184;
b_mant0 = 8'd254; b_mant1 = 8'd114; b_mant2 = 8'd158; b_mant3 = 8'd254;
a_exp0 = 10'd598; a_exp1 = 10'd504; a_exp2 = 10'd994; a_exp3 = 10'd233;
b_exp0 = 10'd203; b_exp1 = 10'd22; b_exp2 = 10'd443; b_exp3 = 10'd254;
a_sign0 = 4'd7; a_sign1 = 4'd2; a_sign2 = 4'd2; a_sign3 = 4'd10;
b_sign0 = 4'd0; b_sign1 = 4'd0; b_sign2 = 4'd6; b_sign3 = 4'd3;
@(posedge clk_i);
a_mant0 = 8'd72; a_mant1 = 8'd190; a_mant2 = 8'd85; a_mant3 = 8'd56;
b_mant0 = 8'd71; b_mant1 = 8'd118; b_mant2 = 8'd3; b_mant3 = 8'd12;
a_exp0 = 10'd605; a_exp1 = 10'd810; a_exp2 = 10'd350; a_exp3 = 10'd744;
b_exp0 = 10'd573; b_exp1 = 10'd147; b_exp2 = 10'd141; b_exp3 = 10'd145;
a_sign0 = 4'd0; a_sign1 = 4'd13; a_sign2 = 4'd0; a_sign3 = 4'd5;
b_sign0 = 4'd5; b_sign1 = 4'd7; b_sign2 = 4'd5; b_sign3 = 4'd7;
@(posedge clk_i);
a_mant0 = 8'd35; a_mant1 = 8'd146; a_mant2 = 8'd195; a_mant3 = 8'd67;
b_mant0 = 8'd210; b_mant1 = 8'd68; b_mant2 = 8'd98; b_mant3 = 8'd1;
a_exp0 = 10'd509; a_exp1 = 10'd576; a_exp2 = 10'd564; a_exp3 = 10'd541;
b_exp0 = 10'd846; b_exp1 = 10'd724; b_exp2 = 10'd672; b_exp3 = 10'd279;
a_sign0 = 4'd9; a_sign1 = 4'd11; a_sign2 = 4'd2; a_sign3 = 4'd6;
b_sign0 = 4'd10; b_sign1 = 4'd7; b_sign2 = 4'd1; b_sign3 = 4'd14;
@(posedge clk_i);
a_mant0 = 8'd26; a_mant1 = 8'd236; a_mant2 = 8'd146; a_mant3 = 8'd69;
b_mant0 = 8'd157; b_mant1 = 8'd221; b_mant2 = 8'd245; b_mant3 = 8'd98;
a_exp0 = 10'd814; a_exp1 = 10'd320; a_exp2 = 10'd757; a_exp3 = 10'd388;
b_exp0 = 10'd482; b_exp1 = 10'd399; b_exp2 = 10'd299; b_exp3 = 10'd122;
a_sign0 = 4'd13; a_sign1 = 4'd13; a_sign2 = 4'd8; a_sign3 = 4'd16;
b_sign0 = 4'd4; b_sign1 = 4'd4; b_sign2 = 4'd15; b_sign3 = 4'd11;
@(posedge clk_i);
shared_exps0 = 8'd155;
shared_exps1 = 8'd135;
a_mant0 = 8'd243; a_mant1 = 8'd20; a_mant2 = 8'd242; a_mant3 = 8'd235;
b_mant0 = 8'd23; b_mant1 = 8'd38; b_mant2 = 8'd224; b_mant3 = 8'd46;
a_exp0 = 10'd985; a_exp1 = 10'd27; a_exp2 = 10'd566; a_exp3 = 10'd330;
b_exp0 = 10'd883; b_exp1 = 10'd203; b_exp2 = 10'd403; b_exp3 = 10'd960;
a_sign0 = 4'd7; a_sign1 = 4'd12; a_sign2 = 4'd10; a_sign3 = 4'd0;
b_sign0 = 4'd5; b_sign1 = 4'd2; b_sign2 = 4'd12; b_sign3 = 4'd2;
@(posedge clk_i);
a_mant0 = 8'd86; a_mant1 = 8'd25; a_mant2 = 8'd219; a_mant3 = 8'd218;
b_mant0 = 8'd39; b_mant1 = 8'd59; b_mant2 = 8'd219; b_mant3 = 8'd156;
a_exp0 = 10'd614; a_exp1 = 10'd451; a_exp2 = 10'd872; a_exp3 = 10'd502;
b_exp0 = 10'd136; b_exp1 = 10'd363; b_exp2 = 10'd692; b_exp3 = 10'd312;
a_sign0 = 4'd6; a_sign1 = 4'd8; a_sign2 = 4'd5; a_sign3 = 4'd14;
b_sign0 = 4'd10; b_sign1 = 4'd4; b_sign2 = 4'd11; b_sign3 = 4'd13;
@(posedge clk_i);
a_mant0 = 8'd57; a_mant1 = 8'd168; a_mant2 = 8'd13; a_mant3 = 8'd237;
b_mant0 = 8'd124; b_mant1 = 8'd92; b_mant2 = 8'd167; b_mant3 = 8'd254;
a_exp0 = 10'd299; a_exp1 = 10'd395; a_exp2 = 10'd929; a_exp3 = 10'd858;
b_exp0 = 10'd165; b_exp1 = 10'd670; b_exp2 = 10'd528; b_exp3 = 10'd91;
a_sign0 = 4'd7; a_sign1 = 4'd5; a_sign2 = 4'd16; a_sign3 = 4'd12;
b_sign0 = 4'd12; b_sign1 = 4'd10; b_sign2 = 4'd10; b_sign3 = 4'd3;
@(posedge clk_i);
a_mant0 = 8'd126; a_mant1 = 8'd189; a_mant2 = 8'd247; a_mant3 = 8'd161;
b_mant0 = 8'd56; b_mant1 = 8'd220; b_mant2 = 8'd31; b_mant3 = 8'd18;
a_exp0 = 10'd304; a_exp1 = 10'd978; a_exp2 = 10'd557; a_exp3 = 10'd542;
b_exp0 = 10'd741; b_exp1 = 10'd598; b_exp2 = 10'd541; b_exp3 = 10'd508;
a_sign0 = 4'd12; a_sign1 = 4'd8; a_sign2 = 4'd4; a_sign3 = 4'd16;
b_sign0 = 4'd14; b_sign1 = 4'd7; b_sign2 = 4'd16; b_sign3 = 4'd15;
@(posedge clk_i);
a_mant0 = 8'd252; a_mant1 = 8'd59; a_mant2 = 8'd113; a_mant3 = 8'd93;
b_mant0 = 8'd221; b_mant1 = 8'd117; b_mant2 = 8'd124; b_mant3 = 8'd99;
a_exp0 = 10'd1005; a_exp1 = 10'd107; a_exp2 = 10'd10; a_exp3 = 10'd932;
b_exp0 = 10'd877; b_exp1 = 10'd277; b_exp2 = 10'd980; b_exp3 = 10'd512;
a_sign0 = 4'd6; a_sign1 = 4'd2; a_sign2 = 4'd14; a_sign3 = 4'd3;
b_sign0 = 4'd10; b_sign1 = 4'd4; b_sign2 = 4'd10; b_sign3 = 4'd1;
@(posedge clk_i);
a_mant0 = 8'd121; a_mant1 = 8'd170; a_mant2 = 8'd165; a_mant3 = 8'd5;
b_mant0 = 8'd36; b_mant1 = 8'd252; b_mant2 = 8'd61; b_mant3 = 8'd92;
a_exp0 = 10'd520; a_exp1 = 10'd68; a_exp2 = 10'd377; a_exp3 = 10'd32;
b_exp0 = 10'd468; b_exp1 = 10'd615; b_exp2 = 10'd376; b_exp3 = 10'd37;
a_sign0 = 4'd1; a_sign1 = 4'd8; a_sign2 = 4'd11; a_sign3 = 4'd8;
b_sign0 = 4'd12; b_sign1 = 4'd9; b_sign2 = 4'd0; b_sign3 = 4'd2;
@(posedge clk_i);
a_mant0 = 8'd198; a_mant1 = 8'd79; a_mant2 = 8'd234; a_mant3 = 8'd249;
b_mant0 = 8'd93; b_mant1 = 8'd56; b_mant2 = 8'd204; b_mant3 = 8'd32;
a_exp0 = 10'd307; a_exp1 = 10'd114; a_exp2 = 10'd868; a_exp3 = 10'd258;
b_exp0 = 10'd581; b_exp1 = 10'd727; b_exp2 = 10'd280; b_exp3 = 10'd250;
a_sign0 = 4'd7; a_sign1 = 4'd10; a_sign2 = 4'd10; a_sign3 = 4'd0;
b_sign0 = 4'd14; b_sign1 = 4'd8; b_sign2 = 4'd7; b_sign3 = 4'd8;
@(posedge clk_i);
a_mant0 = 8'd234; a_mant1 = 8'd214; a_mant2 = 8'd217; a_mant3 = 8'd6;
b_mant0 = 8'd243; b_mant1 = 8'd246; b_mant2 = 8'd141; b_mant3 = 8'd184;
a_exp0 = 10'd144; a_exp1 = 10'd215; a_exp2 = 10'd209; a_exp3 = 10'd543;
b_exp0 = 10'd126; b_exp1 = 10'd33; b_exp2 = 10'd1023; b_exp3 = 10'd869;
a_sign0 = 4'd2; a_sign1 = 4'd6; a_sign2 = 4'd6; a_sign3 = 4'd2;
b_sign0 = 4'd0; b_sign1 = 4'd11; b_sign2 = 4'd3; b_sign3 = 4'd12;
@(posedge clk_i);
shared_exps0 = 8'd136;
shared_exps1 = 8'd134;
rstn = 0;
@(posedge clk_i);
rstn = 1;
a_mant0 = 8'd212; a_mant1 = 8'd94; a_mant2 = 8'd148; a_mant3 = 8'd179;
b_mant0 = 8'd62; b_mant1 = 8'd200; b_mant2 = 8'd255; b_mant3 = 8'd216;
a_exp0 = 10'd436; a_exp1 = 10'd190; a_exp2 = 10'd1006; a_exp3 = 10'd93;
b_exp0 = 10'd107; b_exp1 = 10'd145; b_exp2 = 10'd202; b_exp3 = 10'd519;
a_sign0 = 4'd8; a_sign1 = 4'd6; a_sign2 = 4'd6; a_sign3 = 4'd14;
b_sign0 = 4'd15; b_sign1 = 4'd16; b_sign2 = 4'd1; b_sign3 = 4'd14;
@(posedge clk_i);
a_mant0 = 8'd229; a_mant1 = 8'd17; a_mant2 = 8'd139; a_mant3 = 8'd4;
b_mant0 = 8'd198; b_mant1 = 8'd29; b_mant2 = 8'd194; b_mant3 = 8'd253;
a_exp0 = 10'd330; a_exp1 = 10'd334; a_exp2 = 10'd451; a_exp3 = 10'd546;
b_exp0 = 10'd280; b_exp1 = 10'd967; b_exp2 = 10'd517; b_exp3 = 10'd911;
a_sign0 = 4'd1; a_sign1 = 4'd8; a_sign2 = 4'd6; a_sign3 = 4'd2;
b_sign0 = 4'd5; b_sign1 = 4'd1; b_sign2 = 4'd0; b_sign3 = 4'd0;
@(posedge clk_i);
a_mant0 = 8'd117; a_mant1 = 8'd75; a_mant2 = 8'd40; a_mant3 = 8'd30;
b_mant0 = 8'd37; b_mant1 = 8'd239; b_mant2 = 8'd56; b_mant3 = 8'd31;
a_exp0 = 10'd663; a_exp1 = 10'd948; a_exp2 = 10'd175; a_exp3 = 10'd598;
b_exp0 = 10'd511; b_exp1 = 10'd604; b_exp2 = 10'd591; b_exp3 = 10'd780;
a_sign0 = 4'd5; a_sign1 = 4'd11; a_sign2 = 4'd3; a_sign3 = 4'd13;
b_sign0 = 4'd14; b_sign1 = 4'd14; b_sign2 = 4'd0; b_sign3 = 4'd5;
@(posedge clk_i);
a_mant0 = 8'd38; a_mant1 = 8'd73; a_mant2 = 8'd152; a_mant3 = 8'd235;
b_mant0 = 8'd21; b_mant1 = 8'd45; b_mant2 = 8'd163; b_mant3 = 8'd49;
a_exp0 = 10'd81; a_exp1 = 10'd80; a_exp2 = 10'd955; a_exp3 = 10'd657;
b_exp0 = 10'd805; b_exp1 = 10'd69; b_exp2 = 10'd684; b_exp3 = 10'd626;
a_sign0 = 4'd11; a_sign1 = 4'd12; a_sign2 = 4'd11; a_sign3 = 4'd15;
b_sign0 = 4'd13; b_sign1 = 4'd11; b_sign2 = 4'd2; b_sign3 = 4'd6;
@(posedge clk_i);
a_mant0 = 8'd69; a_mant1 = 8'd118; a_mant2 = 8'd160; a_mant3 = 8'd232;
b_mant0 = 8'd34; b_mant1 = 8'd173; b_mant2 = 8'd153; b_mant3 = 8'd107;
a_exp0 = 10'd243; a_exp1 = 10'd65; a_exp2 = 10'd23; a_exp3 = 10'd609;
b_exp0 = 10'd674; b_exp1 = 10'd759; b_exp2 = 10'd974; b_exp3 = 10'd963;
a_sign0 = 4'd6; a_sign1 = 4'd3; a_sign2 = 4'd15; a_sign3 = 4'd12;
b_sign0 = 4'd13; b_sign1 = 4'd13; b_sign2 = 4'd6; b_sign3 = 4'd4;
@(posedge clk_i);
a_mant0 = 8'd31; a_mant1 = 8'd120; a_mant2 = 8'd6; a_mant3 = 8'd51;
b_mant0 = 8'd52; b_mant1 = 8'd15; b_mant2 = 8'd89; b_mant3 = 8'd203;
a_exp0 = 10'd163; a_exp1 = 10'd704; a_exp2 = 10'd887; a_exp3 = 10'd936;
b_exp0 = 10'd613; b_exp1 = 10'd382; b_exp2 = 10'd909; b_exp3 = 10'd862;
a_sign0 = 4'd7; a_sign1 = 4'd16; a_sign2 = 4'd4; a_sign3 = 4'd2;
b_sign0 = 4'd9; b_sign1 = 4'd4; b_sign2 = 4'd3; b_sign3 = 4'd5;
@(posedge clk_i);
a_mant0 = 8'd22; a_mant1 = 8'd62; a_mant2 = 8'd174; a_mant3 = 8'd202;
b_mant0 = 8'd232; b_mant1 = 8'd67; b_mant2 = 8'd11; b_mant3 = 8'd248;
a_exp0 = 10'd35; a_exp1 = 10'd238; a_exp2 = 10'd186; a_exp3 = 10'd531;
b_exp0 = 10'd921; b_exp1 = 10'd148; b_exp2 = 10'd442; b_exp3 = 10'd250;
a_sign0 = 4'd9; a_sign1 = 4'd6; a_sign2 = 4'd0; a_sign3 = 4'd13;
b_sign0 = 4'd8; b_sign1 = 4'd15; b_sign2 = 4'd3; b_sign3 = 4'd0;
@(posedge clk_i);
shared_exps0 = 8'd137;
shared_exps1 = 8'd138;
a_mant0 = 8'd162; a_mant1 = 8'd229; a_mant2 = 8'd87; a_mant3 = 8'd66;
b_mant0 = 8'd194; b_mant1 = 8'd139; b_mant2 = 8'd88; b_mant3 = 8'd238;
a_exp0 = 10'd12; a_exp1 = 10'd438; a_exp2 = 10'd878; a_exp3 = 10'd285;
b_exp0 = 10'd982; b_exp1 = 10'd515; b_exp2 = 10'd575; b_exp3 = 10'd855;
a_sign0 = 4'd16; a_sign1 = 4'd16; a_sign2 = 4'd4; a_sign3 = 4'd1;
b_sign0 = 4'd14; b_sign1 = 4'd0; b_sign2 = 4'd16; b_sign3 = 4'd3;
@(posedge clk_i);
a_mant0 = 8'd171; a_mant1 = 8'd124; a_mant2 = 8'd129; a_mant3 = 8'd66;
b_mant0 = 8'd145; b_mant1 = 8'd66; b_mant2 = 8'd194; b_mant3 = 8'd88;
a_exp0 = 10'd64; a_exp1 = 10'd913; a_exp2 = 10'd988; a_exp3 = 10'd98;
b_exp0 = 10'd879; b_exp1 = 10'd358; b_exp2 = 10'd274; b_exp3 = 10'd701;
a_sign0 = 4'd11; a_sign1 = 4'd7; a_sign2 = 4'd15; a_sign3 = 4'd11;
b_sign0 = 4'd5; b_sign1 = 4'd10; b_sign2 = 4'd16; b_sign3 = 4'd7;
@(posedge clk_i);
a_mant0 = 8'd223; a_mant1 = 8'd164; a_mant2 = 8'd57; a_mant3 = 8'd2;
b_mant0 = 8'd205; b_mant1 = 8'd155; b_mant2 = 8'd133; b_mant3 = 8'd184;
a_exp0 = 10'd602; a_exp1 = 10'd542; a_exp2 = 10'd676; a_exp3 = 10'd315;
b_exp0 = 10'd336; b_exp1 = 10'd908; b_exp2 = 10'd488; b_exp3 = 10'd741;
a_sign0 = 4'd11; a_sign1 = 4'd14; a_sign2 = 4'd3; a_sign3 = 4'd11;
b_sign0 = 4'd4; b_sign1 = 4'd15; b_sign2 = 4'd15; b_sign3 = 4'd9;
@(posedge clk_i);
a_mant0 = 8'd222; a_mant1 = 8'd255; a_mant2 = 8'd96; a_mant3 = 8'd78;
b_mant0 = 8'd208; b_mant1 = 8'd87; b_mant2 = 8'd126; b_mant3 = 8'd134;
a_exp0 = 10'd389; a_exp1 = 10'd686; a_exp2 = 10'd9; a_exp3 = 10'd626;
b_exp0 = 10'd219; b_exp1 = 10'd542; b_exp2 = 10'd366; b_exp3 = 10'd191;
a_sign0 = 4'd16; a_sign1 = 4'd12; a_sign2 = 4'd9; a_sign3 = 4'd2;
b_sign0 = 4'd16; b_sign1 = 4'd2; b_sign2 = 4'd14; b_sign3 = 4'd4;
@(posedge clk_i);
a_mant0 = 8'd220; a_mant1 = 8'd3; a_mant2 = 8'd37; a_mant3 = 8'd116;
b_mant0 = 8'd102; b_mant1 = 8'd67; b_mant2 = 8'd140; b_mant3 = 8'd156;
a_exp0 = 10'd272; a_exp1 = 10'd323; a_exp2 = 10'd876; a_exp3 = 10'd659;
b_exp0 = 10'd935; b_exp1 = 10'd267; b_exp2 = 10'd371; b_exp3 = 10'd881;
a_sign0 = 4'd1; a_sign1 = 4'd1; a_sign2 = 4'd15; a_sign3 = 4'd8;
b_sign0 = 4'd12; b_sign1 = 4'd3; b_sign2 = 4'd13; b_sign3 = 4'd1;
@(posedge clk_i);
a_mant0 = 8'd250; a_mant1 = 8'd6; a_mant2 = 8'd200; a_mant3 = 8'd4;
b_mant0 = 8'd238; b_mant1 = 8'd162; b_mant2 = 8'd59; b_mant3 = 8'd128;
a_exp0 = 10'd716; a_exp1 = 10'd375; a_exp2 = 10'd776; a_exp3 = 10'd924;
b_exp0 = 10'd476; b_exp1 = 10'd334; b_exp2 = 10'd876; b_exp3 = 10'd48;
a_sign0 = 4'd6; a_sign1 = 4'd1; a_sign2 = 4'd9; a_sign3 = 4'd10;
b_sign0 = 4'd7; b_sign1 = 4'd8; b_sign2 = 4'd10; b_sign3 = 4'd4;
@(posedge clk_i);
a_mant0 = 8'd163; a_mant1 = 8'd187; a_mant2 = 8'd227; a_mant3 = 8'd131;
b_mant0 = 8'd87; b_mant1 = 8'd85; b_mant2 = 8'd174; b_mant3 = 8'd82;
a_exp0 = 10'd968; a_exp1 = 10'd710; a_exp2 = 10'd906; a_exp3 = 10'd674;
b_exp0 = 10'd230; b_exp1 = 10'd810; b_exp2 = 10'd888; b_exp3 = 10'd459;
a_sign0 = 4'd12; a_sign1 = 4'd16; a_sign2 = 4'd13; a_sign3 = 4'd6;
b_sign0 = 4'd1; b_sign1 = 4'd16; b_sign2 = 4'd15; b_sign3 = 4'd10;
@(posedge clk_i);
a_mant0 = 8'd18; a_mant1 = 8'd139; a_mant2 = 8'd206; a_mant3 = 8'd238;
b_mant0 = 8'd24; b_mant1 = 8'd175; b_mant2 = 8'd73; b_mant3 = 8'd49;
a_exp0 = 10'd165; a_exp1 = 10'd375; a_exp2 = 10'd131; a_exp3 = 10'd867;
b_exp0 = 10'd455; b_exp1 = 10'd308; b_exp2 = 10'd671; b_exp3 = 10'd773;
a_sign0 = 4'd7; a_sign1 = 4'd0; a_sign2 = 4'd9; a_sign3 = 4'd5;
b_sign0 = 4'd11; b_sign1 = 4'd14; b_sign2 = 4'd8; b_sign3 = 4'd13;
@(posedge clk_i);
shared_exps0 = 8'd148;
shared_exps1 = 8'd120;
a_mant0 = 8'd55; a_mant1 = 8'd209; a_mant2 = 8'd227; a_mant3 = 8'd102;
b_mant0 = 8'd13; b_mant1 = 8'd135; b_mant2 = 8'd26; b_mant3 = 8'd107;
a_exp0 = 10'd25; a_exp1 = 10'd112; a_exp2 = 10'd732; a_exp3 = 10'd629;
b_exp0 = 10'd106; b_exp1 = 10'd680; b_exp2 = 10'd388; b_exp3 = 10'd990;
a_sign0 = 4'd3; a_sign1 = 4'd9; a_sign2 = 4'd3; a_sign3 = 4'd14;
b_sign0 = 4'd10; b_sign1 = 4'd12; b_sign2 = 4'd7; b_sign3 = 4'd14;
@(posedge clk_i);
a_mant0 = 8'd200; a_mant1 = 8'd39; a_mant2 = 8'd63; a_mant3 = 8'd191;
b_mant0 = 8'd75; b_mant1 = 8'd40; b_mant2 = 8'd219; b_mant3 = 8'd52;
a_exp0 = 10'd165; a_exp1 = 10'd595; a_exp2 = 10'd392; a_exp3 = 10'd1019;
b_exp0 = 10'd856; b_exp1 = 10'd656; b_exp2 = 10'd78; b_exp3 = 10'd203;
a_sign0 = 4'd0; a_sign1 = 4'd8; a_sign2 = 4'd2; a_sign3 = 4'd3;
b_sign0 = 4'd12; b_sign1 = 4'd12; b_sign2 = 4'd13; b_sign3 = 4'd10;
@(posedge clk_i);
a_mant0 = 8'd158; a_mant1 = 8'd98; a_mant2 = 8'd130; a_mant3 = 8'd114;
b_mant0 = 8'd54; b_mant1 = 8'd152; b_mant2 = 8'd9; b_mant3 = 8'd136;
a_exp0 = 10'd545; a_exp1 = 10'd70; a_exp2 = 10'd337; a_exp3 = 10'd890;
b_exp0 = 10'd494; b_exp1 = 10'd731; b_exp2 = 10'd2; b_exp3 = 10'd902;
a_sign0 = 4'd3; a_sign1 = 4'd3; a_sign2 = 4'd12; a_sign3 = 4'd4;
b_sign0 = 4'd14; b_sign1 = 4'd11; b_sign2 = 4'd6; b_sign3 = 4'd3;
@(posedge clk_i);
a_mant0 = 8'd247; a_mant1 = 8'd106; a_mant2 = 8'd173; a_mant3 = 8'd10;
b_mant0 = 8'd60; b_mant1 = 8'd209; b_mant2 = 8'd186; b_mant3 = 8'd106;
a_exp0 = 10'd964; a_exp1 = 10'd976; a_exp2 = 10'd379; a_exp3 = 10'd131;
b_exp0 = 10'd490; b_exp1 = 10'd965; b_exp2 = 10'd357; b_exp3 = 10'd938;
a_sign0 = 4'd0; a_sign1 = 4'd14; a_sign2 = 4'd1; a_sign3 = 4'd12;
b_sign0 = 4'd0; b_sign1 = 4'd12; b_sign2 = 4'd14; b_sign3 = 4'd16;
@(posedge clk_i);
a_mant0 = 8'd218; a_mant1 = 8'd68; a_mant2 = 8'd6; a_mant3 = 8'd6;
b_mant0 = 8'd193; b_mant1 = 8'd165; b_mant2 = 8'd41; b_mant3 = 8'd192;
a_exp0 = 10'd224; a_exp1 = 10'd716; a_exp2 = 10'd681; a_exp3 = 10'd69;
b_exp0 = 10'd831; b_exp1 = 10'd97; b_exp2 = 10'd581; b_exp3 = 10'd465;
a_sign0 = 4'd3; a_sign1 = 4'd14; a_sign2 = 4'd11; a_sign3 = 4'd2;
b_sign0 = 4'd16; b_sign1 = 4'd0; b_sign2 = 4'd13; b_sign3 = 4'd8;
@(posedge clk_i);
a_mant0 = 8'd172; a_mant1 = 8'd41; a_mant2 = 8'd105; a_mant3 = 8'd215;
b_mant0 = 8'd22; b_mant1 = 8'd52; b_mant2 = 8'd118; b_mant3 = 8'd171;
a_exp0 = 10'd241; a_exp1 = 10'd551; a_exp2 = 10'd905; a_exp3 = 10'd384;
b_exp0 = 10'd791; b_exp1 = 10'd824; b_exp2 = 10'd418; b_exp3 = 10'd65;
a_sign0 = 4'd3; a_sign1 = 4'd7; a_sign2 = 4'd13; a_sign3 = 4'd1;
b_sign0 = 4'd9; b_sign1 = 4'd15; b_sign2 = 4'd12; b_sign3 = 4'd7;
@(posedge clk_i);
a_mant0 = 8'd59; a_mant1 = 8'd207; a_mant2 = 8'd144; a_mant3 = 8'd190;
b_mant0 = 8'd171; b_mant1 = 8'd77; b_mant2 = 8'd126; b_mant3 = 8'd229;
a_exp0 = 10'd138; a_exp1 = 10'd142; a_exp2 = 10'd860; a_exp3 = 10'd104;
b_exp0 = 10'd476; b_exp1 = 10'd1019; b_exp2 = 10'd411; b_exp3 = 10'd21;
a_sign0 = 4'd0; a_sign1 = 4'd9; a_sign2 = 4'd3; a_sign3 = 4'd6;
b_sign0 = 4'd16; b_sign1 = 4'd3; b_sign2 = 4'd5; b_sign3 = 4'd10;
@(posedge clk_i);
a_mant0 = 8'd91; a_mant1 = 8'd73; a_mant2 = 8'd139; a_mant3 = 8'd193;
b_mant0 = 8'd110; b_mant1 = 8'd239; b_mant2 = 8'd191; b_mant3 = 8'd116;
a_exp0 = 10'd213; a_exp1 = 10'd513; a_exp2 = 10'd689; a_exp3 = 10'd547;
b_exp0 = 10'd289; b_exp1 = 10'd424; b_exp2 = 10'd580; b_exp3 = 10'd34;
a_sign0 = 4'd15; a_sign1 = 4'd3; a_sign2 = 4'd15; a_sign3 = 4'd4;
b_sign0 = 4'd12; b_sign1 = 4'd4; b_sign2 = 4'd6; b_sign3 = 4'd1;
@(posedge clk_i);
shared_exps0 = 8'd132;
shared_exps1 = 8'd120;
a_mant0 = 8'd141; a_mant1 = 8'd227; a_mant2 = 8'd133; a_mant3 = 8'd253;
b_mant0 = 8'd167; b_mant1 = 8'd15; b_mant2 = 8'd172; b_mant3 = 8'd180;
a_exp0 = 10'd956; a_exp1 = 10'd47; a_exp2 = 10'd238; a_exp3 = 10'd485;
b_exp0 = 10'd88; b_exp1 = 10'd840; b_exp2 = 10'd218; b_exp3 = 10'd357;
a_sign0 = 4'd14; a_sign1 = 4'd2; a_sign2 = 4'd0; a_sign3 = 4'd8;
b_sign0 = 4'd3; b_sign1 = 4'd16; b_sign2 = 4'd11; b_sign3 = 4'd5;
@(posedge clk_i);
a_mant0 = 8'd98; a_mant1 = 8'd241; a_mant2 = 8'd248; a_mant3 = 8'd203;
b_mant0 = 8'd217; b_mant1 = 8'd16; b_mant2 = 8'd167; b_mant3 = 8'd174;
a_exp0 = 10'd710; a_exp1 = 10'd926; a_exp2 = 10'd109; a_exp3 = 10'd416;
b_exp0 = 10'd197; b_exp1 = 10'd402; b_exp2 = 10'd274; b_exp3 = 10'd101;
a_sign0 = 4'd1; a_sign1 = 4'd5; a_sign2 = 4'd1; a_sign3 = 4'd14;
b_sign0 = 4'd6; b_sign1 = 4'd7; b_sign2 = 4'd9; b_sign3 = 4'd13;
@(posedge clk_i);
a_mant0 = 8'd143; a_mant1 = 8'd92; a_mant2 = 8'd169; a_mant3 = 8'd2;
b_mant0 = 8'd57; b_mant1 = 8'd129; b_mant2 = 8'd71; b_mant3 = 8'd230;
a_exp0 = 10'd143; a_exp1 = 10'd490; a_exp2 = 10'd642; a_exp3 = 10'd140;
b_exp0 = 10'd341; b_exp1 = 10'd953; b_exp2 = 10'd608; b_exp3 = 10'd58;
a_sign0 = 4'd0; a_sign1 = 4'd2; a_sign2 = 4'd4; a_sign3 = 4'd5;
b_sign0 = 4'd0; b_sign1 = 4'd10; b_sign2 = 4'd4; b_sign3 = 4'd8;
@(posedge clk_i);
a_mant0 = 8'd223; a_mant1 = 8'd143; a_mant2 = 8'd179; a_mant3 = 8'd243;
b_mant0 = 8'd69; b_mant1 = 8'd181; b_mant2 = 8'd175; b_mant3 = 8'd121;
a_exp0 = 10'd542; a_exp1 = 10'd609; a_exp2 = 10'd214; a_exp3 = 10'd212;
b_exp0 = 10'd930; b_exp1 = 10'd778; b_exp2 = 10'd814; b_exp3 = 10'd726;
a_sign0 = 4'd3; a_sign1 = 4'd8; a_sign2 = 4'd0; a_sign3 = 4'd13;
b_sign0 = 4'd3; b_sign1 = 4'd14; b_sign2 = 4'd12; b_sign3 = 4'd5;
@(posedge clk_i);
a_mant0 = 8'd194; a_mant1 = 8'd99; a_mant2 = 8'd109; a_mant3 = 8'd33;
b_mant0 = 8'd33; b_mant1 = 8'd191; b_mant2 = 8'd159; b_mant3 = 8'd9;
a_exp0 = 10'd311; a_exp1 = 10'd794; a_exp2 = 10'd49; a_exp3 = 10'd782;
b_exp0 = 10'd1013; b_exp1 = 10'd95; b_exp2 = 10'd488; b_exp3 = 10'd460;
a_sign0 = 4'd15; a_sign1 = 4'd12; a_sign2 = 4'd8; a_sign3 = 4'd16;
b_sign0 = 4'd12; b_sign1 = 4'd3; b_sign2 = 4'd13; b_sign3 = 4'd3;
@(posedge clk_i);
a_mant0 = 8'd214; a_mant1 = 8'd2; a_mant2 = 8'd54; a_mant3 = 8'd137;
b_mant0 = 8'd38; b_mant1 = 8'd98; b_mant2 = 8'd209; b_mant3 = 8'd133;
a_exp0 = 10'd861; a_exp1 = 10'd777; a_exp2 = 10'd18; a_exp3 = 10'd863;
b_exp0 = 10'd580; b_exp1 = 10'd743; b_exp2 = 10'd308; b_exp3 = 10'd50;
a_sign0 = 4'd7; a_sign1 = 4'd4; a_sign2 = 4'd2; a_sign3 = 4'd2;
b_sign0 = 4'd3; b_sign1 = 4'd1; b_sign2 = 4'd13; b_sign3 = 4'd4;
@(posedge clk_i);
a_mant0 = 8'd126; a_mant1 = 8'd14; a_mant2 = 8'd146; a_mant3 = 8'd217;
b_mant0 = 8'd68; b_mant1 = 8'd213; b_mant2 = 8'd193; b_mant3 = 8'd165;
a_exp0 = 10'd627; a_exp1 = 10'd483; a_exp2 = 10'd322; a_exp3 = 10'd723;
b_exp0 = 10'd859; b_exp1 = 10'd813; b_exp2 = 10'd420; b_exp3 = 10'd166;
a_sign0 = 4'd8; a_sign1 = 4'd2; a_sign2 = 4'd9; a_sign3 = 4'd10;
b_sign0 = 4'd8; b_sign1 = 4'd13; b_sign2 = 4'd4; b_sign3 = 4'd5;
@(posedge clk_i);
a_mant0 = 8'd220; a_mant1 = 8'd11; a_mant2 = 8'd239; a_mant3 = 8'd58;
b_mant0 = 8'd155; b_mant1 = 8'd196; b_mant2 = 8'd226; b_mant3 = 8'd169;
a_exp0 = 10'd594; a_exp1 = 10'd713; a_exp2 = 10'd401; a_exp3 = 10'd191;
b_exp0 = 10'd754; b_exp1 = 10'd485; b_exp2 = 10'd737; b_exp3 = 10'd667;
a_sign0 = 4'd2; a_sign1 = 4'd16; a_sign2 = 4'd15; a_sign3 = 4'd1;
b_sign0 = 4'd2; b_sign1 = 4'd13; b_sign2 = 4'd2; b_sign3 = 4'd3;
@(posedge clk_i);
shared_exps0 = 8'd147;
shared_exps1 = 8'd146;
rstn = 0;
@(posedge clk_i);
rstn = 1;
a_mant0 = 8'd169; a_mant1 = 8'd141; a_mant2 = 8'd14; a_mant3 = 8'd124;
b_mant0 = 8'd90; b_mant1 = 8'd35; b_mant2 = 8'd234; b_mant3 = 8'd215;
a_exp0 = 10'd85; a_exp1 = 10'd259; a_exp2 = 10'd347; a_exp3 = 10'd932;
b_exp0 = 10'd833; b_exp1 = 10'd372; b_exp2 = 10'd424; b_exp3 = 10'd457;
a_sign0 = 4'd6; a_sign1 = 4'd10; a_sign2 = 4'd3; a_sign3 = 4'd6;
b_sign0 = 4'd2; b_sign1 = 4'd16; b_sign2 = 4'd5; b_sign3 = 4'd10;
@(posedge clk_i);
a_mant0 = 8'd13; a_mant1 = 8'd219; a_mant2 = 8'd122; a_mant3 = 8'd173;
b_mant0 = 8'd118; b_mant1 = 8'd153; b_mant2 = 8'd231; b_mant3 = 8'd65;
a_exp0 = 10'd131; a_exp1 = 10'd902; a_exp2 = 10'd315; a_exp3 = 10'd518;
b_exp0 = 10'd30; b_exp1 = 10'd878; b_exp2 = 10'd716; b_exp3 = 10'd779;
a_sign0 = 4'd3; a_sign1 = 4'd14; a_sign2 = 4'd3; a_sign3 = 4'd4;
b_sign0 = 4'd12; b_sign1 = 4'd14; b_sign2 = 4'd10; b_sign3 = 4'd2;
@(posedge clk_i);
a_mant0 = 8'd58; a_mant1 = 8'd16; a_mant2 = 8'd251; a_mant3 = 8'd26;
b_mant0 = 8'd180; b_mant1 = 8'd116; b_mant2 = 8'd106; b_mant3 = 8'd105;
a_exp0 = 10'd688; a_exp1 = 10'd495; a_exp2 = 10'd417; a_exp3 = 10'd900;
b_exp0 = 10'd255; b_exp1 = 10'd110; b_exp2 = 10'd810; b_exp3 = 10'd739;
a_sign0 = 4'd1; a_sign1 = 4'd4; a_sign2 = 4'd5; a_sign3 = 4'd7;
b_sign0 = 4'd6; b_sign1 = 4'd0; b_sign2 = 4'd16; b_sign3 = 4'd11;
@(posedge clk_i);
a_mant0 = 8'd18; a_mant1 = 8'd174; a_mant2 = 8'd68; a_mant3 = 8'd230;
b_mant0 = 8'd72; b_mant1 = 8'd167; b_mant2 = 8'd112; b_mant3 = 8'd18;
a_exp0 = 10'd510; a_exp1 = 10'd701; a_exp2 = 10'd671; a_exp3 = 10'd548;
b_exp0 = 10'd35; b_exp1 = 10'd277; b_exp2 = 10'd512; b_exp3 = 10'd287;
a_sign0 = 4'd8; a_sign1 = 4'd2; a_sign2 = 4'd2; a_sign3 = 4'd0;
b_sign0 = 4'd0; b_sign1 = 4'd15; b_sign2 = 4'd6; b_sign3 = 4'd8;
@(posedge clk_i);
a_mant0 = 8'd184; a_mant1 = 8'd117; a_mant2 = 8'd140; a_mant3 = 8'd197;
b_mant0 = 8'd121; b_mant1 = 8'd222; b_mant2 = 8'd58; b_mant3 = 8'd221;
a_exp0 = 10'd925; a_exp1 = 10'd995; a_exp2 = 10'd1015; a_exp3 = 10'd47;
b_exp0 = 10'd314; b_exp1 = 10'd318; b_exp2 = 10'd670; b_exp3 = 10'd704;
a_sign0 = 4'd6; a_sign1 = 4'd3; a_sign2 = 4'd10; a_sign3 = 4'd2;
b_sign0 = 4'd2; b_sign1 = 4'd12; b_sign2 = 4'd3; b_sign3 = 4'd12;
@(posedge clk_i);
a_mant0 = 8'd189; a_mant1 = 8'd143; a_mant2 = 8'd81; a_mant3 = 8'd99;
b_mant0 = 8'd169; b_mant1 = 8'd234; b_mant2 = 8'd109; b_mant3 = 8'd64;
a_exp0 = 10'd682; a_exp1 = 10'd748; a_exp2 = 10'd220; a_exp3 = 10'd831;
b_exp0 = 10'd377; b_exp1 = 10'd824; b_exp2 = 10'd844; b_exp3 = 10'd970;
a_sign0 = 4'd14; a_sign1 = 4'd10; a_sign2 = 4'd13; a_sign3 = 4'd4;
b_sign0 = 4'd8; b_sign1 = 4'd11; b_sign2 = 4'd13; b_sign3 = 4'd8;
@(posedge clk_i);
a_mant0 = 8'd58; a_mant1 = 8'd74; a_mant2 = 8'd142; a_mant3 = 8'd249;
b_mant0 = 8'd225; b_mant1 = 8'd10; b_mant2 = 8'd100; b_mant3 = 8'd58;
a_exp0 = 10'd981; a_exp1 = 10'd397; a_exp2 = 10'd961; a_exp3 = 10'd720;
b_exp0 = 10'd788; b_exp1 = 10'd120; b_exp2 = 10'd237; b_exp3 = 10'd942;
a_sign0 = 4'd9; a_sign1 = 4'd10; a_sign2 = 4'd6; a_sign3 = 4'd1;
b_sign0 = 4'd5; b_sign1 = 4'd7; b_sign2 = 4'd6; b_sign3 = 4'd11;
@(posedge clk_i);
shared_exps0 = 8'd153;
shared_exps1 = 8'd97;
a_mant0 = 8'd2; a_mant1 = 8'd133; a_mant2 = 8'd82; a_mant3 = 8'd100;
b_mant0 = 8'd219; b_mant1 = 8'd41; b_mant2 = 8'd87; b_mant3 = 8'd233;
a_exp0 = 10'd396; a_exp1 = 10'd277; a_exp2 = 10'd873; a_exp3 = 10'd706;
b_exp0 = 10'd193; b_exp1 = 10'd811; b_exp2 = 10'd693; b_exp3 = 10'd447;
a_sign0 = 4'd9; a_sign1 = 4'd4; a_sign2 = 4'd1; a_sign3 = 4'd10;
b_sign0 = 4'd15; b_sign1 = 4'd15; b_sign2 = 4'd16; b_sign3 = 4'd10;
@(posedge clk_i);
a_mant0 = 8'd134; a_mant1 = 8'd127; a_mant2 = 8'd65; a_mant3 = 8'd177;
b_mant0 = 8'd26; b_mant1 = 8'd120; b_mant2 = 8'd92; b_mant3 = 8'd58;
a_exp0 = 10'd12; a_exp1 = 10'd235; a_exp2 = 10'd812; a_exp3 = 10'd445;
b_exp0 = 10'd275; b_exp1 = 10'd601; b_exp2 = 10'd584; b_exp3 = 10'd643;
a_sign0 = 4'd3; a_sign1 = 4'd0; a_sign2 = 4'd0; a_sign3 = 4'd13;
b_sign0 = 4'd3; b_sign1 = 4'd13; b_sign2 = 4'd3; b_sign3 = 4'd0;
@(posedge clk_i);
a_mant0 = 8'd209; a_mant1 = 8'd115; a_mant2 = 8'd61; a_mant3 = 8'd51;
b_mant0 = 8'd136; b_mant1 = 8'd204; b_mant2 = 8'd40; b_mant3 = 8'd159;
a_exp0 = 10'd2; a_exp1 = 10'd200; a_exp2 = 10'd572; a_exp3 = 10'd879;
b_exp0 = 10'd677; b_exp1 = 10'd309; b_exp2 = 10'd733; b_exp3 = 10'd717;
a_sign0 = 4'd9; a_sign1 = 4'd14; a_sign2 = 4'd11; a_sign3 = 4'd3;
b_sign0 = 4'd10; b_sign1 = 4'd4; b_sign2 = 4'd9; b_sign3 = 4'd8;
@(posedge clk_i);
a_mant0 = 8'd232; a_mant1 = 8'd8; a_mant2 = 8'd147; a_mant3 = 8'd151;
b_mant0 = 8'd217; b_mant1 = 8'd80; b_mant2 = 8'd214; b_mant3 = 8'd230;
a_exp0 = 10'd337; a_exp1 = 10'd680; a_exp2 = 10'd696; a_exp3 = 10'd36;
b_exp0 = 10'd896; b_exp1 = 10'd506; b_exp2 = 10'd125; b_exp3 = 10'd827;
a_sign0 = 4'd7; a_sign1 = 4'd0; a_sign2 = 4'd0; a_sign3 = 4'd3;
b_sign0 = 4'd6; b_sign1 = 4'd5; b_sign2 = 4'd11; b_sign3 = 4'd8;
@(posedge clk_i);
a_mant0 = 8'd230; a_mant1 = 8'd211; a_mant2 = 8'd127; a_mant3 = 8'd225;
b_mant0 = 8'd231; b_mant1 = 8'd95; b_mant2 = 8'd218; b_mant3 = 8'd83;
a_exp0 = 10'd781; a_exp1 = 10'd923; a_exp2 = 10'd933; a_exp3 = 10'd986;
b_exp0 = 10'd83; b_exp1 = 10'd922; b_exp2 = 10'd36; b_exp3 = 10'd467;
a_sign0 = 4'd6; a_sign1 = 4'd8; a_sign2 = 4'd16; a_sign3 = 4'd13;
b_sign0 = 4'd2; b_sign1 = 4'd3; b_sign2 = 4'd13; b_sign3 = 4'd1;
@(posedge clk_i);
a_mant0 = 8'd132; a_mant1 = 8'd236; a_mant2 = 8'd233; a_mant3 = 8'd25;
b_mant0 = 8'd192; b_mant1 = 8'd141; b_mant2 = 8'd200; b_mant3 = 8'd239;
a_exp0 = 10'd31; a_exp1 = 10'd781; a_exp2 = 10'd100; a_exp3 = 10'd540;
b_exp0 = 10'd485; b_exp1 = 10'd127; b_exp2 = 10'd328; b_exp3 = 10'd680;
a_sign0 = 4'd8; a_sign1 = 4'd9; a_sign2 = 4'd12; a_sign3 = 4'd4;
b_sign0 = 4'd1; b_sign1 = 4'd10; b_sign2 = 4'd3; b_sign3 = 4'd2;
@(posedge clk_i);
a_mant0 = 8'd138; a_mant1 = 8'd42; a_mant2 = 8'd1; a_mant3 = 8'd248;
b_mant0 = 8'd94; b_mant1 = 8'd49; b_mant2 = 8'd171; b_mant3 = 8'd172;
a_exp0 = 10'd459; a_exp1 = 10'd585; a_exp2 = 10'd76; a_exp3 = 10'd198;
b_exp0 = 10'd306; b_exp1 = 10'd1013; b_exp2 = 10'd894; b_exp3 = 10'd470;
a_sign0 = 4'd14; a_sign1 = 4'd11; a_sign2 = 4'd3; a_sign3 = 4'd8;
b_sign0 = 4'd1; b_sign1 = 4'd2; b_sign2 = 4'd11; b_sign3 = 4'd2;
@(posedge clk_i);
a_mant0 = 8'd42; a_mant1 = 8'd234; a_mant2 = 8'd185; a_mant3 = 8'd167;
b_mant0 = 8'd110; b_mant1 = 8'd11; b_mant2 = 8'd217; b_mant3 = 8'd49;
a_exp0 = 10'd258; a_exp1 = 10'd531; a_exp2 = 10'd818; a_exp3 = 10'd835;
b_exp0 = 10'd878; b_exp1 = 10'd235; b_exp2 = 10'd881; b_exp3 = 10'd441;
a_sign0 = 4'd11; a_sign1 = 4'd8; a_sign2 = 4'd11; a_sign3 = 4'd0;
b_sign0 = 4'd5; b_sign1 = 4'd2; b_sign2 = 4'd14; b_sign3 = 4'd15;
@(posedge clk_i);
shared_exps0 = 8'd113;
shared_exps1 = 8'd142;
a_mant0 = 8'd10; a_mant1 = 8'd195; a_mant2 = 8'd25; a_mant3 = 8'd249;
b_mant0 = 8'd4; b_mant1 = 8'd228; b_mant2 = 8'd117; b_mant3 = 8'd117;
a_exp0 = 10'd166; a_exp1 = 10'd814; a_exp2 = 10'd577; a_exp3 = 10'd684;
b_exp0 = 10'd126; b_exp1 = 10'd930; b_exp2 = 10'd920; b_exp3 = 10'd442;
a_sign0 = 4'd16; a_sign1 = 4'd10; a_sign2 = 4'd15; a_sign3 = 4'd2;
b_sign0 = 4'd9; b_sign1 = 4'd8; b_sign2 = 4'd11; b_sign3 = 4'd12;
@(posedge clk_i);
a_mant0 = 8'd78; a_mant1 = 8'd16; a_mant2 = 8'd36; a_mant3 = 8'd156;
b_mant0 = 8'd160; b_mant1 = 8'd189; b_mant2 = 8'd9; b_mant3 = 8'd222;
a_exp0 = 10'd741; a_exp1 = 10'd574; a_exp2 = 10'd375; a_exp3 = 10'd661;
b_exp0 = 10'd631; b_exp1 = 10'd343; b_exp2 = 10'd777; b_exp3 = 10'd307;
a_sign0 = 4'd13; a_sign1 = 4'd7; a_sign2 = 4'd4; a_sign3 = 4'd6;
b_sign0 = 4'd1; b_sign1 = 4'd8; b_sign2 = 4'd6; b_sign3 = 4'd9;
@(posedge clk_i);
a_mant0 = 8'd169; a_mant1 = 8'd139; a_mant2 = 8'd224; a_mant3 = 8'd154;
b_mant0 = 8'd23; b_mant1 = 8'd229; b_mant2 = 8'd122; b_mant3 = 8'd204;
a_exp0 = 10'd997; a_exp1 = 10'd22; a_exp2 = 10'd37; a_exp3 = 10'd437;
b_exp0 = 10'd821; b_exp1 = 10'd848; b_exp2 = 10'd743; b_exp3 = 10'd176;
a_sign0 = 4'd12; a_sign1 = 4'd13; a_sign2 = 4'd8; a_sign3 = 4'd1;
b_sign0 = 4'd15; b_sign1 = 4'd16; b_sign2 = 4'd2; b_sign3 = 4'd12;
@(posedge clk_i);
a_mant0 = 8'd219; a_mant1 = 8'd241; a_mant2 = 8'd231; a_mant3 = 8'd225;
b_mant0 = 8'd147; b_mant1 = 8'd109; b_mant2 = 8'd136; b_mant3 = 8'd156;
a_exp0 = 10'd112; a_exp1 = 10'd964; a_exp2 = 10'd879; a_exp3 = 10'd453;
b_exp0 = 10'd498; b_exp1 = 10'd822; b_exp2 = 10'd44; b_exp3 = 10'd892;
a_sign0 = 4'd4; a_sign1 = 4'd16; a_sign2 = 4'd5; a_sign3 = 4'd2;
b_sign0 = 4'd11; b_sign1 = 4'd9; b_sign2 = 4'd14; b_sign3 = 4'd13;
@(posedge clk_i);
a_mant0 = 8'd145; a_mant1 = 8'd248; a_mant2 = 8'd130; a_mant3 = 8'd253;
b_mant0 = 8'd153; b_mant1 = 8'd205; b_mant2 = 8'd187; b_mant3 = 8'd26;
a_exp0 = 10'd163; a_exp1 = 10'd95; a_exp2 = 10'd772; a_exp3 = 10'd163;
b_exp0 = 10'd60; b_exp1 = 10'd207; b_exp2 = 10'd824; b_exp3 = 10'd494;
a_sign0 = 4'd2; a_sign1 = 4'd6; a_sign2 = 4'd7; a_sign3 = 4'd7;
b_sign0 = 4'd7; b_sign1 = 4'd1; b_sign2 = 4'd8; b_sign3 = 4'd13;
@(posedge clk_i);
a_mant0 = 8'd155; a_mant1 = 8'd175; a_mant2 = 8'd5; a_mant3 = 8'd222;
b_mant0 = 8'd176; b_mant1 = 8'd157; b_mant2 = 8'd124; b_mant3 = 8'd4;
a_exp0 = 10'd990; a_exp1 = 10'd915; a_exp2 = 10'd484; a_exp3 = 10'd909;
b_exp0 = 10'd801; b_exp1 = 10'd1004; b_exp2 = 10'd691; b_exp3 = 10'd602;
a_sign0 = 4'd7; a_sign1 = 4'd10; a_sign2 = 4'd1; a_sign3 = 4'd15;
b_sign0 = 4'd11; b_sign1 = 4'd11; b_sign2 = 4'd13; b_sign3 = 4'd3;
@(posedge clk_i);
a_mant0 = 8'd159; a_mant1 = 8'd169; a_mant2 = 8'd121; a_mant3 = 8'd19;
b_mant0 = 8'd233; b_mant1 = 8'd246; b_mant2 = 8'd202; b_mant3 = 8'd111;
a_exp0 = 10'd479; a_exp1 = 10'd999; a_exp2 = 10'd592; a_exp3 = 10'd684;
b_exp0 = 10'd974; b_exp1 = 10'd366; b_exp2 = 10'd278; b_exp3 = 10'd904;
a_sign0 = 4'd0; a_sign1 = 4'd0; a_sign2 = 4'd9; a_sign3 = 4'd0;
b_sign0 = 4'd9; b_sign1 = 4'd12; b_sign2 = 4'd14; b_sign3 = 4'd16;
@(posedge clk_i);
a_mant0 = 8'd156; a_mant1 = 8'd188; a_mant2 = 8'd135; a_mant3 = 8'd111;
b_mant0 = 8'd168; b_mant1 = 8'd78; b_mant2 = 8'd180; b_mant3 = 8'd151;
a_exp0 = 10'd489; a_exp1 = 10'd826; a_exp2 = 10'd243; a_exp3 = 10'd620;
b_exp0 = 10'd509; b_exp1 = 10'd380; b_exp2 = 10'd102; b_exp3 = 10'd1015;
a_sign0 = 4'd11; a_sign1 = 4'd16; a_sign2 = 4'd4; a_sign3 = 4'd11;
b_sign0 = 4'd11; b_sign1 = 4'd4; b_sign2 = 4'd15; b_sign3 = 4'd14;
@(posedge clk_i);
shared_exps0 = 8'd124;
shared_exps1 = 8'd137;
a_mant0 = 8'd78; a_mant1 = 8'd7; a_mant2 = 8'd65; a_mant3 = 8'd120;
b_mant0 = 8'd73; b_mant1 = 8'd246; b_mant2 = 8'd92; b_mant3 = 8'd177;
a_exp0 = 10'd1010; a_exp1 = 10'd472; a_exp2 = 10'd126; a_exp3 = 10'd661;
b_exp0 = 10'd727; b_exp1 = 10'd518; b_exp2 = 10'd459; b_exp3 = 10'd97;
a_sign0 = 4'd7; a_sign1 = 4'd2; a_sign2 = 4'd10; a_sign3 = 4'd12;
b_sign0 = 4'd13; b_sign1 = 4'd2; b_sign2 = 4'd3; b_sign3 = 4'd4;
@(posedge clk_i);
a_mant0 = 8'd40; a_mant1 = 8'd114; a_mant2 = 8'd47; a_mant3 = 8'd35;
b_mant0 = 8'd175; b_mant1 = 8'd36; b_mant2 = 8'd195; b_mant3 = 8'd60;
a_exp0 = 10'd533; a_exp1 = 10'd314; a_exp2 = 10'd83; a_exp3 = 10'd568;
b_exp0 = 10'd507; b_exp1 = 10'd574; b_exp2 = 10'd328; b_exp3 = 10'd539;
a_sign0 = 4'd2; a_sign1 = 4'd16; a_sign2 = 4'd2; a_sign3 = 4'd12;
b_sign0 = 4'd3; b_sign1 = 4'd6; b_sign2 = 4'd14; b_sign3 = 4'd0;
@(posedge clk_i);
a_mant0 = 8'd166; a_mant1 = 8'd246; a_mant2 = 8'd123; a_mant3 = 8'd22;
b_mant0 = 8'd73; b_mant1 = 8'd31; b_mant2 = 8'd197; b_mant3 = 8'd167;
a_exp0 = 10'd836; a_exp1 = 10'd848; a_exp2 = 10'd25; a_exp3 = 10'd722;
b_exp0 = 10'd396; b_exp1 = 10'd323; b_exp2 = 10'd350; b_exp3 = 10'd172;
a_sign0 = 4'd16; a_sign1 = 4'd15; a_sign2 = 4'd1; a_sign3 = 4'd11;
b_sign0 = 4'd3; b_sign1 = 4'd13; b_sign2 = 4'd3; b_sign3 = 4'd6;
@(posedge clk_i);
a_mant0 = 8'd227; a_mant1 = 8'd52; a_mant2 = 8'd8; a_mant3 = 8'd171;
b_mant0 = 8'd141; b_mant1 = 8'd145; b_mant2 = 8'd132; b_mant3 = 8'd36;
a_exp0 = 10'd651; a_exp1 = 10'd200; a_exp2 = 10'd54; a_exp3 = 10'd24;
b_exp0 = 10'd197; b_exp1 = 10'd965; b_exp2 = 10'd601; b_exp3 = 10'd855;
a_sign0 = 4'd16; a_sign1 = 4'd6; a_sign2 = 4'd10; a_sign3 = 4'd10;
b_sign0 = 4'd16; b_sign1 = 4'd8; b_sign2 = 4'd11; b_sign3 = 4'd3;
@(posedge clk_i);
a_mant0 = 8'd86; a_mant1 = 8'd213; a_mant2 = 8'd8; a_mant3 = 8'd73;
b_mant0 = 8'd112; b_mant1 = 8'd134; b_mant2 = 8'd197; b_mant3 = 8'd84;
a_exp0 = 10'd15; a_exp1 = 10'd535; a_exp2 = 10'd936; a_exp3 = 10'd489;
b_exp0 = 10'd999; b_exp1 = 10'd19; b_exp2 = 10'd472; b_exp3 = 10'd659;
a_sign0 = 4'd1; a_sign1 = 4'd10; a_sign2 = 4'd8; a_sign3 = 4'd0;
b_sign0 = 4'd14; b_sign1 = 4'd1; b_sign2 = 4'd4; b_sign3 = 4'd7;
@(posedge clk_i);
a_mant0 = 8'd62; a_mant1 = 8'd239; a_mant2 = 8'd221; a_mant3 = 8'd168;
b_mant0 = 8'd94; b_mant1 = 8'd141; b_mant2 = 8'd216; b_mant3 = 8'd83;
a_exp0 = 10'd475; a_exp1 = 10'd131; a_exp2 = 10'd794; a_exp3 = 10'd674;
b_exp0 = 10'd156; b_exp1 = 10'd412; b_exp2 = 10'd629; b_exp3 = 10'd238;
a_sign0 = 4'd7; a_sign1 = 4'd5; a_sign2 = 4'd16; a_sign3 = 4'd1;
b_sign0 = 4'd6; b_sign1 = 4'd5; b_sign2 = 4'd6; b_sign3 = 4'd9;
@(posedge clk_i);
a_mant0 = 8'd141; a_mant1 = 8'd112; a_mant2 = 8'd215; a_mant3 = 8'd4;
b_mant0 = 8'd68; b_mant1 = 8'd62; b_mant2 = 8'd186; b_mant3 = 8'd44;
a_exp0 = 10'd708; a_exp1 = 10'd934; a_exp2 = 10'd552; a_exp3 = 10'd630;
b_exp0 = 10'd918; b_exp1 = 10'd804; b_exp2 = 10'd285; b_exp3 = 10'd716;
a_sign0 = 4'd7; a_sign1 = 4'd3; a_sign2 = 4'd3; a_sign3 = 4'd0;
b_sign0 = 4'd9; b_sign1 = 4'd4; b_sign2 = 4'd9; b_sign3 = 4'd5;
@(posedge clk_i);
a_mant0 = 8'd70; a_mant1 = 8'd146; a_mant2 = 8'd14; a_mant3 = 8'd54;
b_mant0 = 8'd148; b_mant1 = 8'd63; b_mant2 = 8'd44; b_mant3 = 8'd203;
a_exp0 = 10'd683; a_exp1 = 10'd332; a_exp2 = 10'd438; a_exp3 = 10'd282;
b_exp0 = 10'd534; b_exp1 = 10'd59; b_exp2 = 10'd807; b_exp3 = 10'd769;
a_sign0 = 4'd0; a_sign1 = 4'd10; a_sign2 = 4'd15; a_sign3 = 4'd7;
b_sign0 = 4'd12; b_sign1 = 4'd1; b_sign2 = 4'd11; b_sign3 = 4'd9;
@(posedge clk_i);
shared_exps0 = 8'd115;
shared_exps1 = 8'd129;
rstn = 0;
@(posedge clk_i);
rstn = 1;
a_mant0 = 8'd126; a_mant1 = 8'd172; a_mant2 = 8'd22; a_mant3 = 8'd202;
b_mant0 = 8'd238; b_mant1 = 8'd168; b_mant2 = 8'd213; b_mant3 = 8'd136;
a_exp0 = 10'd911; a_exp1 = 10'd698; a_exp2 = 10'd577; a_exp3 = 10'd224;
b_exp0 = 10'd387; b_exp1 = 10'd1014; b_exp2 = 10'd840; b_exp3 = 10'd164;
a_sign0 = 4'd0; a_sign1 = 4'd15; a_sign2 = 4'd15; a_sign3 = 4'd8;
b_sign0 = 4'd13; b_sign1 = 4'd9; b_sign2 = 4'd13; b_sign3 = 4'd5;
@(posedge clk_i);
a_mant0 = 8'd0; a_mant1 = 8'd191; a_mant2 = 8'd225; a_mant3 = 8'd237;
b_mant0 = 8'd226; b_mant1 = 8'd2; b_mant2 = 8'd24; b_mant3 = 8'd64;
a_exp0 = 10'd304; a_exp1 = 10'd204; a_exp2 = 10'd875; a_exp3 = 10'd502;
b_exp0 = 10'd3; b_exp1 = 10'd309; b_exp2 = 10'd574; b_exp3 = 10'd863;
a_sign0 = 4'd7; a_sign1 = 4'd13; a_sign2 = 4'd13; a_sign3 = 4'd12;
b_sign0 = 4'd2; b_sign1 = 4'd1; b_sign2 = 4'd2; b_sign3 = 4'd6;
@(posedge clk_i);
a_mant0 = 8'd23; a_mant1 = 8'd63; a_mant2 = 8'd141; a_mant3 = 8'd132;
b_mant0 = 8'd121; b_mant1 = 8'd160; b_mant2 = 8'd39; b_mant3 = 8'd54;
a_exp0 = 10'd391; a_exp1 = 10'd768; a_exp2 = 10'd491; a_exp3 = 10'd350;
b_exp0 = 10'd114; b_exp1 = 10'd659; b_exp2 = 10'd349; b_exp3 = 10'd326;
a_sign0 = 4'd9; a_sign1 = 4'd15; a_sign2 = 4'd9; a_sign3 = 4'd1;
b_sign0 = 4'd11; b_sign1 = 4'd15; b_sign2 = 4'd2; b_sign3 = 4'd5;
@(posedge clk_i);
a_mant0 = 8'd0; a_mant1 = 8'd24; a_mant2 = 8'd212; a_mant3 = 8'd136;
b_mant0 = 8'd175; b_mant1 = 8'd8; b_mant2 = 8'd87; b_mant3 = 8'd221;
a_exp0 = 10'd916; a_exp1 = 10'd185; a_exp2 = 10'd522; a_exp3 = 10'd0;
b_exp0 = 10'd59; b_exp1 = 10'd885; b_exp2 = 10'd37; b_exp3 = 10'd258;
a_sign0 = 4'd12; a_sign1 = 4'd16; a_sign2 = 4'd1; a_sign3 = 4'd0;
b_sign0 = 4'd8; b_sign1 = 4'd3; b_sign2 = 4'd10; b_sign3 = 4'd8;
@(posedge clk_i);
a_mant0 = 8'd15; a_mant1 = 8'd86; a_mant2 = 8'd254; a_mant3 = 8'd149;
b_mant0 = 8'd148; b_mant1 = 8'd238; b_mant2 = 8'd144; b_mant3 = 8'd35;
a_exp0 = 10'd749; a_exp1 = 10'd604; a_exp2 = 10'd998; a_exp3 = 10'd483;
b_exp0 = 10'd60; b_exp1 = 10'd904; b_exp2 = 10'd38; b_exp3 = 10'd933;
a_sign0 = 4'd15; a_sign1 = 4'd6; a_sign2 = 4'd6; a_sign3 = 4'd4;
b_sign0 = 4'd12; b_sign1 = 4'd3; b_sign2 = 4'd7; b_sign3 = 4'd12;
@(posedge clk_i);
a_mant0 = 8'd192; a_mant1 = 8'd174; a_mant2 = 8'd39; a_mant3 = 8'd45;
b_mant0 = 8'd92; b_mant1 = 8'd168; b_mant2 = 8'd141; b_mant3 = 8'd63;
a_exp0 = 10'd18; a_exp1 = 10'd725; a_exp2 = 10'd569; a_exp3 = 10'd823;
b_exp0 = 10'd872; b_exp1 = 10'd932; b_exp2 = 10'd128; b_exp3 = 10'd129;
a_sign0 = 4'd6; a_sign1 = 4'd3; a_sign2 = 4'd1; a_sign3 = 4'd3;
b_sign0 = 4'd5; b_sign1 = 4'd16; b_sign2 = 4'd0; b_sign3 = 4'd6;
@(posedge clk_i);
a_mant0 = 8'd42; a_mant1 = 8'd111; a_mant2 = 8'd120; a_mant3 = 8'd192;
b_mant0 = 8'd57; b_mant1 = 8'd152; b_mant2 = 8'd243; b_mant3 = 8'd136;
a_exp0 = 10'd588; a_exp1 = 10'd73; a_exp2 = 10'd326; a_exp3 = 10'd1007;
b_exp0 = 10'd854; b_exp1 = 10'd956; b_exp2 = 10'd725; b_exp3 = 10'd633;
a_sign0 = 4'd4; a_sign1 = 4'd11; a_sign2 = 4'd7; a_sign3 = 4'd5;
b_sign0 = 4'd9; b_sign1 = 4'd15; b_sign2 = 4'd13; b_sign3 = 4'd12;
@(posedge clk_i);
shared_exps0 = 8'd123;
shared_exps1 = 8'd125;
a_mant0 = 8'd89; a_mant1 = 8'd162; a_mant2 = 8'd81; a_mant3 = 8'd211;
b_mant0 = 8'd203; b_mant1 = 8'd187; b_mant2 = 8'd168; b_mant3 = 8'd198;
a_exp0 = 10'd582; a_exp1 = 10'd414; a_exp2 = 10'd831; a_exp3 = 10'd469;
b_exp0 = 10'd935; b_exp1 = 10'd815; b_exp2 = 10'd801; b_exp3 = 10'd624;
a_sign0 = 4'd5; a_sign1 = 4'd11; a_sign2 = 4'd0; a_sign3 = 4'd8;
b_sign0 = 4'd11; b_sign1 = 4'd9; b_sign2 = 4'd5; b_sign3 = 4'd8;
@(posedge clk_i);
a_mant0 = 8'd98; a_mant1 = 8'd171; a_mant2 = 8'd230; a_mant3 = 8'd214;
b_mant0 = 8'd131; b_mant1 = 8'd202; b_mant2 = 8'd38; b_mant3 = 8'd104;
a_exp0 = 10'd305; a_exp1 = 10'd975; a_exp2 = 10'd811; a_exp3 = 10'd746;
b_exp0 = 10'd383; b_exp1 = 10'd517; b_exp2 = 10'd655; b_exp3 = 10'd902;
a_sign0 = 4'd2; a_sign1 = 4'd5; a_sign2 = 4'd14; a_sign3 = 4'd15;
b_sign0 = 4'd6; b_sign1 = 4'd7; b_sign2 = 4'd13; b_sign3 = 4'd4;
@(posedge clk_i);
a_mant0 = 8'd31; a_mant1 = 8'd103; a_mant2 = 8'd100; a_mant3 = 8'd179;
b_mant0 = 8'd100; b_mant1 = 8'd140; b_mant2 = 8'd113; b_mant3 = 8'd27;
a_exp0 = 10'd246; a_exp1 = 10'd38; a_exp2 = 10'd82; a_exp3 = 10'd920;
b_exp0 = 10'd688; b_exp1 = 10'd873; b_exp2 = 10'd38; b_exp3 = 10'd697;
a_sign0 = 4'd8; a_sign1 = 4'd9; a_sign2 = 4'd0; a_sign3 = 4'd3;
b_sign0 = 4'd0; b_sign1 = 4'd9; b_sign2 = 4'd11; b_sign3 = 4'd11;
@(posedge clk_i);
a_mant0 = 8'd159; a_mant1 = 8'd150; a_mant2 = 8'd205; a_mant3 = 8'd61;
b_mant0 = 8'd200; b_mant1 = 8'd48; b_mant2 = 8'd182; b_mant3 = 8'd233;
a_exp0 = 10'd408; a_exp1 = 10'd878; a_exp2 = 10'd841; a_exp3 = 10'd999;
b_exp0 = 10'd316; b_exp1 = 10'd440; b_exp2 = 10'd196; b_exp3 = 10'd764;
a_sign0 = 4'd11; a_sign1 = 4'd5; a_sign2 = 4'd7; a_sign3 = 4'd8;
b_sign0 = 4'd9; b_sign1 = 4'd14; b_sign2 = 4'd13; b_sign3 = 4'd14;
@(posedge clk_i);
a_mant0 = 8'd243; a_mant1 = 8'd248; a_mant2 = 8'd139; a_mant3 = 8'd187;
b_mant0 = 8'd143; b_mant1 = 8'd14; b_mant2 = 8'd2; b_mant3 = 8'd74;
a_exp0 = 10'd430; a_exp1 = 10'd164; a_exp2 = 10'd50; a_exp3 = 10'd564;
b_exp0 = 10'd221; b_exp1 = 10'd321; b_exp2 = 10'd766; b_exp3 = 10'd845;
a_sign0 = 4'd9; a_sign1 = 4'd16; a_sign2 = 4'd10; a_sign3 = 4'd6;
b_sign0 = 4'd14; b_sign1 = 4'd0; b_sign2 = 4'd9; b_sign3 = 4'd1;
@(posedge clk_i);
a_mant0 = 8'd167; a_mant1 = 8'd70; a_mant2 = 8'd115; a_mant3 = 8'd49;
b_mant0 = 8'd28; b_mant1 = 8'd218; b_mant2 = 8'd80; b_mant3 = 8'd238;
a_exp0 = 10'd482; a_exp1 = 10'd241; a_exp2 = 10'd697; a_exp3 = 10'd559;
b_exp0 = 10'd656; b_exp1 = 10'd307; b_exp2 = 10'd89; b_exp3 = 10'd142;
a_sign0 = 4'd6; a_sign1 = 4'd12; a_sign2 = 4'd14; a_sign3 = 4'd9;
b_sign0 = 4'd5; b_sign1 = 4'd13; b_sign2 = 4'd7; b_sign3 = 4'd7;
@(posedge clk_i);
a_mant0 = 8'd241; a_mant1 = 8'd223; a_mant2 = 8'd227; a_mant3 = 8'd32;
b_mant0 = 8'd230; b_mant1 = 8'd85; b_mant2 = 8'd227; b_mant3 = 8'd35;
a_exp0 = 10'd271; a_exp1 = 10'd704; a_exp2 = 10'd858; a_exp3 = 10'd281;
b_exp0 = 10'd812; b_exp1 = 10'd396; b_exp2 = 10'd414; b_exp3 = 10'd482;
a_sign0 = 4'd15; a_sign1 = 4'd11; a_sign2 = 4'd10; a_sign3 = 4'd15;
b_sign0 = 4'd4; b_sign1 = 4'd16; b_sign2 = 4'd10; b_sign3 = 4'd11;
@(posedge clk_i);
a_mant0 = 8'd162; a_mant1 = 8'd117; a_mant2 = 8'd80; a_mant3 = 8'd249;
b_mant0 = 8'd241; b_mant1 = 8'd70; b_mant2 = 8'd122; b_mant3 = 8'd99;
a_exp0 = 10'd752; a_exp1 = 10'd293; a_exp2 = 10'd893; a_exp3 = 10'd927;
b_exp0 = 10'd494; b_exp1 = 10'd169; b_exp2 = 10'd448; b_exp3 = 10'd528;
a_sign0 = 4'd6; a_sign1 = 4'd2; a_sign2 = 4'd0; a_sign3 = 4'd10;
b_sign0 = 4'd5; b_sign1 = 4'd12; b_sign2 = 4'd4; b_sign3 = 4'd8;
@(posedge clk_i);
shared_exps0 = 8'd124;
shared_exps1 = 8'd124;
a_mant0 = 8'd191; a_mant1 = 8'd126; a_mant2 = 8'd208; a_mant3 = 8'd59;
b_mant0 = 8'd92; b_mant1 = 8'd209; b_mant2 = 8'd0; b_mant3 = 8'd253;
a_exp0 = 10'd321; a_exp1 = 10'd975; a_exp2 = 10'd270; a_exp3 = 10'd48;
b_exp0 = 10'd209; b_exp1 = 10'd201; b_exp2 = 10'd128; b_exp3 = 10'd634;
a_sign0 = 4'd4; a_sign1 = 4'd16; a_sign2 = 4'd12; a_sign3 = 4'd6;
b_sign0 = 4'd6; b_sign1 = 4'd7; b_sign2 = 4'd5; b_sign3 = 4'd2;
@(posedge clk_i);
a_mant0 = 8'd2; a_mant1 = 8'd183; a_mant2 = 8'd12; a_mant3 = 8'd24;
b_mant0 = 8'd229; b_mant1 = 8'd44; b_mant2 = 8'd28; b_mant3 = 8'd1;
a_exp0 = 10'd52; a_exp1 = 10'd739; a_exp2 = 10'd250; a_exp3 = 10'd76;
b_exp0 = 10'd714; b_exp1 = 10'd285; b_exp2 = 10'd789; b_exp3 = 10'd760;
a_sign0 = 4'd9; a_sign1 = 4'd12; a_sign2 = 4'd2; a_sign3 = 4'd8;
b_sign0 = 4'd11; b_sign1 = 4'd5; b_sign2 = 4'd7; b_sign3 = 4'd11;
@(posedge clk_i);
a_mant0 = 8'd152; a_mant1 = 8'd169; a_mant2 = 8'd245; a_mant3 = 8'd70;
b_mant0 = 8'd110; b_mant1 = 8'd238; b_mant2 = 8'd136; b_mant3 = 8'd237;
a_exp0 = 10'd24; a_exp1 = 10'd447; a_exp2 = 10'd709; a_exp3 = 10'd718;
b_exp0 = 10'd695; b_exp1 = 10'd460; b_exp2 = 10'd353; b_exp3 = 10'd623;
a_sign0 = 4'd9; a_sign1 = 4'd11; a_sign2 = 4'd3; a_sign3 = 4'd3;
b_sign0 = 4'd1; b_sign1 = 4'd14; b_sign2 = 4'd16; b_sign3 = 4'd13;
@(posedge clk_i);
a_mant0 = 8'd125; a_mant1 = 8'd144; a_mant2 = 8'd191; a_mant3 = 8'd37;
b_mant0 = 8'd154; b_mant1 = 8'd218; b_mant2 = 8'd144; b_mant3 = 8'd225;
a_exp0 = 10'd450; a_exp1 = 10'd484; a_exp2 = 10'd826; a_exp3 = 10'd693;
b_exp0 = 10'd119; b_exp1 = 10'd319; b_exp2 = 10'd16; b_exp3 = 10'd468;
a_sign0 = 4'd0; a_sign1 = 4'd11; a_sign2 = 4'd9; a_sign3 = 4'd0;
b_sign0 = 4'd12; b_sign1 = 4'd2; b_sign2 = 4'd0; b_sign3 = 4'd16;
@(posedge clk_i);
a_mant0 = 8'd164; a_mant1 = 8'd19; a_mant2 = 8'd86; a_mant3 = 8'd78;
b_mant0 = 8'd3; b_mant1 = 8'd187; b_mant2 = 8'd93; b_mant3 = 8'd172;
a_exp0 = 10'd962; a_exp1 = 10'd235; a_exp2 = 10'd312; a_exp3 = 10'd722;
b_exp0 = 10'd202; b_exp1 = 10'd80; b_exp2 = 10'd827; b_exp3 = 10'd321;
a_sign0 = 4'd0; a_sign1 = 4'd15; a_sign2 = 4'd5; a_sign3 = 4'd0;
b_sign0 = 4'd0; b_sign1 = 4'd6; b_sign2 = 4'd3; b_sign3 = 4'd14;
@(posedge clk_i);
a_mant0 = 8'd228; a_mant1 = 8'd128; a_mant2 = 8'd120; a_mant3 = 8'd127;
b_mant0 = 8'd161; b_mant1 = 8'd110; b_mant2 = 8'd194; b_mant3 = 8'd198;
a_exp0 = 10'd812; a_exp1 = 10'd12; a_exp2 = 10'd989; a_exp3 = 10'd50;
b_exp0 = 10'd466; b_exp1 = 10'd817; b_exp2 = 10'd366; b_exp3 = 10'd354;
a_sign0 = 4'd9; a_sign1 = 4'd7; a_sign2 = 4'd13; a_sign3 = 4'd10;
b_sign0 = 4'd9; b_sign1 = 4'd12; b_sign2 = 4'd2; b_sign3 = 4'd5;
@(posedge clk_i);
a_mant0 = 8'd139; a_mant1 = 8'd143; a_mant2 = 8'd238; a_mant3 = 8'd55;
b_mant0 = 8'd248; b_mant1 = 8'd154; b_mant2 = 8'd202; b_mant3 = 8'd154;
a_exp0 = 10'd720; a_exp1 = 10'd82; a_exp2 = 10'd242; a_exp3 = 10'd486;
b_exp0 = 10'd1002; b_exp1 = 10'd878; b_exp2 = 10'd809; b_exp3 = 10'd840;
a_sign0 = 4'd0; a_sign1 = 4'd16; a_sign2 = 4'd11; a_sign3 = 4'd9;
b_sign0 = 4'd7; b_sign1 = 4'd0; b_sign2 = 4'd9; b_sign3 = 4'd7;
@(posedge clk_i);
a_mant0 = 8'd142; a_mant1 = 8'd14; a_mant2 = 8'd120; a_mant3 = 8'd26;
b_mant0 = 8'd33; b_mant1 = 8'd19; b_mant2 = 8'd220; b_mant3 = 8'd147;
a_exp0 = 10'd1004; a_exp1 = 10'd538; a_exp2 = 10'd722; a_exp3 = 10'd1000;
b_exp0 = 10'd658; b_exp1 = 10'd651; b_exp2 = 10'd81; b_exp3 = 10'd192;
a_sign0 = 4'd7; a_sign1 = 4'd9; a_sign2 = 4'd14; a_sign3 = 4'd2;
b_sign0 = 4'd8; b_sign1 = 4'd13; b_sign2 = 4'd16; b_sign3 = 4'd10;
@(posedge clk_i);
shared_exps0 = 8'd139;
shared_exps1 = 8'd144;
a_mant0 = 8'd0; a_mant1 = 8'd42; a_mant2 = 8'd106; a_mant3 = 8'd87;
b_mant0 = 8'd221; b_mant1 = 8'd123; b_mant2 = 8'd57; b_mant3 = 8'd1;
a_exp0 = 10'd888; a_exp1 = 10'd497; a_exp2 = 10'd893; a_exp3 = 10'd908;
b_exp0 = 10'd283; b_exp1 = 10'd570; b_exp2 = 10'd1; b_exp3 = 10'd943;
a_sign0 = 4'd7; a_sign1 = 4'd3; a_sign2 = 4'd16; a_sign3 = 4'd7;
b_sign0 = 4'd8; b_sign1 = 4'd5; b_sign2 = 4'd15; b_sign3 = 4'd2;
@(posedge clk_i);
a_mant0 = 8'd142; a_mant1 = 8'd148; a_mant2 = 8'd4; a_mant3 = 8'd24;
b_mant0 = 8'd49; b_mant1 = 8'd181; b_mant2 = 8'd180; b_mant3 = 8'd238;
a_exp0 = 10'd767; a_exp1 = 10'd100; a_exp2 = 10'd211; a_exp3 = 10'd615;
b_exp0 = 10'd134; b_exp1 = 10'd380; b_exp2 = 10'd258; b_exp3 = 10'd495;
a_sign0 = 4'd13; a_sign1 = 4'd1; a_sign2 = 4'd4; a_sign3 = 4'd7;
b_sign0 = 4'd4; b_sign1 = 4'd9; b_sign2 = 4'd15; b_sign3 = 4'd3;
@(posedge clk_i);
a_mant0 = 8'd32; a_mant1 = 8'd94; a_mant2 = 8'd35; a_mant3 = 8'd16;
b_mant0 = 8'd22; b_mant1 = 8'd179; b_mant2 = 8'd210; b_mant3 = 8'd1;
a_exp0 = 10'd992; a_exp1 = 10'd803; a_exp2 = 10'd349; a_exp3 = 10'd209;
b_exp0 = 10'd314; b_exp1 = 10'd780; b_exp2 = 10'd910; b_exp3 = 10'd510;
a_sign0 = 4'd8; a_sign1 = 4'd8; a_sign2 = 4'd2; a_sign3 = 4'd8;
b_sign0 = 4'd9; b_sign1 = 4'd15; b_sign2 = 4'd12; b_sign3 = 4'd0;
@(posedge clk_i);
a_mant0 = 8'd84; a_mant1 = 8'd18; a_mant2 = 8'd199; a_mant3 = 8'd17;
b_mant0 = 8'd47; b_mant1 = 8'd98; b_mant2 = 8'd203; b_mant3 = 8'd64;
a_exp0 = 10'd556; a_exp1 = 10'd556; a_exp2 = 10'd356; a_exp3 = 10'd937;
b_exp0 = 10'd704; b_exp1 = 10'd157; b_exp2 = 10'd23; b_exp3 = 10'd456;
a_sign0 = 4'd13; a_sign1 = 4'd11; a_sign2 = 4'd2; a_sign3 = 4'd10;
b_sign0 = 4'd16; b_sign1 = 4'd4; b_sign2 = 4'd10; b_sign3 = 4'd2;
@(posedge clk_i);
a_mant0 = 8'd160; a_mant1 = 8'd157; a_mant2 = 8'd152; a_mant3 = 8'd103;
b_mant0 = 8'd7; b_mant1 = 8'd248; b_mant2 = 8'd105; b_mant3 = 8'd31;
a_exp0 = 10'd340; a_exp1 = 10'd942; a_exp2 = 10'd985; a_exp3 = 10'd891;
b_exp0 = 10'd570; b_exp1 = 10'd767; b_exp2 = 10'd14; b_exp3 = 10'd906;
a_sign0 = 4'd2; a_sign1 = 4'd15; a_sign2 = 4'd5; a_sign3 = 4'd13;
b_sign0 = 4'd3; b_sign1 = 4'd6; b_sign2 = 4'd1; b_sign3 = 4'd15;
@(posedge clk_i);
a_mant0 = 8'd39; a_mant1 = 8'd85; a_mant2 = 8'd135; a_mant3 = 8'd105;
b_mant0 = 8'd105; b_mant1 = 8'd157; b_mant2 = 8'd177; b_mant3 = 8'd102;
a_exp0 = 10'd288; a_exp1 = 10'd560; a_exp2 = 10'd116; a_exp3 = 10'd619;
b_exp0 = 10'd33; b_exp1 = 10'd938; b_exp2 = 10'd267; b_exp3 = 10'd700;
a_sign0 = 4'd12; a_sign1 = 4'd0; a_sign2 = 4'd4; a_sign3 = 4'd3;
b_sign0 = 4'd15; b_sign1 = 4'd3; b_sign2 = 4'd15; b_sign3 = 4'd11;
@(posedge clk_i);
a_mant0 = 8'd149; a_mant1 = 8'd138; a_mant2 = 8'd159; a_mant3 = 8'd131;
b_mant0 = 8'd41; b_mant1 = 8'd116; b_mant2 = 8'd137; b_mant3 = 8'd207;
a_exp0 = 10'd229; a_exp1 = 10'd841; a_exp2 = 10'd335; a_exp3 = 10'd697;
b_exp0 = 10'd820; b_exp1 = 10'd145; b_exp2 = 10'd24; b_exp3 = 10'd1005;
a_sign0 = 4'd2; a_sign1 = 4'd9; a_sign2 = 4'd2; a_sign3 = 4'd0;
b_sign0 = 4'd7; b_sign1 = 4'd15; b_sign2 = 4'd9; b_sign3 = 4'd15;
@(posedge clk_i);
a_mant0 = 8'd164; a_mant1 = 8'd197; a_mant2 = 8'd109; a_mant3 = 8'd134;
b_mant0 = 8'd146; b_mant1 = 8'd196; b_mant2 = 8'd68; b_mant3 = 8'd111;
a_exp0 = 10'd349; a_exp1 = 10'd103; a_exp2 = 10'd496; a_exp3 = 10'd906;
b_exp0 = 10'd937; b_exp1 = 10'd606; b_exp2 = 10'd11; b_exp3 = 10'd847;
a_sign0 = 4'd1; a_sign1 = 4'd4; a_sign2 = 4'd10; a_sign3 = 4'd16;
b_sign0 = 4'd15; b_sign1 = 4'd9; b_sign2 = 4'd14; b_sign3 = 4'd0;
@(posedge clk_i);
shared_exps0 = 8'd120;
shared_exps1 = 8'd129;
rstn = 0;
@(posedge clk_i);
rstn = 1;
a_mant0 = 8'd96; a_mant1 = 8'd225; a_mant2 = 8'd240; a_mant3 = 8'd14;
b_mant0 = 8'd36; b_mant1 = 8'd100; b_mant2 = 8'd61; b_mant3 = 8'd60;
a_exp0 = 10'd575; a_exp1 = 10'd605; a_exp2 = 10'd257; a_exp3 = 10'd357;
b_exp0 = 10'd541; b_exp1 = 10'd353; b_exp2 = 10'd967; b_exp3 = 10'd1018;
a_sign0 = 4'd9; a_sign1 = 4'd12; a_sign2 = 4'd9; a_sign3 = 4'd13;
b_sign0 = 4'd11; b_sign1 = 4'd6; b_sign2 = 4'd14; b_sign3 = 4'd7;
@(posedge clk_i);
a_mant0 = 8'd250; a_mant1 = 8'd233; a_mant2 = 8'd133; a_mant3 = 8'd239;
b_mant0 = 8'd254; b_mant1 = 8'd24; b_mant2 = 8'd211; b_mant3 = 8'd41;
a_exp0 = 10'd205; a_exp1 = 10'd684; a_exp2 = 10'd29; a_exp3 = 10'd186;
b_exp0 = 10'd507; b_exp1 = 10'd688; b_exp2 = 10'd115; b_exp3 = 10'd404;
a_sign0 = 4'd5; a_sign1 = 4'd7; a_sign2 = 4'd0; a_sign3 = 4'd14;
b_sign0 = 4'd12; b_sign1 = 4'd0; b_sign2 = 4'd7; b_sign3 = 4'd0;
@(posedge clk_i);
a_mant0 = 8'd145; a_mant1 = 8'd33; a_mant2 = 8'd9; a_mant3 = 8'd111;
b_mant0 = 8'd61; b_mant1 = 8'd217; b_mant2 = 8'd253; b_mant3 = 8'd128;
a_exp0 = 10'd330; a_exp1 = 10'd65; a_exp2 = 10'd227; a_exp3 = 10'd812;
b_exp0 = 10'd635; b_exp1 = 10'd481; b_exp2 = 10'd708; b_exp3 = 10'd275;
a_sign0 = 4'd15; a_sign1 = 4'd15; a_sign2 = 4'd15; a_sign3 = 4'd11;
b_sign0 = 4'd11; b_sign1 = 4'd10; b_sign2 = 4'd7; b_sign3 = 4'd2;
@(posedge clk_i);
a_mant0 = 8'd22; a_mant1 = 8'd3; a_mant2 = 8'd86; a_mant3 = 8'd97;
b_mant0 = 8'd3; b_mant1 = 8'd94; b_mant2 = 8'd89; b_mant3 = 8'd70;
a_exp0 = 10'd798; a_exp1 = 10'd824; a_exp2 = 10'd610; a_exp3 = 10'd308;
b_exp0 = 10'd1000; b_exp1 = 10'd520; b_exp2 = 10'd263; b_exp3 = 10'd976;
a_sign0 = 4'd2; a_sign1 = 4'd12; a_sign2 = 4'd5; a_sign3 = 4'd9;
b_sign0 = 4'd10; b_sign1 = 4'd13; b_sign2 = 4'd8; b_sign3 = 4'd2;
@(posedge clk_i);
a_mant0 = 8'd49; a_mant1 = 8'd158; a_mant2 = 8'd210; a_mant3 = 8'd102;
b_mant0 = 8'd203; b_mant1 = 8'd61; b_mant2 = 8'd109; b_mant3 = 8'd232;
a_exp0 = 10'd376; a_exp1 = 10'd528; a_exp2 = 10'd517; a_exp3 = 10'd793;
b_exp0 = 10'd247; b_exp1 = 10'd585; b_exp2 = 10'd631; b_exp3 = 10'd76;
a_sign0 = 4'd4; a_sign1 = 4'd6; a_sign2 = 4'd1; a_sign3 = 4'd8;
b_sign0 = 4'd0; b_sign1 = 4'd0; b_sign2 = 4'd15; b_sign3 = 4'd10;
@(posedge clk_i);
a_mant0 = 8'd0; a_mant1 = 8'd15; a_mant2 = 8'd247; a_mant3 = 8'd211;
b_mant0 = 8'd136; b_mant1 = 8'd197; b_mant2 = 8'd80; b_mant3 = 8'd44;
a_exp0 = 10'd122; a_exp1 = 10'd887; a_exp2 = 10'd210; a_exp3 = 10'd931;
b_exp0 = 10'd248; b_exp1 = 10'd471; b_exp2 = 10'd872; b_exp3 = 10'd353;
a_sign0 = 4'd10; a_sign1 = 4'd11; a_sign2 = 4'd13; a_sign3 = 4'd6;
b_sign0 = 4'd6; b_sign1 = 4'd15; b_sign2 = 4'd12; b_sign3 = 4'd8;
@(posedge clk_i);
a_mant0 = 8'd39; a_mant1 = 8'd34; a_mant2 = 8'd239; a_mant3 = 8'd221;
b_mant0 = 8'd85; b_mant1 = 8'd178; b_mant2 = 8'd99; b_mant3 = 8'd88;
a_exp0 = 10'd384; a_exp1 = 10'd682; a_exp2 = 10'd519; a_exp3 = 10'd561;
b_exp0 = 10'd702; b_exp1 = 10'd647; b_exp2 = 10'd869; b_exp3 = 10'd778;
a_sign0 = 4'd13; a_sign1 = 4'd1; a_sign2 = 4'd14; a_sign3 = 4'd13;
b_sign0 = 4'd5; b_sign1 = 4'd1; b_sign2 = 4'd12; b_sign3 = 4'd7;
@(posedge clk_i);
shared_exps0 = 8'd108;
shared_exps1 = 8'd143;
a_mant0 = 8'd47; a_mant1 = 8'd97; a_mant2 = 8'd55; a_mant3 = 8'd138;
b_mant0 = 8'd147; b_mant1 = 8'd224; b_mant2 = 8'd91; b_mant3 = 8'd197;
a_exp0 = 10'd1005; a_exp1 = 10'd359; a_exp2 = 10'd93; a_exp3 = 10'd673;
b_exp0 = 10'd211; b_exp1 = 10'd2; b_exp2 = 10'd434; b_exp3 = 10'd944;
a_sign0 = 4'd1; a_sign1 = 4'd14; a_sign2 = 4'd3; a_sign3 = 4'd10;
b_sign0 = 4'd10; b_sign1 = 4'd4; b_sign2 = 4'd6; b_sign3 = 4'd9;
@(posedge clk_i);
a_mant0 = 8'd93; a_mant1 = 8'd177; a_mant2 = 8'd24; a_mant3 = 8'd134;
b_mant0 = 8'd252; b_mant1 = 8'd144; b_mant2 = 8'd83; b_mant3 = 8'd119;
a_exp0 = 10'd12; a_exp1 = 10'd802; a_exp2 = 10'd167; a_exp3 = 10'd285;
b_exp0 = 10'd1014; b_exp1 = 10'd197; b_exp2 = 10'd966; b_exp3 = 10'd477;
a_sign0 = 4'd9; a_sign1 = 4'd1; a_sign2 = 4'd1; a_sign3 = 4'd3;
b_sign0 = 4'd11; b_sign1 = 4'd8; b_sign2 = 4'd8; b_sign3 = 4'd15;
@(posedge clk_i);
a_mant0 = 8'd245; a_mant1 = 8'd156; a_mant2 = 8'd205; a_mant3 = 8'd153;
b_mant0 = 8'd91; b_mant1 = 8'd53; b_mant2 = 8'd0; b_mant3 = 8'd215;
a_exp0 = 10'd494; a_exp1 = 10'd397; a_exp2 = 10'd880; a_exp3 = 10'd75;
b_exp0 = 10'd427; b_exp1 = 10'd93; b_exp2 = 10'd818; b_exp3 = 10'd620;
a_sign0 = 4'd0; a_sign1 = 4'd10; a_sign2 = 4'd7; a_sign3 = 4'd2;
b_sign0 = 4'd0; b_sign1 = 4'd11; b_sign2 = 4'd0; b_sign3 = 4'd14;
@(posedge clk_i);
a_mant0 = 8'd166; a_mant1 = 8'd171; a_mant2 = 8'd3; a_mant3 = 8'd58;
b_mant0 = 8'd239; b_mant1 = 8'd72; b_mant2 = 8'd182; b_mant3 = 8'd10;
a_exp0 = 10'd667; a_exp1 = 10'd837; a_exp2 = 10'd298; a_exp3 = 10'd896;
b_exp0 = 10'd1004; b_exp1 = 10'd396; b_exp2 = 10'd93; b_exp3 = 10'd450;
a_sign0 = 4'd13; a_sign1 = 4'd7; a_sign2 = 4'd8; a_sign3 = 4'd15;
b_sign0 = 4'd0; b_sign1 = 4'd11; b_sign2 = 4'd1; b_sign3 = 4'd12;
@(posedge clk_i);
a_mant0 = 8'd229; a_mant1 = 8'd218; a_mant2 = 8'd147; a_mant3 = 8'd124;
b_mant0 = 8'd111; b_mant1 = 8'd146; b_mant2 = 8'd247; b_mant3 = 8'd19;
a_exp0 = 10'd873; a_exp1 = 10'd134; a_exp2 = 10'd98; a_exp3 = 10'd844;
b_exp0 = 10'd579; b_exp1 = 10'd847; b_exp2 = 10'd870; b_exp3 = 10'd823;
a_sign0 = 4'd14; a_sign1 = 4'd6; a_sign2 = 4'd0; a_sign3 = 4'd4;
b_sign0 = 4'd0; b_sign1 = 4'd9; b_sign2 = 4'd16; b_sign3 = 4'd10;
@(posedge clk_i);
a_mant0 = 8'd143; a_mant1 = 8'd228; a_mant2 = 8'd236; a_mant3 = 8'd163;
b_mant0 = 8'd177; b_mant1 = 8'd33; b_mant2 = 8'd66; b_mant3 = 8'd234;
a_exp0 = 10'd170; a_exp1 = 10'd103; a_exp2 = 10'd971; a_exp3 = 10'd254;
b_exp0 = 10'd545; b_exp1 = 10'd1023; b_exp2 = 10'd550; b_exp3 = 10'd901;
a_sign0 = 4'd16; a_sign1 = 4'd9; a_sign2 = 4'd11; a_sign3 = 4'd8;
b_sign0 = 4'd5; b_sign1 = 4'd5; b_sign2 = 4'd0; b_sign3 = 4'd8;
@(posedge clk_i);
a_mant0 = 8'd53; a_mant1 = 8'd183; a_mant2 = 8'd30; a_mant3 = 8'd7;
b_mant0 = 8'd133; b_mant1 = 8'd216; b_mant2 = 8'd136; b_mant3 = 8'd187;
a_exp0 = 10'd359; a_exp1 = 10'd953; a_exp2 = 10'd813; a_exp3 = 10'd181;
b_exp0 = 10'd1011; b_exp1 = 10'd647; b_exp2 = 10'd898; b_exp3 = 10'd801;
a_sign0 = 4'd13; a_sign1 = 4'd14; a_sign2 = 4'd1; a_sign3 = 4'd3;
b_sign0 = 4'd13; b_sign1 = 4'd8; b_sign2 = 4'd3; b_sign3 = 4'd7;
@(posedge clk_i);
a_mant0 = 8'd27; a_mant1 = 8'd78; a_mant2 = 8'd71; a_mant3 = 8'd213;
b_mant0 = 8'd130; b_mant1 = 8'd96; b_mant2 = 8'd99; b_mant3 = 8'd230;
a_exp0 = 10'd700; a_exp1 = 10'd229; a_exp2 = 10'd508; a_exp3 = 10'd846;
b_exp0 = 10'd332; b_exp1 = 10'd712; b_exp2 = 10'd198; b_exp3 = 10'd496;
a_sign0 = 4'd16; a_sign1 = 4'd6; a_sign2 = 4'd0; a_sign3 = 4'd9;
b_sign0 = 4'd11; b_sign1 = 4'd12; b_sign2 = 4'd16; b_sign3 = 4'd10;
@(posedge clk_i);
shared_exps0 = 8'd94;
shared_exps1 = 8'd137;
a_mant0 = 8'd99; a_mant1 = 8'd120; a_mant2 = 8'd15; a_mant3 = 8'd209;
b_mant0 = 8'd141; b_mant1 = 8'd54; b_mant2 = 8'd105; b_mant3 = 8'd177;
a_exp0 = 10'd542; a_exp1 = 10'd883; a_exp2 = 10'd617; a_exp3 = 10'd91;
b_exp0 = 10'd577; b_exp1 = 10'd153; b_exp2 = 10'd374; b_exp3 = 10'd135;
a_sign0 = 4'd14; a_sign1 = 4'd12; a_sign2 = 4'd3; a_sign3 = 4'd0;
b_sign0 = 4'd5; b_sign1 = 4'd3; b_sign2 = 4'd14; b_sign3 = 4'd5;
@(posedge clk_i);
a_mant0 = 8'd107; a_mant1 = 8'd219; a_mant2 = 8'd75; a_mant3 = 8'd96;
b_mant0 = 8'd156; b_mant1 = 8'd37; b_mant2 = 8'd81; b_mant3 = 8'd10;
a_exp0 = 10'd132; a_exp1 = 10'd124; a_exp2 = 10'd830; a_exp3 = 10'd97;
b_exp0 = 10'd575; b_exp1 = 10'd61; b_exp2 = 10'd536; b_exp3 = 10'd82;
a_sign0 = 4'd16; a_sign1 = 4'd9; a_sign2 = 4'd6; a_sign3 = 4'd2;
b_sign0 = 4'd15; b_sign1 = 4'd4; b_sign2 = 4'd8; b_sign3 = 4'd5;
@(posedge clk_i);
a_mant0 = 8'd110; a_mant1 = 8'd8; a_mant2 = 8'd28; a_mant3 = 8'd61;
b_mant0 = 8'd241; b_mant1 = 8'd89; b_mant2 = 8'd235; b_mant3 = 8'd225;
a_exp0 = 10'd732; a_exp1 = 10'd28; a_exp2 = 10'd1022; a_exp3 = 10'd929;
b_exp0 = 10'd338; b_exp1 = 10'd668; b_exp2 = 10'd489; b_exp3 = 10'd122;
a_sign0 = 4'd12; a_sign1 = 4'd10; a_sign2 = 4'd5; a_sign3 = 4'd0;
b_sign0 = 4'd12; b_sign1 = 4'd13; b_sign2 = 4'd11; b_sign3 = 4'd9;
@(posedge clk_i);
a_mant0 = 8'd65; a_mant1 = 8'd170; a_mant2 = 8'd21; a_mant3 = 8'd110;
b_mant0 = 8'd59; b_mant1 = 8'd110; b_mant2 = 8'd9; b_mant3 = 8'd199;
a_exp0 = 10'd449; a_exp1 = 10'd386; a_exp2 = 10'd147; a_exp3 = 10'd965;
b_exp0 = 10'd533; b_exp1 = 10'd47; b_exp2 = 10'd606; b_exp3 = 10'd1010;
a_sign0 = 4'd11; a_sign1 = 4'd2; a_sign2 = 4'd2; a_sign3 = 4'd6;
b_sign0 = 4'd3; b_sign1 = 4'd15; b_sign2 = 4'd6; b_sign3 = 4'd14;
@(posedge clk_i);
a_mant0 = 8'd210; a_mant1 = 8'd17; a_mant2 = 8'd5; a_mant3 = 8'd76;
b_mant0 = 8'd233; b_mant1 = 8'd88; b_mant2 = 8'd129; b_mant3 = 8'd238;
a_exp0 = 10'd849; a_exp1 = 10'd496; a_exp2 = 10'd408; a_exp3 = 10'd704;
b_exp0 = 10'd323; b_exp1 = 10'd146; b_exp2 = 10'd252; b_exp3 = 10'd686;
a_sign0 = 4'd15; a_sign1 = 4'd13; a_sign2 = 4'd6; a_sign3 = 4'd15;
b_sign0 = 4'd3; b_sign1 = 4'd10; b_sign2 = 4'd6; b_sign3 = 4'd0;
@(posedge clk_i);
a_mant0 = 8'd85; a_mant1 = 8'd187; a_mant2 = 8'd182; a_mant3 = 8'd109;
b_mant0 = 8'd253; b_mant1 = 8'd170; b_mant2 = 8'd243; b_mant3 = 8'd32;
a_exp0 = 10'd97; a_exp1 = 10'd1004; a_exp2 = 10'd934; a_exp3 = 10'd331;
b_exp0 = 10'd60; b_exp1 = 10'd822; b_exp2 = 10'd385; b_exp3 = 10'd411;
a_sign0 = 4'd5; a_sign1 = 4'd5; a_sign2 = 4'd14; a_sign3 = 4'd14;
b_sign0 = 4'd12; b_sign1 = 4'd4; b_sign2 = 4'd0; b_sign3 = 4'd12;
@(posedge clk_i);
a_mant0 = 8'd195; a_mant1 = 8'd248; a_mant2 = 8'd33; a_mant3 = 8'd96;
b_mant0 = 8'd175; b_mant1 = 8'd244; b_mant2 = 8'd124; b_mant3 = 8'd94;
a_exp0 = 10'd267; a_exp1 = 10'd787; a_exp2 = 10'd942; a_exp3 = 10'd612;
b_exp0 = 10'd770; b_exp1 = 10'd1005; b_exp2 = 10'd907; b_exp3 = 10'd350;
a_sign0 = 4'd10; a_sign1 = 4'd15; a_sign2 = 4'd10; a_sign3 = 4'd1;
b_sign0 = 4'd10; b_sign1 = 4'd3; b_sign2 = 4'd1; b_sign3 = 4'd8;
@(posedge clk_i);
a_mant0 = 8'd137; a_mant1 = 8'd243; a_mant2 = 8'd240; a_mant3 = 8'd24;
b_mant0 = 8'd254; b_mant1 = 8'd134; b_mant2 = 8'd48; b_mant3 = 8'd75;
a_exp0 = 10'd173; a_exp1 = 10'd330; a_exp2 = 10'd977; a_exp3 = 10'd855;
b_exp0 = 10'd492; b_exp1 = 10'd338; b_exp2 = 10'd57; b_exp3 = 10'd223;
a_sign0 = 4'd12; a_sign1 = 4'd1; a_sign2 = 4'd11; a_sign3 = 4'd5;
b_sign0 = 4'd11; b_sign1 = 4'd14; b_sign2 = 4'd6; b_sign3 = 4'd1;
@(posedge clk_i);
shared_exps0 = 8'd103;
shared_exps1 = 8'd113;
a_mant0 = 8'd132; a_mant1 = 8'd222; a_mant2 = 8'd41; a_mant3 = 8'd100;
b_mant0 = 8'd107; b_mant1 = 8'd47; b_mant2 = 8'd129; b_mant3 = 8'd132;
a_exp0 = 10'd972; a_exp1 = 10'd746; a_exp2 = 10'd824; a_exp3 = 10'd963;
b_exp0 = 10'd685; b_exp1 = 10'd399; b_exp2 = 10'd906; b_exp3 = 10'd183;
a_sign0 = 4'd5; a_sign1 = 4'd0; a_sign2 = 4'd7; a_sign3 = 4'd9;
b_sign0 = 4'd14; b_sign1 = 4'd12; b_sign2 = 4'd0; b_sign3 = 4'd8;
@(posedge clk_i);
a_mant0 = 8'd189; a_mant1 = 8'd155; a_mant2 = 8'd89; a_mant3 = 8'd170;
b_mant0 = 8'd13; b_mant1 = 8'd25; b_mant2 = 8'd139; b_mant3 = 8'd179;
a_exp0 = 10'd192; a_exp1 = 10'd249; a_exp2 = 10'd164; a_exp3 = 10'd694;
b_exp0 = 10'd316; b_exp1 = 10'd908; b_exp2 = 10'd913; b_exp3 = 10'd18;
a_sign0 = 4'd15; a_sign1 = 4'd9; a_sign2 = 4'd7; a_sign3 = 4'd4;
b_sign0 = 4'd13; b_sign1 = 4'd0; b_sign2 = 4'd4; b_sign3 = 4'd8;
@(posedge clk_i);
a_mant0 = 8'd110; a_mant1 = 8'd24; a_mant2 = 8'd98; a_mant3 = 8'd127;
b_mant0 = 8'd55; b_mant1 = 8'd39; b_mant2 = 8'd9; b_mant3 = 8'd89;
a_exp0 = 10'd27; a_exp1 = 10'd99; a_exp2 = 10'd722; a_exp3 = 10'd989;
b_exp0 = 10'd700; b_exp1 = 10'd983; b_exp2 = 10'd464; b_exp3 = 10'd300;
a_sign0 = 4'd9; a_sign1 = 4'd1; a_sign2 = 4'd12; a_sign3 = 4'd5;
b_sign0 = 4'd10; b_sign1 = 4'd3; b_sign2 = 4'd12; b_sign3 = 4'd13;
@(posedge clk_i);
a_mant0 = 8'd218; a_mant1 = 8'd251; a_mant2 = 8'd254; a_mant3 = 8'd95;
b_mant0 = 8'd219; b_mant1 = 8'd234; b_mant2 = 8'd15; b_mant3 = 8'd70;
a_exp0 = 10'd742; a_exp1 = 10'd624; a_exp2 = 10'd827; a_exp3 = 10'd360;
b_exp0 = 10'd868; b_exp1 = 10'd125; b_exp2 = 10'd649; b_exp3 = 10'd550;
a_sign0 = 4'd16; a_sign1 = 4'd10; a_sign2 = 4'd4; a_sign3 = 4'd0;
b_sign0 = 4'd0; b_sign1 = 4'd10; b_sign2 = 4'd10; b_sign3 = 4'd11;
@(posedge clk_i);
a_mant0 = 8'd79; a_mant1 = 8'd227; a_mant2 = 8'd184; a_mant3 = 8'd120;
b_mant0 = 8'd170; b_mant1 = 8'd52; b_mant2 = 8'd72; b_mant3 = 8'd118;
a_exp0 = 10'd712; a_exp1 = 10'd162; a_exp2 = 10'd625; a_exp3 = 10'd271;
b_exp0 = 10'd112; b_exp1 = 10'd1019; b_exp2 = 10'd128; b_exp3 = 10'd312;
a_sign0 = 4'd6; a_sign1 = 4'd6; a_sign2 = 4'd0; a_sign3 = 4'd6;
b_sign0 = 4'd1; b_sign1 = 4'd1; b_sign2 = 4'd11; b_sign3 = 4'd4;
@(posedge clk_i);
a_mant0 = 8'd218; a_mant1 = 8'd255; a_mant2 = 8'd255; a_mant3 = 8'd252;
b_mant0 = 8'd191; b_mant1 = 8'd221; b_mant2 = 8'd100; b_mant3 = 8'd170;
a_exp0 = 10'd978; a_exp1 = 10'd17; a_exp2 = 10'd347; a_exp3 = 10'd115;
b_exp0 = 10'd737; b_exp1 = 10'd243; b_exp2 = 10'd933; b_exp3 = 10'd882;
a_sign0 = 4'd8; a_sign1 = 4'd16; a_sign2 = 4'd15; a_sign3 = 4'd10;
b_sign0 = 4'd16; b_sign1 = 4'd2; b_sign2 = 4'd1; b_sign3 = 4'd1;
@(posedge clk_i);
a_mant0 = 8'd42; a_mant1 = 8'd115; a_mant2 = 8'd178; a_mant3 = 8'd184;
b_mant0 = 8'd98; b_mant1 = 8'd144; b_mant2 = 8'd114; b_mant3 = 8'd205;
a_exp0 = 10'd292; a_exp1 = 10'd20; a_exp2 = 10'd326; a_exp3 = 10'd38;
b_exp0 = 10'd808; b_exp1 = 10'd578; b_exp2 = 10'd759; b_exp3 = 10'd948;
a_sign0 = 4'd1; a_sign1 = 4'd14; a_sign2 = 4'd10; a_sign3 = 4'd12;
b_sign0 = 4'd3; b_sign1 = 4'd0; b_sign2 = 4'd7; b_sign3 = 4'd6;
@(posedge clk_i);
a_mant0 = 8'd130; a_mant1 = 8'd238; a_mant2 = 8'd201; a_mant3 = 8'd63;
b_mant0 = 8'd81; b_mant1 = 8'd183; b_mant2 = 8'd171; b_mant3 = 8'd158;
a_exp0 = 10'd4; a_exp1 = 10'd845; a_exp2 = 10'd818; a_exp3 = 10'd294;
b_exp0 = 10'd756; b_exp1 = 10'd861; b_exp2 = 10'd692; b_exp3 = 10'd688;
a_sign0 = 4'd13; a_sign1 = 4'd3; a_sign2 = 4'd4; a_sign3 = 4'd14;
b_sign0 = 4'd12; b_sign1 = 4'd7; b_sign2 = 4'd13; b_sign3 = 4'd13;
@(posedge clk_i);
shared_exps0 = 8'd101;
shared_exps1 = 8'd135;
rstn = 0;
@(posedge clk_i);
rstn = 1;
a_mant0 = 8'd7; a_mant1 = 8'd245; a_mant2 = 8'd201; a_mant3 = 8'd207;
b_mant0 = 8'd164; b_mant1 = 8'd214; b_mant2 = 8'd182; b_mant3 = 8'd55;
a_exp0 = 10'd1023; a_exp1 = 10'd301; a_exp2 = 10'd804; a_exp3 = 10'd716;
b_exp0 = 10'd639; b_exp1 = 10'd87; b_exp2 = 10'd226; b_exp3 = 10'd750;
a_sign0 = 4'd2; a_sign1 = 4'd11; a_sign2 = 4'd2; a_sign3 = 4'd6;
b_sign0 = 4'd9; b_sign1 = 4'd3; b_sign2 = 4'd4; b_sign3 = 4'd3;
@(posedge clk_i);
a_mant0 = 8'd199; a_mant1 = 8'd187; a_mant2 = 8'd25; a_mant3 = 8'd140;
b_mant0 = 8'd177; b_mant1 = 8'd145; b_mant2 = 8'd83; b_mant3 = 8'd24;
a_exp0 = 10'd709; a_exp1 = 10'd889; a_exp2 = 10'd99; a_exp3 = 10'd292;
b_exp0 = 10'd668; b_exp1 = 10'd221; b_exp2 = 10'd45; b_exp3 = 10'd133;
a_sign0 = 4'd12; a_sign1 = 4'd15; a_sign2 = 4'd3; a_sign3 = 4'd12;
b_sign0 = 4'd4; b_sign1 = 4'd11; b_sign2 = 4'd1; b_sign3 = 4'd1;
@(posedge clk_i);
a_mant0 = 8'd177; a_mant1 = 8'd92; a_mant2 = 8'd101; a_mant3 = 8'd207;
b_mant0 = 8'd131; b_mant1 = 8'd204; b_mant2 = 8'd108; b_mant3 = 8'd91;
a_exp0 = 10'd842; a_exp1 = 10'd190; a_exp2 = 10'd724; a_exp3 = 10'd542;
b_exp0 = 10'd54; b_exp1 = 10'd183; b_exp2 = 10'd579; b_exp3 = 10'd268;
a_sign0 = 4'd5; a_sign1 = 4'd7; a_sign2 = 4'd13; a_sign3 = 4'd13;
b_sign0 = 4'd4; b_sign1 = 4'd2; b_sign2 = 4'd3; b_sign3 = 4'd10;
@(posedge clk_i);
a_mant0 = 8'd123; a_mant1 = 8'd123; a_mant2 = 8'd91; a_mant3 = 8'd62;
b_mant0 = 8'd83; b_mant1 = 8'd32; b_mant2 = 8'd237; b_mant3 = 8'd103;
a_exp0 = 10'd472; a_exp1 = 10'd242; a_exp2 = 10'd282; a_exp3 = 10'd745;
b_exp0 = 10'd164; b_exp1 = 10'd794; b_exp2 = 10'd1015; b_exp3 = 10'd311;
a_sign0 = 4'd10; a_sign1 = 4'd2; a_sign2 = 4'd8; a_sign3 = 4'd15;
b_sign0 = 4'd9; b_sign1 = 4'd1; b_sign2 = 4'd12; b_sign3 = 4'd9;
@(posedge clk_i);
a_mant0 = 8'd65; a_mant1 = 8'd192; a_mant2 = 8'd57; a_mant3 = 8'd226;
b_mant0 = 8'd162; b_mant1 = 8'd27; b_mant2 = 8'd203; b_mant3 = 8'd9;
a_exp0 = 10'd722; a_exp1 = 10'd651; a_exp2 = 10'd357; a_exp3 = 10'd276;
b_exp0 = 10'd678; b_exp1 = 10'd442; b_exp2 = 10'd46; b_exp3 = 10'd670;
a_sign0 = 4'd4; a_sign1 = 4'd11; a_sign2 = 4'd4; a_sign3 = 4'd11;
b_sign0 = 4'd8; b_sign1 = 4'd2; b_sign2 = 4'd9; b_sign3 = 4'd0;
@(posedge clk_i);
a_mant0 = 8'd212; a_mant1 = 8'd92; a_mant2 = 8'd76; a_mant3 = 8'd243;
b_mant0 = 8'd34; b_mant1 = 8'd106; b_mant2 = 8'd218; b_mant3 = 8'd27;
a_exp0 = 10'd554; a_exp1 = 10'd912; a_exp2 = 10'd513; a_exp3 = 10'd208;
b_exp0 = 10'd883; b_exp1 = 10'd568; b_exp2 = 10'd954; b_exp3 = 10'd826;
a_sign0 = 4'd4; a_sign1 = 4'd7; a_sign2 = 4'd14; a_sign3 = 4'd12;
b_sign0 = 4'd7; b_sign1 = 4'd5; b_sign2 = 4'd7; b_sign3 = 4'd16;
@(posedge clk_i);
a_mant0 = 8'd147; a_mant1 = 8'd222; a_mant2 = 8'd163; a_mant3 = 8'd210;
b_mant0 = 8'd102; b_mant1 = 8'd134; b_mant2 = 8'd229; b_mant3 = 8'd146;
a_exp0 = 10'd659; a_exp1 = 10'd607; a_exp2 = 10'd555; a_exp3 = 10'd620;
b_exp0 = 10'd286; b_exp1 = 10'd258; b_exp2 = 10'd645; b_exp3 = 10'd345;
a_sign0 = 4'd4; a_sign1 = 4'd6; a_sign2 = 4'd14; a_sign3 = 4'd11;
b_sign0 = 4'd2; b_sign1 = 4'd0; b_sign2 = 4'd10; b_sign3 = 4'd14;
@(posedge clk_i);
shared_exps0 = 8'd140;
shared_exps1 = 8'd114;
a_mant0 = 8'd216; a_mant1 = 8'd212; a_mant2 = 8'd182; a_mant3 = 8'd45;
b_mant0 = 8'd179; b_mant1 = 8'd252; b_mant2 = 8'd177; b_mant3 = 8'd102;
a_exp0 = 10'd235; a_exp1 = 10'd780; a_exp2 = 10'd743; a_exp3 = 10'd399;
b_exp0 = 10'd963; b_exp1 = 10'd55; b_exp2 = 10'd331; b_exp3 = 10'd841;
a_sign0 = 4'd5; a_sign1 = 4'd5; a_sign2 = 4'd7; a_sign3 = 4'd7;
b_sign0 = 4'd4; b_sign1 = 4'd5; b_sign2 = 4'd16; b_sign3 = 4'd8;
@(posedge clk_i);
a_mant0 = 8'd129; a_mant1 = 8'd23; a_mant2 = 8'd191; a_mant3 = 8'd126;
b_mant0 = 8'd226; b_mant1 = 8'd70; b_mant2 = 8'd14; b_mant3 = 8'd200;
a_exp0 = 10'd16; a_exp1 = 10'd400; a_exp2 = 10'd831; a_exp3 = 10'd134;
b_exp0 = 10'd463; b_exp1 = 10'd130; b_exp2 = 10'd599; b_exp3 = 10'd688;
a_sign0 = 4'd4; a_sign1 = 4'd11; a_sign2 = 4'd5; a_sign3 = 4'd16;
b_sign0 = 4'd15; b_sign1 = 4'd8; b_sign2 = 4'd6; b_sign3 = 4'd7;
@(posedge clk_i);
a_mant0 = 8'd82; a_mant1 = 8'd155; a_mant2 = 8'd143; a_mant3 = 8'd74;
b_mant0 = 8'd78; b_mant1 = 8'd254; b_mant2 = 8'd178; b_mant3 = 8'd33;
a_exp0 = 10'd786; a_exp1 = 10'd597; a_exp2 = 10'd104; a_exp3 = 10'd852;
b_exp0 = 10'd917; b_exp1 = 10'd584; b_exp2 = 10'd637; b_exp3 = 10'd936;
a_sign0 = 4'd3; a_sign1 = 4'd1; a_sign2 = 4'd8; a_sign3 = 4'd3;
b_sign0 = 4'd3; b_sign1 = 4'd6; b_sign2 = 4'd16; b_sign3 = 4'd10;
@(posedge clk_i);
a_mant0 = 8'd215; a_mant1 = 8'd118; a_mant2 = 8'd252; a_mant3 = 8'd114;
b_mant0 = 8'd152; b_mant1 = 8'd204; b_mant2 = 8'd186; b_mant3 = 8'd81;
a_exp0 = 10'd101; a_exp1 = 10'd551; a_exp2 = 10'd79; a_exp3 = 10'd950;
b_exp0 = 10'd776; b_exp1 = 10'd325; b_exp2 = 10'd972; b_exp3 = 10'd944;
a_sign0 = 4'd4; a_sign1 = 4'd7; a_sign2 = 4'd8; a_sign3 = 4'd10;
b_sign0 = 4'd1; b_sign1 = 4'd5; b_sign2 = 4'd0; b_sign3 = 4'd10;
@(posedge clk_i);
a_mant0 = 8'd133; a_mant1 = 8'd145; a_mant2 = 8'd251; a_mant3 = 8'd218;
b_mant0 = 8'd163; b_mant1 = 8'd23; b_mant2 = 8'd41; b_mant3 = 8'd213;
a_exp0 = 10'd1010; a_exp1 = 10'd687; a_exp2 = 10'd555; a_exp3 = 10'd765;
b_exp0 = 10'd746; b_exp1 = 10'd972; b_exp2 = 10'd990; b_exp3 = 10'd254;
a_sign0 = 4'd14; a_sign1 = 4'd8; a_sign2 = 4'd13; a_sign3 = 4'd3;
b_sign0 = 4'd12; b_sign1 = 4'd13; b_sign2 = 4'd8; b_sign3 = 4'd3;
@(posedge clk_i);
a_mant0 = 8'd7; a_mant1 = 8'd15; a_mant2 = 8'd134; a_mant3 = 8'd247;
b_mant0 = 8'd242; b_mant1 = 8'd200; b_mant2 = 8'd206; b_mant3 = 8'd6;
a_exp0 = 10'd816; a_exp1 = 10'd19; a_exp2 = 10'd364; a_exp3 = 10'd845;
b_exp0 = 10'd425; b_exp1 = 10'd662; b_exp2 = 10'd737; b_exp3 = 10'd469;
a_sign0 = 4'd6; a_sign1 = 4'd0; a_sign2 = 4'd3; a_sign3 = 4'd13;
b_sign0 = 4'd15; b_sign1 = 4'd6; b_sign2 = 4'd15; b_sign3 = 4'd5;
@(posedge clk_i);
a_mant0 = 8'd208; a_mant1 = 8'd209; a_mant2 = 8'd109; a_mant3 = 8'd188;
b_mant0 = 8'd93; b_mant1 = 8'd27; b_mant2 = 8'd61; b_mant3 = 8'd96;
a_exp0 = 10'd576; a_exp1 = 10'd759; a_exp2 = 10'd395; a_exp3 = 10'd948;
b_exp0 = 10'd536; b_exp1 = 10'd804; b_exp2 = 10'd410; b_exp3 = 10'd152;
a_sign0 = 4'd12; a_sign1 = 4'd10; a_sign2 = 4'd9; a_sign3 = 4'd2;
b_sign0 = 4'd9; b_sign1 = 4'd1; b_sign2 = 4'd9; b_sign3 = 4'd12;
@(posedge clk_i);
a_mant0 = 8'd129; a_mant1 = 8'd89; a_mant2 = 8'd143; a_mant3 = 8'd150;
b_mant0 = 8'd199; b_mant1 = 8'd251; b_mant2 = 8'd41; b_mant3 = 8'd178;
a_exp0 = 10'd92; a_exp1 = 10'd802; a_exp2 = 10'd504; a_exp3 = 10'd665;
b_exp0 = 10'd252; b_exp1 = 10'd515; b_exp2 = 10'd921; b_exp3 = 10'd304;
a_sign0 = 4'd0; a_sign1 = 4'd7; a_sign2 = 4'd5; a_sign3 = 4'd5;
b_sign0 = 4'd3; b_sign1 = 4'd6; b_sign2 = 4'd15; b_sign3 = 4'd15;
@(posedge clk_i);
shared_exps0 = 8'd128;
shared_exps1 = 8'd117;
a_mant0 = 8'd182; a_mant1 = 8'd223; a_mant2 = 8'd86; a_mant3 = 8'd35;
b_mant0 = 8'd85; b_mant1 = 8'd60; b_mant2 = 8'd228; b_mant3 = 8'd231;
a_exp0 = 10'd844; a_exp1 = 10'd142; a_exp2 = 10'd474; a_exp3 = 10'd862;
b_exp0 = 10'd975; b_exp1 = 10'd422; b_exp2 = 10'd967; b_exp3 = 10'd271;
a_sign0 = 4'd13; a_sign1 = 4'd2; a_sign2 = 4'd15; a_sign3 = 4'd6;
b_sign0 = 4'd14; b_sign1 = 4'd12; b_sign2 = 4'd6; b_sign3 = 4'd10;
@(posedge clk_i);
a_mant0 = 8'd200; a_mant1 = 8'd41; a_mant2 = 8'd16; a_mant3 = 8'd57;
b_mant0 = 8'd183; b_mant1 = 8'd43; b_mant2 = 8'd40; b_mant3 = 8'd119;
a_exp0 = 10'd938; a_exp1 = 10'd698; a_exp2 = 10'd817; a_exp3 = 10'd837;
b_exp0 = 10'd758; b_exp1 = 10'd125; b_exp2 = 10'd931; b_exp3 = 10'd36;
a_sign0 = 4'd11; a_sign1 = 4'd10; a_sign2 = 4'd14; a_sign3 = 4'd3;
b_sign0 = 4'd11; b_sign1 = 4'd1; b_sign2 = 4'd0; b_sign3 = 4'd15;
@(posedge clk_i);
a_mant0 = 8'd22; a_mant1 = 8'd20; a_mant2 = 8'd246; a_mant3 = 8'd101;
b_mant0 = 8'd73; b_mant1 = 8'd137; b_mant2 = 8'd254; b_mant3 = 8'd120;
a_exp0 = 10'd58; a_exp1 = 10'd919; a_exp2 = 10'd739; a_exp3 = 10'd598;
b_exp0 = 10'd298; b_exp1 = 10'd121; b_exp2 = 10'd703; b_exp3 = 10'd405;
a_sign0 = 4'd0; a_sign1 = 4'd5; a_sign2 = 4'd1; a_sign3 = 4'd14;
b_sign0 = 4'd1; b_sign1 = 4'd2; b_sign2 = 4'd3; b_sign3 = 4'd8;
@(posedge clk_i);
a_mant0 = 8'd44; a_mant1 = 8'd12; a_mant2 = 8'd60; a_mant3 = 8'd131;
b_mant0 = 8'd71; b_mant1 = 8'd18; b_mant2 = 8'd206; b_mant3 = 8'd222;
a_exp0 = 10'd689; a_exp1 = 10'd597; a_exp2 = 10'd915; a_exp3 = 10'd494;
b_exp0 = 10'd794; b_exp1 = 10'd130; b_exp2 = 10'd356; b_exp3 = 10'd1000;
a_sign0 = 4'd3; a_sign1 = 4'd4; a_sign2 = 4'd0; a_sign3 = 4'd12;
b_sign0 = 4'd11; b_sign1 = 4'd12; b_sign2 = 4'd12; b_sign3 = 4'd6;
@(posedge clk_i);
a_mant0 = 8'd178; a_mant1 = 8'd45; a_mant2 = 8'd205; a_mant3 = 8'd11;
b_mant0 = 8'd215; b_mant1 = 8'd51; b_mant2 = 8'd133; b_mant3 = 8'd251;
a_exp0 = 10'd556; a_exp1 = 10'd33; a_exp2 = 10'd418; a_exp3 = 10'd577;
b_exp0 = 10'd391; b_exp1 = 10'd198; b_exp2 = 10'd128; b_exp3 = 10'd141;
a_sign0 = 4'd9; a_sign1 = 4'd7; a_sign2 = 4'd15; a_sign3 = 4'd15;
b_sign0 = 4'd11; b_sign1 = 4'd0; b_sign2 = 4'd15; b_sign3 = 4'd6;
@(posedge clk_i);
a_mant0 = 8'd103; a_mant1 = 8'd15; a_mant2 = 8'd188; a_mant3 = 8'd52;
b_mant0 = 8'd222; b_mant1 = 8'd79; b_mant2 = 8'd20; b_mant3 = 8'd213;
a_exp0 = 10'd6; a_exp1 = 10'd505; a_exp2 = 10'd635; a_exp3 = 10'd66;
b_exp0 = 10'd554; b_exp1 = 10'd401; b_exp2 = 10'd661; b_exp3 = 10'd692;
a_sign0 = 4'd16; a_sign1 = 4'd6; a_sign2 = 4'd6; a_sign3 = 4'd13;
b_sign0 = 4'd11; b_sign1 = 4'd0; b_sign2 = 4'd4; b_sign3 = 4'd15;
@(posedge clk_i);
a_mant0 = 8'd203; a_mant1 = 8'd72; a_mant2 = 8'd159; a_mant3 = 8'd237;
b_mant0 = 8'd57; b_mant1 = 8'd60; b_mant2 = 8'd216; b_mant3 = 8'd14;
a_exp0 = 10'd219; a_exp1 = 10'd335; a_exp2 = 10'd715; a_exp3 = 10'd750;
b_exp0 = 10'd325; b_exp1 = 10'd512; b_exp2 = 10'd39; b_exp3 = 10'd218;
a_sign0 = 4'd6; a_sign1 = 4'd12; a_sign2 = 4'd11; a_sign3 = 4'd7;
b_sign0 = 4'd7; b_sign1 = 4'd11; b_sign2 = 4'd12; b_sign3 = 4'd8;
@(posedge clk_i);
a_mant0 = 8'd216; a_mant1 = 8'd53; a_mant2 = 8'd13; a_mant3 = 8'd173;
b_mant0 = 8'd11; b_mant1 = 8'd167; b_mant2 = 8'd26; b_mant3 = 8'd58;
a_exp0 = 10'd172; a_exp1 = 10'd855; a_exp2 = 10'd428; a_exp3 = 10'd761;
b_exp0 = 10'd682; b_exp1 = 10'd691; b_exp2 = 10'd887; b_exp3 = 10'd554;
a_sign0 = 4'd6; a_sign1 = 4'd6; a_sign2 = 4'd2; a_sign3 = 4'd7;
b_sign0 = 4'd12; b_sign1 = 4'd6; b_sign2 = 4'd14; b_sign3 = 4'd9;
@(posedge clk_i);
shared_exps0 = 8'd116;
shared_exps1 = 8'd116;
a_mant0 = 8'd18; a_mant1 = 8'd1; a_mant2 = 8'd48; a_mant3 = 8'd104;
b_mant0 = 8'd14; b_mant1 = 8'd192; b_mant2 = 8'd73; b_mant3 = 8'd0;
a_exp0 = 10'd377; a_exp1 = 10'd953; a_exp2 = 10'd932; a_exp3 = 10'd712;
b_exp0 = 10'd939; b_exp1 = 10'd141; b_exp2 = 10'd480; b_exp3 = 10'd175;
a_sign0 = 4'd0; a_sign1 = 4'd7; a_sign2 = 4'd2; a_sign3 = 4'd10;
b_sign0 = 4'd15; b_sign1 = 4'd5; b_sign2 = 4'd3; b_sign3 = 4'd5;
@(posedge clk_i);
a_mant0 = 8'd219; a_mant1 = 8'd174; a_mant2 = 8'd60; a_mant3 = 8'd9;
b_mant0 = 8'd171; b_mant1 = 8'd39; b_mant2 = 8'd109; b_mant3 = 8'd132;
a_exp0 = 10'd854; a_exp1 = 10'd75; a_exp2 = 10'd310; a_exp3 = 10'd548;
b_exp0 = 10'd906; b_exp1 = 10'd645; b_exp2 = 10'd621; b_exp3 = 10'd363;
a_sign0 = 4'd11; a_sign1 = 4'd3; a_sign2 = 4'd1; a_sign3 = 4'd0;
b_sign0 = 4'd4; b_sign1 = 4'd14; b_sign2 = 4'd9; b_sign3 = 4'd3;
@(posedge clk_i);
a_mant0 = 8'd173; a_mant1 = 8'd1; a_mant2 = 8'd134; a_mant3 = 8'd184;
b_mant0 = 8'd156; b_mant1 = 8'd186; b_mant2 = 8'd115; b_mant3 = 8'd228;
a_exp0 = 10'd107; a_exp1 = 10'd444; a_exp2 = 10'd1020; a_exp3 = 10'd786;
b_exp0 = 10'd429; b_exp1 = 10'd117; b_exp2 = 10'd482; b_exp3 = 10'd798;
a_sign0 = 4'd7; a_sign1 = 4'd12; a_sign2 = 4'd3; a_sign3 = 4'd9;
b_sign0 = 4'd7; b_sign1 = 4'd6; b_sign2 = 4'd5; b_sign3 = 4'd12;
@(posedge clk_i);
a_mant0 = 8'd228; a_mant1 = 8'd204; a_mant2 = 8'd128; a_mant3 = 8'd155;
b_mant0 = 8'd167; b_mant1 = 8'd13; b_mant2 = 8'd0; b_mant3 = 8'd151;
a_exp0 = 10'd613; a_exp1 = 10'd913; a_exp2 = 10'd96; a_exp3 = 10'd293;
b_exp0 = 10'd146; b_exp1 = 10'd687; b_exp2 = 10'd661; b_exp3 = 10'd830;
a_sign0 = 4'd10; a_sign1 = 4'd10; a_sign2 = 4'd14; a_sign3 = 4'd7;
b_sign0 = 4'd9; b_sign1 = 4'd14; b_sign2 = 4'd4; b_sign3 = 4'd7;
@(posedge clk_i);
a_mant0 = 8'd208; a_mant1 = 8'd158; a_mant2 = 8'd8; a_mant3 = 8'd3;
b_mant0 = 8'd239; b_mant1 = 8'd12; b_mant2 = 8'd89; b_mant3 = 8'd23;
a_exp0 = 10'd572; a_exp1 = 10'd709; a_exp2 = 10'd412; a_exp3 = 10'd458;
b_exp0 = 10'd961; b_exp1 = 10'd274; b_exp2 = 10'd884; b_exp3 = 10'd501;
a_sign0 = 4'd8; a_sign1 = 4'd8; a_sign2 = 4'd14; a_sign3 = 4'd11;
b_sign0 = 4'd5; b_sign1 = 4'd2; b_sign2 = 4'd4; b_sign3 = 4'd7;
@(posedge clk_i);
a_mant0 = 8'd125; a_mant1 = 8'd143; a_mant2 = 8'd104; a_mant3 = 8'd33;
b_mant0 = 8'd53; b_mant1 = 8'd80; b_mant2 = 8'd5; b_mant3 = 8'd133;
a_exp0 = 10'd784; a_exp1 = 10'd169; a_exp2 = 10'd4; a_exp3 = 10'd280;
b_exp0 = 10'd869; b_exp1 = 10'd534; b_exp2 = 10'd919; b_exp3 = 10'd140;
a_sign0 = 4'd12; a_sign1 = 4'd5; a_sign2 = 4'd9; a_sign3 = 4'd9;
b_sign0 = 4'd6; b_sign1 = 4'd6; b_sign2 = 4'd2; b_sign3 = 4'd8;
@(posedge clk_i);
a_mant0 = 8'd177; a_mant1 = 8'd7; a_mant2 = 8'd137; a_mant3 = 8'd126;
b_mant0 = 8'd133; b_mant1 = 8'd79; b_mant2 = 8'd124; b_mant3 = 8'd148;
a_exp0 = 10'd568; a_exp1 = 10'd804; a_exp2 = 10'd719; a_exp3 = 10'd161;
b_exp0 = 10'd274; b_exp1 = 10'd1013; b_exp2 = 10'd174; b_exp3 = 10'd108;
a_sign0 = 4'd0; a_sign1 = 4'd5; a_sign2 = 4'd1; a_sign3 = 4'd4;
b_sign0 = 4'd12; b_sign1 = 4'd0; b_sign2 = 4'd12; b_sign3 = 4'd9;
@(posedge clk_i);
a_mant0 = 8'd135; a_mant1 = 8'd125; a_mant2 = 8'd51; a_mant3 = 8'd36;
b_mant0 = 8'd41; b_mant1 = 8'd44; b_mant2 = 8'd59; b_mant3 = 8'd124;
a_exp0 = 10'd875; a_exp1 = 10'd197; a_exp2 = 10'd831; a_exp3 = 10'd799;
b_exp0 = 10'd428; b_exp1 = 10'd289; b_exp2 = 10'd160; b_exp3 = 10'd634;
a_sign0 = 4'd5; a_sign1 = 4'd8; a_sign2 = 4'd9; a_sign3 = 4'd2;
b_sign0 = 4'd15; b_sign1 = 4'd15; b_sign2 = 4'd9; b_sign3 = 4'd14;
@(posedge clk_i);
shared_exps0 = 8'd104;
shared_exps1 = 8'd108;
rstn = 0;
@(posedge clk_i);
rstn = 1;
a_mant0 = 8'd151; a_mant1 = 8'd132; a_mant2 = 8'd33; a_mant3 = 8'd36;
b_mant0 = 8'd137; b_mant1 = 8'd108; b_mant2 = 8'd29; b_mant3 = 8'd28;
a_exp0 = 10'd596; a_exp1 = 10'd985; a_exp2 = 10'd127; a_exp3 = 10'd146;
b_exp0 = 10'd196; b_exp1 = 10'd53; b_exp2 = 10'd614; b_exp3 = 10'd99;
a_sign0 = 4'd5; a_sign1 = 4'd1; a_sign2 = 4'd4; a_sign3 = 4'd2;
b_sign0 = 4'd13; b_sign1 = 4'd8; b_sign2 = 4'd8; b_sign3 = 4'd14;
@(posedge clk_i);
a_mant0 = 8'd94; a_mant1 = 8'd6; a_mant2 = 8'd206; a_mant3 = 8'd236;
b_mant0 = 8'd154; b_mant1 = 8'd97; b_mant2 = 8'd153; b_mant3 = 8'd65;
a_exp0 = 10'd682; a_exp1 = 10'd428; a_exp2 = 10'd144; a_exp3 = 10'd847;
b_exp0 = 10'd854; b_exp1 = 10'd249; b_exp2 = 10'd484; b_exp3 = 10'd88;
a_sign0 = 4'd6; a_sign1 = 4'd3; a_sign2 = 4'd2; a_sign3 = 4'd9;
b_sign0 = 4'd12; b_sign1 = 4'd0; b_sign2 = 4'd10; b_sign3 = 4'd4;
@(posedge clk_i);
a_mant0 = 8'd116; a_mant1 = 8'd223; a_mant2 = 8'd186; a_mant3 = 8'd21;
b_mant0 = 8'd107; b_mant1 = 8'd105; b_mant2 = 8'd105; b_mant3 = 8'd79;
a_exp0 = 10'd830; a_exp1 = 10'd469; a_exp2 = 10'd587; a_exp3 = 10'd666;
b_exp0 = 10'd866; b_exp1 = 10'd297; b_exp2 = 10'd580; b_exp3 = 10'd862;
a_sign0 = 4'd10; a_sign1 = 4'd5; a_sign2 = 4'd7; a_sign3 = 4'd4;
b_sign0 = 4'd6; b_sign1 = 4'd1; b_sign2 = 4'd3; b_sign3 = 4'd14;
@(posedge clk_i);
a_mant0 = 8'd158; a_mant1 = 8'd189; a_mant2 = 8'd17; a_mant3 = 8'd37;
b_mant0 = 8'd209; b_mant1 = 8'd113; b_mant2 = 8'd213; b_mant3 = 8'd30;
a_exp0 = 10'd355; a_exp1 = 10'd460; a_exp2 = 10'd557; a_exp3 = 10'd268;
b_exp0 = 10'd671; b_exp1 = 10'd326; b_exp2 = 10'd903; b_exp3 = 10'd237;
a_sign0 = 4'd1; a_sign1 = 4'd6; a_sign2 = 4'd0; a_sign3 = 4'd2;
b_sign0 = 4'd0; b_sign1 = 4'd4; b_sign2 = 4'd0; b_sign3 = 4'd10;
@(posedge clk_i);
a_mant0 = 8'd169; a_mant1 = 8'd8; a_mant2 = 8'd54; a_mant3 = 8'd228;
b_mant0 = 8'd34; b_mant1 = 8'd233; b_mant2 = 8'd91; b_mant3 = 8'd193;
a_exp0 = 10'd435; a_exp1 = 10'd40; a_exp2 = 10'd667; a_exp3 = 10'd694;
b_exp0 = 10'd129; b_exp1 = 10'd287; b_exp2 = 10'd234; b_exp3 = 10'd190;
a_sign0 = 4'd14; a_sign1 = 4'd0; a_sign2 = 4'd11; a_sign3 = 4'd13;
b_sign0 = 4'd12; b_sign1 = 4'd9; b_sign2 = 4'd4; b_sign3 = 4'd3;
@(posedge clk_i);
a_mant0 = 8'd234; a_mant1 = 8'd185; a_mant2 = 8'd59; a_mant3 = 8'd104;
b_mant0 = 8'd23; b_mant1 = 8'd210; b_mant2 = 8'd184; b_mant3 = 8'd95;
a_exp0 = 10'd373; a_exp1 = 10'd172; a_exp2 = 10'd697; a_exp3 = 10'd463;
b_exp0 = 10'd62; b_exp1 = 10'd424; b_exp2 = 10'd475; b_exp3 = 10'd529;
a_sign0 = 4'd7; a_sign1 = 4'd3; a_sign2 = 4'd7; a_sign3 = 4'd15;
b_sign0 = 4'd14; b_sign1 = 4'd6; b_sign2 = 4'd4; b_sign3 = 4'd3;
@(posedge clk_i);
a_mant0 = 8'd139; a_mant1 = 8'd206; a_mant2 = 8'd75; a_mant3 = 8'd205;
b_mant0 = 8'd95; b_mant1 = 8'd242; b_mant2 = 8'd46; b_mant3 = 8'd28;
a_exp0 = 10'd797; a_exp1 = 10'd557; a_exp2 = 10'd749; a_exp3 = 10'd377;
b_exp0 = 10'd581; b_exp1 = 10'd1000; b_exp2 = 10'd297; b_exp3 = 10'd272;
a_sign0 = 4'd8; a_sign1 = 4'd16; a_sign2 = 4'd12; a_sign3 = 4'd16;
b_sign0 = 4'd15; b_sign1 = 4'd5; b_sign2 = 4'd11; b_sign3 = 4'd5;
@(posedge clk_i);
shared_exps0 = 8'd118;
shared_exps1 = 8'd150;
a_mant0 = 8'd175; a_mant1 = 8'd243; a_mant2 = 8'd65; a_mant3 = 8'd241;
b_mant0 = 8'd172; b_mant1 = 8'd92; b_mant2 = 8'd244; b_mant3 = 8'd251;
a_exp0 = 10'd679; a_exp1 = 10'd167; a_exp2 = 10'd184; a_exp3 = 10'd907;
b_exp0 = 10'd602; b_exp1 = 10'd125; b_exp2 = 10'd349; b_exp3 = 10'd427;
a_sign0 = 4'd12; a_sign1 = 4'd4; a_sign2 = 4'd0; a_sign3 = 4'd5;
b_sign0 = 4'd6; b_sign1 = 4'd7; b_sign2 = 4'd0; b_sign3 = 4'd7;
@(posedge clk_i);
a_mant0 = 8'd136; a_mant1 = 8'd51; a_mant2 = 8'd95; a_mant3 = 8'd55;
b_mant0 = 8'd229; b_mant1 = 8'd247; b_mant2 = 8'd233; b_mant3 = 8'd21;
a_exp0 = 10'd800; a_exp1 = 10'd276; a_exp2 = 10'd422; a_exp3 = 10'd255;
b_exp0 = 10'd827; b_exp1 = 10'd198; b_exp2 = 10'd870; b_exp3 = 10'd893;
a_sign0 = 4'd1; a_sign1 = 4'd16; a_sign2 = 4'd4; a_sign3 = 4'd15;
b_sign0 = 4'd3; b_sign1 = 4'd0; b_sign2 = 4'd2; b_sign3 = 4'd10;
@(posedge clk_i);
a_mant0 = 8'd139; a_mant1 = 8'd235; a_mant2 = 8'd9; a_mant3 = 8'd128;
b_mant0 = 8'd29; b_mant1 = 8'd110; b_mant2 = 8'd73; b_mant3 = 8'd68;
a_exp0 = 10'd658; a_exp1 = 10'd837; a_exp2 = 10'd249; a_exp3 = 10'd548;
b_exp0 = 10'd750; b_exp1 = 10'd151; b_exp2 = 10'd188; b_exp3 = 10'd678;
a_sign0 = 4'd0; a_sign1 = 4'd7; a_sign2 = 4'd4; a_sign3 = 4'd8;
b_sign0 = 4'd11; b_sign1 = 4'd8; b_sign2 = 4'd5; b_sign3 = 4'd9;
@(posedge clk_i);
a_mant0 = 8'd190; a_mant1 = 8'd61; a_mant2 = 8'd144; a_mant3 = 8'd124;
b_mant0 = 8'd212; b_mant1 = 8'd21; b_mant2 = 8'd54; b_mant3 = 8'd23;
a_exp0 = 10'd817; a_exp1 = 10'd92; a_exp2 = 10'd398; a_exp3 = 10'd929;
b_exp0 = 10'd408; b_exp1 = 10'd880; b_exp2 = 10'd706; b_exp3 = 10'd297;
a_sign0 = 4'd2; a_sign1 = 4'd4; a_sign2 = 4'd1; a_sign3 = 4'd14;
b_sign0 = 4'd15; b_sign1 = 4'd10; b_sign2 = 4'd3; b_sign3 = 4'd13;
@(posedge clk_i);
a_mant0 = 8'd58; a_mant1 = 8'd146; a_mant2 = 8'd239; a_mant3 = 8'd148;
b_mant0 = 8'd27; b_mant1 = 8'd203; b_mant2 = 8'd141; b_mant3 = 8'd129;
a_exp0 = 10'd554; a_exp1 = 10'd419; a_exp2 = 10'd224; a_exp3 = 10'd304;
b_exp0 = 10'd782; b_exp1 = 10'd263; b_exp2 = 10'd802; b_exp3 = 10'd560;
a_sign0 = 4'd13; a_sign1 = 4'd10; a_sign2 = 4'd8; a_sign3 = 4'd11;
b_sign0 = 4'd13; b_sign1 = 4'd1; b_sign2 = 4'd3; b_sign3 = 4'd15;
@(posedge clk_i);
a_mant0 = 8'd144; a_mant1 = 8'd33; a_mant2 = 8'd18; a_mant3 = 8'd50;
b_mant0 = 8'd200; b_mant1 = 8'd39; b_mant2 = 8'd151; b_mant3 = 8'd173;
a_exp0 = 10'd785; a_exp1 = 10'd681; a_exp2 = 10'd420; a_exp3 = 10'd222;
b_exp0 = 10'd983; b_exp1 = 10'd1002; b_exp2 = 10'd856; b_exp3 = 10'd141;
a_sign0 = 4'd2; a_sign1 = 4'd7; a_sign2 = 4'd11; a_sign3 = 4'd16;
b_sign0 = 4'd13; b_sign1 = 4'd0; b_sign2 = 4'd1; b_sign3 = 4'd12;
@(posedge clk_i);
a_mant0 = 8'd137; a_mant1 = 8'd108; a_mant2 = 8'd50; a_mant3 = 8'd113;
b_mant0 = 8'd185; b_mant1 = 8'd148; b_mant2 = 8'd80; b_mant3 = 8'd24;
a_exp0 = 10'd478; a_exp1 = 10'd400; a_exp2 = 10'd52; a_exp3 = 10'd747;
b_exp0 = 10'd739; b_exp1 = 10'd504; b_exp2 = 10'd682; b_exp3 = 10'd901;
a_sign0 = 4'd11; a_sign1 = 4'd2; a_sign2 = 4'd11; a_sign3 = 4'd12;
b_sign0 = 4'd13; b_sign1 = 4'd13; b_sign2 = 4'd3; b_sign3 = 4'd9;
@(posedge clk_i);
a_mant0 = 8'd33; a_mant1 = 8'd236; a_mant2 = 8'd130; a_mant3 = 8'd120;
b_mant0 = 8'd172; b_mant1 = 8'd7; b_mant2 = 8'd146; b_mant3 = 8'd134;
a_exp0 = 10'd372; a_exp1 = 10'd104; a_exp2 = 10'd77; a_exp3 = 10'd579;
b_exp0 = 10'd990; b_exp1 = 10'd937; b_exp2 = 10'd992; b_exp3 = 10'd753;
a_sign0 = 4'd3; a_sign1 = 4'd0; a_sign2 = 4'd9; a_sign3 = 4'd11;
b_sign0 = 4'd6; b_sign1 = 4'd3; b_sign2 = 4'd11; b_sign3 = 4'd12;
@(posedge clk_i);
shared_exps0 = 8'd111;
shared_exps1 = 8'd112;
a_mant0 = 8'd152; a_mant1 = 8'd34; a_mant2 = 8'd18; a_mant3 = 8'd166;
b_mant0 = 8'd224; b_mant1 = 8'd123; b_mant2 = 8'd204; b_mant3 = 8'd159;
a_exp0 = 10'd606; a_exp1 = 10'd32; a_exp2 = 10'd527; a_exp3 = 10'd17;
b_exp0 = 10'd717; b_exp1 = 10'd681; b_exp2 = 10'd345; b_exp3 = 10'd5;
a_sign0 = 4'd8; a_sign1 = 4'd4; a_sign2 = 4'd2; a_sign3 = 4'd13;
b_sign0 = 4'd10; b_sign1 = 4'd6; b_sign2 = 4'd11; b_sign3 = 4'd11;
@(posedge clk_i);
a_mant0 = 8'd0; a_mant1 = 8'd246; a_mant2 = 8'd247; a_mant3 = 8'd200;
b_mant0 = 8'd241; b_mant1 = 8'd33; b_mant2 = 8'd42; b_mant3 = 8'd55;
a_exp0 = 10'd86; a_exp1 = 10'd564; a_exp2 = 10'd996; a_exp3 = 10'd455;
b_exp0 = 10'd68; b_exp1 = 10'd38; b_exp2 = 10'd360; b_exp3 = 10'd772;
a_sign0 = 4'd13; a_sign1 = 4'd2; a_sign2 = 4'd9; a_sign3 = 4'd16;
b_sign0 = 4'd3; b_sign1 = 4'd1; b_sign2 = 4'd6; b_sign3 = 4'd16;
@(posedge clk_i);
a_mant0 = 8'd191; a_mant1 = 8'd15; a_mant2 = 8'd242; a_mant3 = 8'd130;
b_mant0 = 8'd2; b_mant1 = 8'd148; b_mant2 = 8'd10; b_mant3 = 8'd213;
a_exp0 = 10'd906; a_exp1 = 10'd42; a_exp2 = 10'd456; a_exp3 = 10'd562;
b_exp0 = 10'd579; b_exp1 = 10'd535; b_exp2 = 10'd691; b_exp3 = 10'd215;
a_sign0 = 4'd10; a_sign1 = 4'd6; a_sign2 = 4'd13; a_sign3 = 4'd10;
b_sign0 = 4'd15; b_sign1 = 4'd5; b_sign2 = 4'd4; b_sign3 = 4'd5;
@(posedge clk_i);
a_mant0 = 8'd158; a_mant1 = 8'd239; a_mant2 = 8'd47; a_mant3 = 8'd232;
b_mant0 = 8'd205; b_mant1 = 8'd44; b_mant2 = 8'd157; b_mant3 = 8'd177;
a_exp0 = 10'd465; a_exp1 = 10'd303; a_exp2 = 10'd11; a_exp3 = 10'd352;
b_exp0 = 10'd647; b_exp1 = 10'd1019; b_exp2 = 10'd789; b_exp3 = 10'd150;
a_sign0 = 4'd16; a_sign1 = 4'd15; a_sign2 = 4'd11; a_sign3 = 4'd2;
b_sign0 = 4'd13; b_sign1 = 4'd10; b_sign2 = 4'd6; b_sign3 = 4'd7;
@(posedge clk_i);
a_mant0 = 8'd135; a_mant1 = 8'd212; a_mant2 = 8'd1; a_mant3 = 8'd26;
b_mant0 = 8'd88; b_mant1 = 8'd97; b_mant2 = 8'd94; b_mant3 = 8'd10;
a_exp0 = 10'd712; a_exp1 = 10'd864; a_exp2 = 10'd447; a_exp3 = 10'd637;
b_exp0 = 10'd450; b_exp1 = 10'd315; b_exp2 = 10'd394; b_exp3 = 10'd862;
a_sign0 = 4'd4; a_sign1 = 4'd7; a_sign2 = 4'd16; a_sign3 = 4'd5;
b_sign0 = 4'd2; b_sign1 = 4'd6; b_sign2 = 4'd9; b_sign3 = 4'd15;
@(posedge clk_i);
a_mant0 = 8'd140; a_mant1 = 8'd87; a_mant2 = 8'd180; a_mant3 = 8'd250;
b_mant0 = 8'd94; b_mant1 = 8'd41; b_mant2 = 8'd237; b_mant3 = 8'd103;
a_exp0 = 10'd81; a_exp1 = 10'd397; a_exp2 = 10'd365; a_exp3 = 10'd492;
b_exp0 = 10'd829; b_exp1 = 10'd888; b_exp2 = 10'd614; b_exp3 = 10'd658;
a_sign0 = 4'd7; a_sign1 = 4'd2; a_sign2 = 4'd9; a_sign3 = 4'd2;
b_sign0 = 4'd3; b_sign1 = 4'd7; b_sign2 = 4'd6; b_sign3 = 4'd4;
@(posedge clk_i);
a_mant0 = 8'd128; a_mant1 = 8'd137; a_mant2 = 8'd235; a_mant3 = 8'd122;
b_mant0 = 8'd238; b_mant1 = 8'd167; b_mant2 = 8'd39; b_mant3 = 8'd232;
a_exp0 = 10'd43; a_exp1 = 10'd725; a_exp2 = 10'd215; a_exp3 = 10'd829;
b_exp0 = 10'd254; b_exp1 = 10'd49; b_exp2 = 10'd326; b_exp3 = 10'd791;
a_sign0 = 4'd8; a_sign1 = 4'd5; a_sign2 = 4'd3; a_sign3 = 4'd15;
b_sign0 = 4'd2; b_sign1 = 4'd15; b_sign2 = 4'd0; b_sign3 = 4'd9;
@(posedge clk_i);
a_mant0 = 8'd129; a_mant1 = 8'd104; a_mant2 = 8'd69; a_mant3 = 8'd91;
b_mant0 = 8'd107; b_mant1 = 8'd0; b_mant2 = 8'd164; b_mant3 = 8'd72;
a_exp0 = 10'd470; a_exp1 = 10'd500; a_exp2 = 10'd53; a_exp3 = 10'd222;
b_exp0 = 10'd940; b_exp1 = 10'd286; b_exp2 = 10'd490; b_exp3 = 10'd178;
a_sign0 = 4'd9; a_sign1 = 4'd12; a_sign2 = 4'd9; a_sign3 = 4'd6;
b_sign0 = 4'd13; b_sign1 = 4'd12; b_sign2 = 4'd3; b_sign3 = 4'd14;
@(posedge clk_i);
shared_exps0 = 8'd149;
shared_exps1 = 8'd133;
a_mant0 = 8'd94; a_mant1 = 8'd90; a_mant2 = 8'd21; a_mant3 = 8'd163;
b_mant0 = 8'd83; b_mant1 = 8'd232; b_mant2 = 8'd116; b_mant3 = 8'd132;
a_exp0 = 10'd200; a_exp1 = 10'd583; a_exp2 = 10'd26; a_exp3 = 10'd194;
b_exp0 = 10'd335; b_exp1 = 10'd573; b_exp2 = 10'd455; b_exp3 = 10'd216;
a_sign0 = 4'd14; a_sign1 = 4'd4; a_sign2 = 4'd4; a_sign3 = 4'd12;
b_sign0 = 4'd0; b_sign1 = 4'd15; b_sign2 = 4'd8; b_sign3 = 4'd11;
@(posedge clk_i);
a_mant0 = 8'd109; a_mant1 = 8'd239; a_mant2 = 8'd140; a_mant3 = 8'd69;
b_mant0 = 8'd19; b_mant1 = 8'd46; b_mant2 = 8'd52; b_mant3 = 8'd238;
a_exp0 = 10'd226; a_exp1 = 10'd566; a_exp2 = 10'd529; a_exp3 = 10'd280;
b_exp0 = 10'd816; b_exp1 = 10'd471; b_exp2 = 10'd265; b_exp3 = 10'd192;
a_sign0 = 4'd2; a_sign1 = 4'd0; a_sign2 = 4'd16; a_sign3 = 4'd1;
b_sign0 = 4'd5; b_sign1 = 4'd5; b_sign2 = 4'd7; b_sign3 = 4'd1;
@(posedge clk_i);
a_mant0 = 8'd24; a_mant1 = 8'd219; a_mant2 = 8'd167; a_mant3 = 8'd106;
b_mant0 = 8'd216; b_mant1 = 8'd156; b_mant2 = 8'd8; b_mant3 = 8'd95;
a_exp0 = 10'd689; a_exp1 = 10'd441; a_exp2 = 10'd910; a_exp3 = 10'd682;
b_exp0 = 10'd303; b_exp1 = 10'd967; b_exp2 = 10'd208; b_exp3 = 10'd483;
a_sign0 = 4'd14; a_sign1 = 4'd0; a_sign2 = 4'd13; a_sign3 = 4'd6;
b_sign0 = 4'd5; b_sign1 = 4'd3; b_sign2 = 4'd15; b_sign3 = 4'd11;
@(posedge clk_i);
a_mant0 = 8'd238; a_mant1 = 8'd50; a_mant2 = 8'd100; a_mant3 = 8'd254;
b_mant0 = 8'd242; b_mant1 = 8'd68; b_mant2 = 8'd40; b_mant3 = 8'd56;
a_exp0 = 10'd246; a_exp1 = 10'd768; a_exp2 = 10'd87; a_exp3 = 10'd114;
b_exp0 = 10'd878; b_exp1 = 10'd308; b_exp2 = 10'd310; b_exp3 = 10'd521;
a_sign0 = 4'd11; a_sign1 = 4'd11; a_sign2 = 4'd9; a_sign3 = 4'd7;
b_sign0 = 4'd7; b_sign1 = 4'd5; b_sign2 = 4'd8; b_sign3 = 4'd9;
@(posedge clk_i);
a_mant0 = 8'd200; a_mant1 = 8'd243; a_mant2 = 8'd212; a_mant3 = 8'd69;
b_mant0 = 8'd22; b_mant1 = 8'd206; b_mant2 = 8'd17; b_mant3 = 8'd170;
a_exp0 = 10'd39; a_exp1 = 10'd22; a_exp2 = 10'd349; a_exp3 = 10'd950;
b_exp0 = 10'd489; b_exp1 = 10'd1001; b_exp2 = 10'd184; b_exp3 = 10'd1001;
a_sign0 = 4'd14; a_sign1 = 4'd14; a_sign2 = 4'd7; a_sign3 = 4'd6;
b_sign0 = 4'd7; b_sign1 = 4'd14; b_sign2 = 4'd8; b_sign3 = 4'd0;
@(posedge clk_i);
a_mant0 = 8'd134; a_mant1 = 8'd9; a_mant2 = 8'd160; a_mant3 = 8'd161;
b_mant0 = 8'd164; b_mant1 = 8'd141; b_mant2 = 8'd132; b_mant3 = 8'd214;
a_exp0 = 10'd623; a_exp1 = 10'd243; a_exp2 = 10'd754; a_exp3 = 10'd457;
b_exp0 = 10'd233; b_exp1 = 10'd510; b_exp2 = 10'd471; b_exp3 = 10'd279;
a_sign0 = 4'd4; a_sign1 = 4'd4; a_sign2 = 4'd16; a_sign3 = 4'd0;
b_sign0 = 4'd16; b_sign1 = 4'd6; b_sign2 = 4'd11; b_sign3 = 4'd9;
@(posedge clk_i);
a_mant0 = 8'd171; a_mant1 = 8'd213; a_mant2 = 8'd111; a_mant3 = 8'd119;
b_mant0 = 8'd88; b_mant1 = 8'd1; b_mant2 = 8'd54; b_mant3 = 8'd247;
a_exp0 = 10'd1004; a_exp1 = 10'd118; a_exp2 = 10'd59; a_exp3 = 10'd684;
b_exp0 = 10'd914; b_exp1 = 10'd72; b_exp2 = 10'd146; b_exp3 = 10'd929;
a_sign0 = 4'd5; a_sign1 = 4'd1; a_sign2 = 4'd12; a_sign3 = 4'd15;
b_sign0 = 4'd14; b_sign1 = 4'd4; b_sign2 = 4'd10; b_sign3 = 4'd15;
@(posedge clk_i);
a_mant0 = 8'd184; a_mant1 = 8'd3; a_mant2 = 8'd26; a_mant3 = 8'd161;
b_mant0 = 8'd110; b_mant1 = 8'd5; b_mant2 = 8'd52; b_mant3 = 8'd51;
a_exp0 = 10'd231; a_exp1 = 10'd885; a_exp2 = 10'd406; a_exp3 = 10'd837;
b_exp0 = 10'd993; b_exp1 = 10'd594; b_exp2 = 10'd177; b_exp3 = 10'd659;
a_sign0 = 4'd6; a_sign1 = 4'd5; a_sign2 = 4'd1; a_sign3 = 4'd12;
b_sign0 = 4'd4; b_sign1 = 4'd4; b_sign2 = 4'd16; b_sign3 = 4'd9;
@(posedge clk_i);
shared_exps0 = 8'd134;
shared_exps1 = 8'd134;
rstn = 0;
@(posedge clk_i);
rstn = 1;
a_mant0 = 8'd61; a_mant1 = 8'd11; a_mant2 = 8'd79; a_mant3 = 8'd173;
b_mant0 = 8'd34; b_mant1 = 8'd168; b_mant2 = 8'd67; b_mant3 = 8'd171;
a_exp0 = 10'd296; a_exp1 = 10'd714; a_exp2 = 10'd464; a_exp3 = 10'd515;
b_exp0 = 10'd562; b_exp1 = 10'd329; b_exp2 = 10'd50; b_exp3 = 10'd477;
a_sign0 = 4'd6; a_sign1 = 4'd11; a_sign2 = 4'd15; a_sign3 = 4'd3;
b_sign0 = 4'd8; b_sign1 = 4'd15; b_sign2 = 4'd2; b_sign3 = 4'd12;
@(posedge clk_i);
a_mant0 = 8'd191; a_mant1 = 8'd39; a_mant2 = 8'd65; a_mant3 = 8'd22;
b_mant0 = 8'd155; b_mant1 = 8'd173; b_mant2 = 8'd36; b_mant3 = 8'd147;
a_exp0 = 10'd574; a_exp1 = 10'd360; a_exp2 = 10'd57; a_exp3 = 10'd747;
b_exp0 = 10'd111; b_exp1 = 10'd557; b_exp2 = 10'd742; b_exp3 = 10'd162;
a_sign0 = 4'd6; a_sign1 = 4'd7; a_sign2 = 4'd15; a_sign3 = 4'd0;
b_sign0 = 4'd1; b_sign1 = 4'd10; b_sign2 = 4'd12; b_sign3 = 4'd11;
@(posedge clk_i);
a_mant0 = 8'd70; a_mant1 = 8'd5; a_mant2 = 8'd25; a_mant3 = 8'd218;
b_mant0 = 8'd180; b_mant1 = 8'd31; b_mant2 = 8'd97; b_mant3 = 8'd101;
a_exp0 = 10'd808; a_exp1 = 10'd579; a_exp2 = 10'd970; a_exp3 = 10'd46;
b_exp0 = 10'd336; b_exp1 = 10'd920; b_exp2 = 10'd1018; b_exp3 = 10'd428;
a_sign0 = 4'd11; a_sign1 = 4'd14; a_sign2 = 4'd6; a_sign3 = 4'd5;
b_sign0 = 4'd10; b_sign1 = 4'd15; b_sign2 = 4'd12; b_sign3 = 4'd3;
@(posedge clk_i);
a_mant0 = 8'd249; a_mant1 = 8'd20; a_mant2 = 8'd74; a_mant3 = 8'd157;
b_mant0 = 8'd255; b_mant1 = 8'd149; b_mant2 = 8'd69; b_mant3 = 8'd67;
a_exp0 = 10'd818; a_exp1 = 10'd105; a_exp2 = 10'd178; a_exp3 = 10'd554;
b_exp0 = 10'd821; b_exp1 = 10'd1006; b_exp2 = 10'd569; b_exp3 = 10'd624;
a_sign0 = 4'd0; a_sign1 = 4'd16; a_sign2 = 4'd14; a_sign3 = 4'd7;
b_sign0 = 4'd15; b_sign1 = 4'd14; b_sign2 = 4'd13; b_sign3 = 4'd1;
@(posedge clk_i);
a_mant0 = 8'd78; a_mant1 = 8'd150; a_mant2 = 8'd169; a_mant3 = 8'd191;
b_mant0 = 8'd187; b_mant1 = 8'd115; b_mant2 = 8'd120; b_mant3 = 8'd169;
a_exp0 = 10'd998; a_exp1 = 10'd1022; a_exp2 = 10'd144; a_exp3 = 10'd775;
b_exp0 = 10'd713; b_exp1 = 10'd245; b_exp2 = 10'd91; b_exp3 = 10'd737;
a_sign0 = 4'd1; a_sign1 = 4'd6; a_sign2 = 4'd15; a_sign3 = 4'd9;
b_sign0 = 4'd12; b_sign1 = 4'd0; b_sign2 = 4'd13; b_sign3 = 4'd2;
@(posedge clk_i);
a_mant0 = 8'd206; a_mant1 = 8'd169; a_mant2 = 8'd86; a_mant3 = 8'd162;
b_mant0 = 8'd216; b_mant1 = 8'd195; b_mant2 = 8'd233; b_mant3 = 8'd245;
a_exp0 = 10'd225; a_exp1 = 10'd405; a_exp2 = 10'd719; a_exp3 = 10'd381;
b_exp0 = 10'd198; b_exp1 = 10'd185; b_exp2 = 10'd565; b_exp3 = 10'd391;
a_sign0 = 4'd9; a_sign1 = 4'd7; a_sign2 = 4'd9; a_sign3 = 4'd10;
b_sign0 = 4'd1; b_sign1 = 4'd5; b_sign2 = 4'd14; b_sign3 = 4'd8;
@(posedge clk_i);
a_mant0 = 8'd223; a_mant1 = 8'd245; a_mant2 = 8'd178; a_mant3 = 8'd168;
b_mant0 = 8'd4; b_mant1 = 8'd197; b_mant2 = 8'd91; b_mant3 = 8'd45;
a_exp0 = 10'd900; a_exp1 = 10'd294; a_exp2 = 10'd585; a_exp3 = 10'd426;
b_exp0 = 10'd162; b_exp1 = 10'd967; b_exp2 = 10'd688; b_exp3 = 10'd331;
a_sign0 = 4'd3; a_sign1 = 4'd1; a_sign2 = 4'd11; a_sign3 = 4'd13;
b_sign0 = 4'd16; b_sign1 = 4'd9; b_sign2 = 4'd13; b_sign3 = 4'd7;
@(posedge clk_i);
shared_exps0 = 8'd125;
shared_exps1 = 8'd152;
a_mant0 = 8'd10; a_mant1 = 8'd23; a_mant2 = 8'd200; a_mant3 = 8'd137;
b_mant0 = 8'd28; b_mant1 = 8'd11; b_mant2 = 8'd88; b_mant3 = 8'd51;
a_exp0 = 10'd211; a_exp1 = 10'd733; a_exp2 = 10'd658; a_exp3 = 10'd841;
b_exp0 = 10'd425; b_exp1 = 10'd542; b_exp2 = 10'd647; b_exp3 = 10'd330;
a_sign0 = 4'd9; a_sign1 = 4'd3; a_sign2 = 4'd2; a_sign3 = 4'd3;
b_sign0 = 4'd7; b_sign1 = 4'd11; b_sign2 = 4'd13; b_sign3 = 4'd9;
@(posedge clk_i);
a_mant0 = 8'd137; a_mant1 = 8'd192; a_mant2 = 8'd205; a_mant3 = 8'd53;
b_mant0 = 8'd42; b_mant1 = 8'd166; b_mant2 = 8'd243; b_mant3 = 8'd40;
a_exp0 = 10'd779; a_exp1 = 10'd406; a_exp2 = 10'd674; a_exp3 = 10'd7;
b_exp0 = 10'd283; b_exp1 = 10'd679; b_exp2 = 10'd689; b_exp3 = 10'd601;
a_sign0 = 4'd12; a_sign1 = 4'd15; a_sign2 = 4'd2; a_sign3 = 4'd13;
b_sign0 = 4'd1; b_sign1 = 4'd11; b_sign2 = 4'd2; b_sign3 = 4'd3;
@(posedge clk_i);
a_mant0 = 8'd223; a_mant1 = 8'd225; a_mant2 = 8'd129; a_mant3 = 8'd220;
b_mant0 = 8'd142; b_mant1 = 8'd132; b_mant2 = 8'd120; b_mant3 = 8'd61;
a_exp0 = 10'd687; a_exp1 = 10'd40; a_exp2 = 10'd875; a_exp3 = 10'd72;
b_exp0 = 10'd462; b_exp1 = 10'd355; b_exp2 = 10'd332; b_exp3 = 10'd191;
a_sign0 = 4'd0; a_sign1 = 4'd8; a_sign2 = 4'd1; a_sign3 = 4'd6;
b_sign0 = 4'd7; b_sign1 = 4'd3; b_sign2 = 4'd14; b_sign3 = 4'd5;
@(posedge clk_i);
a_mant0 = 8'd27; a_mant1 = 8'd96; a_mant2 = 8'd55; a_mant3 = 8'd145;
b_mant0 = 8'd15; b_mant1 = 8'd136; b_mant2 = 8'd85; b_mant3 = 8'd228;
a_exp0 = 10'd151; a_exp1 = 10'd786; a_exp2 = 10'd146; a_exp3 = 10'd210;
b_exp0 = 10'd692; b_exp1 = 10'd189; b_exp2 = 10'd895; b_exp3 = 10'd782;
a_sign0 = 4'd9; a_sign1 = 4'd6; a_sign2 = 4'd5; a_sign3 = 4'd16;
b_sign0 = 4'd5; b_sign1 = 4'd3; b_sign2 = 4'd9; b_sign3 = 4'd6;
@(posedge clk_i);
a_mant0 = 8'd254; a_mant1 = 8'd19; a_mant2 = 8'd159; a_mant3 = 8'd59;
b_mant0 = 8'd216; b_mant1 = 8'd34; b_mant2 = 8'd213; b_mant3 = 8'd32;
a_exp0 = 10'd50; a_exp1 = 10'd387; a_exp2 = 10'd93; a_exp3 = 10'd203;
b_exp0 = 10'd308; b_exp1 = 10'd403; b_exp2 = 10'd1018; b_exp3 = 10'd117;
a_sign0 = 4'd3; a_sign1 = 4'd11; a_sign2 = 4'd4; a_sign3 = 4'd1;
b_sign0 = 4'd9; b_sign1 = 4'd15; b_sign2 = 4'd15; b_sign3 = 4'd9;
@(posedge clk_i);
a_mant0 = 8'd100; a_mant1 = 8'd169; a_mant2 = 8'd212; a_mant3 = 8'd126;
b_mant0 = 8'd188; b_mant1 = 8'd215; b_mant2 = 8'd89; b_mant3 = 8'd11;
a_exp0 = 10'd697; a_exp1 = 10'd923; a_exp2 = 10'd836; a_exp3 = 10'd607;
b_exp0 = 10'd984; b_exp1 = 10'd368; b_exp2 = 10'd993; b_exp3 = 10'd717;
a_sign0 = 4'd13; a_sign1 = 4'd2; a_sign2 = 4'd10; a_sign3 = 4'd2;
b_sign0 = 4'd1; b_sign1 = 4'd16; b_sign2 = 4'd12; b_sign3 = 4'd4;
@(posedge clk_i);
a_mant0 = 8'd88; a_mant1 = 8'd2; a_mant2 = 8'd174; a_mant3 = 8'd76;
b_mant0 = 8'd193; b_mant1 = 8'd252; b_mant2 = 8'd107; b_mant3 = 8'd0;
a_exp0 = 10'd387; a_exp1 = 10'd664; a_exp2 = 10'd922; a_exp3 = 10'd167;
b_exp0 = 10'd889; b_exp1 = 10'd66; b_exp2 = 10'd165; b_exp3 = 10'd245;
a_sign0 = 4'd3; a_sign1 = 4'd3; a_sign2 = 4'd10; a_sign3 = 4'd13;
b_sign0 = 4'd2; b_sign1 = 4'd3; b_sign2 = 4'd12; b_sign3 = 4'd7;
@(posedge clk_i);
a_mant0 = 8'd242; a_mant1 = 8'd124; a_mant2 = 8'd207; a_mant3 = 8'd40;
b_mant0 = 8'd241; b_mant1 = 8'd63; b_mant2 = 8'd159; b_mant3 = 8'd42;
a_exp0 = 10'd753; a_exp1 = 10'd385; a_exp2 = 10'd846; a_exp3 = 10'd216;
b_exp0 = 10'd859; b_exp1 = 10'd752; b_exp2 = 10'd105; b_exp3 = 10'd250;
a_sign0 = 4'd12; a_sign1 = 4'd11; a_sign2 = 4'd12; a_sign3 = 4'd5;
b_sign0 = 4'd1; b_sign1 = 4'd10; b_sign2 = 4'd7; b_sign3 = 4'd7;
@(posedge clk_i);
shared_exps0 = 8'd137;
shared_exps1 = 8'd138;
a_mant0 = 8'd211; a_mant1 = 8'd80; a_mant2 = 8'd212; a_mant3 = 8'd226;
b_mant0 = 8'd29; b_mant1 = 8'd168; b_mant2 = 8'd52; b_mant3 = 8'd244;
a_exp0 = 10'd759; a_exp1 = 10'd702; a_exp2 = 10'd620; a_exp3 = 10'd516;
b_exp0 = 10'd323; b_exp1 = 10'd616; b_exp2 = 10'd38; b_exp3 = 10'd689;
a_sign0 = 4'd7; a_sign1 = 4'd8; a_sign2 = 4'd1; a_sign3 = 4'd11;
b_sign0 = 4'd10; b_sign1 = 4'd7; b_sign2 = 4'd8; b_sign3 = 4'd6;
@(posedge clk_i);
a_mant0 = 8'd233; a_mant1 = 8'd232; a_mant2 = 8'd0; a_mant3 = 8'd54;
b_mant0 = 8'd123; b_mant1 = 8'd115; b_mant2 = 8'd112; b_mant3 = 8'd251;
a_exp0 = 10'd393; a_exp1 = 10'd521; a_exp2 = 10'd83; a_exp3 = 10'd712;
b_exp0 = 10'd83; b_exp1 = 10'd676; b_exp2 = 10'd916; b_exp3 = 10'd288;
a_sign0 = 4'd16; a_sign1 = 4'd7; a_sign2 = 4'd5; a_sign3 = 4'd6;
b_sign0 = 4'd4; b_sign1 = 4'd12; b_sign2 = 4'd15; b_sign3 = 4'd14;
@(posedge clk_i);
a_mant0 = 8'd54; a_mant1 = 8'd113; a_mant2 = 8'd79; a_mant3 = 8'd6;
b_mant0 = 8'd169; b_mant1 = 8'd71; b_mant2 = 8'd186; b_mant3 = 8'd215;
a_exp0 = 10'd453; a_exp1 = 10'd965; a_exp2 = 10'd717; a_exp3 = 10'd758;
b_exp0 = 10'd797; b_exp1 = 10'd834; b_exp2 = 10'd986; b_exp3 = 10'd573;
a_sign0 = 4'd5; a_sign1 = 4'd12; a_sign2 = 4'd7; a_sign3 = 4'd14;
b_sign0 = 4'd14; b_sign1 = 4'd7; b_sign2 = 4'd15; b_sign3 = 4'd4;
@(posedge clk_i);
a_mant0 = 8'd3; a_mant1 = 8'd165; a_mant2 = 8'd98; a_mant3 = 8'd106;
b_mant0 = 8'd239; b_mant1 = 8'd250; b_mant2 = 8'd220; b_mant3 = 8'd7;
a_exp0 = 10'd633; a_exp1 = 10'd373; a_exp2 = 10'd723; a_exp3 = 10'd892;
b_exp0 = 10'd399; b_exp1 = 10'd9; b_exp2 = 10'd843; b_exp3 = 10'd419;
a_sign0 = 4'd5; a_sign1 = 4'd2; a_sign2 = 4'd0; a_sign3 = 4'd11;
b_sign0 = 4'd7; b_sign1 = 4'd16; b_sign2 = 4'd3; b_sign3 = 4'd15;
@(posedge clk_i);
a_mant0 = 8'd3; a_mant1 = 8'd251; a_mant2 = 8'd108; a_mant3 = 8'd40;
b_mant0 = 8'd203; b_mant1 = 8'd60; b_mant2 = 8'd182; b_mant3 = 8'd132;
a_exp0 = 10'd631; a_exp1 = 10'd274; a_exp2 = 10'd689; a_exp3 = 10'd1006;
b_exp0 = 10'd957; b_exp1 = 10'd723; b_exp2 = 10'd111; b_exp3 = 10'd181;
a_sign0 = 4'd10; a_sign1 = 4'd11; a_sign2 = 4'd4; a_sign3 = 4'd4;
b_sign0 = 4'd6; b_sign1 = 4'd0; b_sign2 = 4'd16; b_sign3 = 4'd10;
@(posedge clk_i);
a_mant0 = 8'd215; a_mant1 = 8'd191; a_mant2 = 8'd175; a_mant3 = 8'd175;
b_mant0 = 8'd3; b_mant1 = 8'd150; b_mant2 = 8'd230; b_mant3 = 8'd188;
a_exp0 = 10'd437; a_exp1 = 10'd484; a_exp2 = 10'd867; a_exp3 = 10'd98;
b_exp0 = 10'd647; b_exp1 = 10'd375; b_exp2 = 10'd3; b_exp3 = 10'd360;
a_sign0 = 4'd8; a_sign1 = 4'd4; a_sign2 = 4'd3; a_sign3 = 4'd12;
b_sign0 = 4'd3; b_sign1 = 4'd0; b_sign2 = 4'd1; b_sign3 = 4'd14;
@(posedge clk_i);
a_mant0 = 8'd132; a_mant1 = 8'd121; a_mant2 = 8'd216; a_mant3 = 8'd150;
b_mant0 = 8'd205; b_mant1 = 8'd68; b_mant2 = 8'd97; b_mant3 = 8'd60;
a_exp0 = 10'd470; a_exp1 = 10'd68; a_exp2 = 10'd503; a_exp3 = 10'd258;
b_exp0 = 10'd226; b_exp1 = 10'd481; b_exp2 = 10'd816; b_exp3 = 10'd755;
a_sign0 = 4'd6; a_sign1 = 4'd9; a_sign2 = 4'd9; a_sign3 = 4'd7;
b_sign0 = 4'd1; b_sign1 = 4'd0; b_sign2 = 4'd12; b_sign3 = 4'd4;
@(posedge clk_i);
a_mant0 = 8'd245; a_mant1 = 8'd227; a_mant2 = 8'd133; a_mant3 = 8'd146;
b_mant0 = 8'd245; b_mant1 = 8'd99; b_mant2 = 8'd31; b_mant3 = 8'd46;
a_exp0 = 10'd469; a_exp1 = 10'd161; a_exp2 = 10'd674; a_exp3 = 10'd884;
b_exp0 = 10'd509; b_exp1 = 10'd598; b_exp2 = 10'd706; b_exp3 = 10'd217;
a_sign0 = 4'd10; a_sign1 = 4'd2; a_sign2 = 4'd0; a_sign3 = 4'd2;
b_sign0 = 4'd11; b_sign1 = 4'd14; b_sign2 = 4'd0; b_sign3 = 4'd2;
@(posedge clk_i);
shared_exps0 = 8'd90;
shared_exps1 = 8'd138;
a_mant0 = 8'd109; a_mant1 = 8'd27; a_mant2 = 8'd145; a_mant3 = 8'd234;
b_mant0 = 8'd88; b_mant1 = 8'd68; b_mant2 = 8'd186; b_mant3 = 8'd48;
a_exp0 = 10'd254; a_exp1 = 10'd591; a_exp2 = 10'd8; a_exp3 = 10'd713;
b_exp0 = 10'd285; b_exp1 = 10'd64; b_exp2 = 10'd791; b_exp3 = 10'd276;
a_sign0 = 4'd11; a_sign1 = 4'd3; a_sign2 = 4'd6; a_sign3 = 4'd7;
b_sign0 = 4'd6; b_sign1 = 4'd11; b_sign2 = 4'd15; b_sign3 = 4'd13;
@(posedge clk_i);
a_mant0 = 8'd90; a_mant1 = 8'd76; a_mant2 = 8'd115; a_mant3 = 8'd62;
b_mant0 = 8'd153; b_mant1 = 8'd170; b_mant2 = 8'd174; b_mant3 = 8'd173;
a_exp0 = 10'd181; a_exp1 = 10'd109; a_exp2 = 10'd910; a_exp3 = 10'd684;
b_exp0 = 10'd128; b_exp1 = 10'd528; b_exp2 = 10'd438; b_exp3 = 10'd838;
a_sign0 = 4'd9; a_sign1 = 4'd0; a_sign2 = 4'd16; a_sign3 = 4'd9;
b_sign0 = 4'd1; b_sign1 = 4'd12; b_sign2 = 4'd15; b_sign3 = 4'd8;
@(posedge clk_i);
a_mant0 = 8'd215; a_mant1 = 8'd34; a_mant2 = 8'd101; a_mant3 = 8'd253;
b_mant0 = 8'd185; b_mant1 = 8'd147; b_mant2 = 8'd142; b_mant3 = 8'd55;
a_exp0 = 10'd85; a_exp1 = 10'd425; a_exp2 = 10'd772; a_exp3 = 10'd245;
b_exp0 = 10'd931; b_exp1 = 10'd104; b_exp2 = 10'd289; b_exp3 = 10'd717;
a_sign0 = 4'd16; a_sign1 = 4'd1; a_sign2 = 4'd16; a_sign3 = 4'd8;
b_sign0 = 4'd10; b_sign1 = 4'd1; b_sign2 = 4'd11; b_sign3 = 4'd16;
@(posedge clk_i);
a_mant0 = 8'd164; a_mant1 = 8'd86; a_mant2 = 8'd201; a_mant3 = 8'd160;
b_mant0 = 8'd244; b_mant1 = 8'd90; b_mant2 = 8'd39; b_mant3 = 8'd202;
a_exp0 = 10'd551; a_exp1 = 10'd698; a_exp2 = 10'd787; a_exp3 = 10'd792;
b_exp0 = 10'd828; b_exp1 = 10'd70; b_exp2 = 10'd800; b_exp3 = 10'd553;
a_sign0 = 4'd2; a_sign1 = 4'd14; a_sign2 = 4'd16; a_sign3 = 4'd4;
b_sign0 = 4'd4; b_sign1 = 4'd7; b_sign2 = 4'd7; b_sign3 = 4'd11;
@(posedge clk_i);
a_mant0 = 8'd227; a_mant1 = 8'd139; a_mant2 = 8'd40; a_mant3 = 8'd201;
b_mant0 = 8'd31; b_mant1 = 8'd207; b_mant2 = 8'd242; b_mant3 = 8'd241;
a_exp0 = 10'd716; a_exp1 = 10'd571; a_exp2 = 10'd777; a_exp3 = 10'd616;
b_exp0 = 10'd534; b_exp1 = 10'd89; b_exp2 = 10'd743; b_exp3 = 10'd248;
a_sign0 = 4'd4; a_sign1 = 4'd3; a_sign2 = 4'd5; a_sign3 = 4'd0;
b_sign0 = 4'd5; b_sign1 = 4'd12; b_sign2 = 4'd11; b_sign3 = 4'd12;
@(posedge clk_i);
a_mant0 = 8'd69; a_mant1 = 8'd177; a_mant2 = 8'd204; a_mant3 = 8'd122;
b_mant0 = 8'd63; b_mant1 = 8'd7; b_mant2 = 8'd158; b_mant3 = 8'd238;
a_exp0 = 10'd242; a_exp1 = 10'd537; a_exp2 = 10'd470; a_exp3 = 10'd961;
b_exp0 = 10'd864; b_exp1 = 10'd685; b_exp2 = 10'd839; b_exp3 = 10'd187;
a_sign0 = 4'd7; a_sign1 = 4'd4; a_sign2 = 4'd14; a_sign3 = 4'd12;
b_sign0 = 4'd8; b_sign1 = 4'd4; b_sign2 = 4'd7; b_sign3 = 4'd13;
@(posedge clk_i);
a_mant0 = 8'd20; a_mant1 = 8'd128; a_mant2 = 8'd21; a_mant3 = 8'd145;
b_mant0 = 8'd231; b_mant1 = 8'd225; b_mant2 = 8'd21; b_mant3 = 8'd121;
a_exp0 = 10'd670; a_exp1 = 10'd101; a_exp2 = 10'd438; a_exp3 = 10'd173;
b_exp0 = 10'd883; b_exp1 = 10'd294; b_exp2 = 10'd626; b_exp3 = 10'd545;
a_sign0 = 4'd4; a_sign1 = 4'd16; a_sign2 = 4'd7; a_sign3 = 4'd9;
b_sign0 = 4'd0; b_sign1 = 4'd11; b_sign2 = 4'd5; b_sign3 = 4'd11;
@(posedge clk_i);
a_mant0 = 8'd107; a_mant1 = 8'd205; a_mant2 = 8'd37; a_mant3 = 8'd33;
b_mant0 = 8'd182; b_mant1 = 8'd113; b_mant2 = 8'd189; b_mant3 = 8'd84;
a_exp0 = 10'd525; a_exp1 = 10'd510; a_exp2 = 10'd795; a_exp3 = 10'd30;
b_exp0 = 10'd837; b_exp1 = 10'd186; b_exp2 = 10'd332; b_exp3 = 10'd638;
a_sign0 = 4'd1; a_sign1 = 4'd0; a_sign2 = 4'd10; a_sign3 = 4'd4;
b_sign0 = 4'd2; b_sign1 = 4'd8; b_sign2 = 4'd0; b_sign3 = 4'd13;
@(posedge clk_i);
shared_exps0 = 8'd143;
shared_exps1 = 8'd102;
rstn = 0;
@(posedge clk_i);
rstn = 1;
a_mant0 = 8'd141; a_mant1 = 8'd147; a_mant2 = 8'd52; a_mant3 = 8'd66;
b_mant0 = 8'd85; b_mant1 = 8'd22; b_mant2 = 8'd87; b_mant3 = 8'd69;
a_exp0 = 10'd77; a_exp1 = 10'd925; a_exp2 = 10'd422; a_exp3 = 10'd695;
b_exp0 = 10'd24; b_exp1 = 10'd1000; b_exp2 = 10'd201; b_exp3 = 10'd743;
a_sign0 = 4'd1; a_sign1 = 4'd2; a_sign2 = 4'd15; a_sign3 = 4'd15;
b_sign0 = 4'd8; b_sign1 = 4'd6; b_sign2 = 4'd16; b_sign3 = 4'd14;
@(posedge clk_i);
a_mant0 = 8'd238; a_mant1 = 8'd136; a_mant2 = 8'd204; a_mant3 = 8'd224;
b_mant0 = 8'd99; b_mant1 = 8'd21; b_mant2 = 8'd6; b_mant3 = 8'd73;
a_exp0 = 10'd972; a_exp1 = 10'd43; a_exp2 = 10'd920; a_exp3 = 10'd876;
b_exp0 = 10'd433; b_exp1 = 10'd812; b_exp2 = 10'd462; b_exp3 = 10'd752;
a_sign0 = 4'd0; a_sign1 = 4'd15; a_sign2 = 4'd9; a_sign3 = 4'd14;
b_sign0 = 4'd0; b_sign1 = 4'd2; b_sign2 = 4'd13; b_sign3 = 4'd8;
@(posedge clk_i);
a_mant0 = 8'd251; a_mant1 = 8'd187; a_mant2 = 8'd65; a_mant3 = 8'd216;
b_mant0 = 8'd91; b_mant1 = 8'd134; b_mant2 = 8'd78; b_mant3 = 8'd207;
a_exp0 = 10'd333; a_exp1 = 10'd943; a_exp2 = 10'd551; a_exp3 = 10'd133;
b_exp0 = 10'd995; b_exp1 = 10'd611; b_exp2 = 10'd530; b_exp3 = 10'd460;
a_sign0 = 4'd13; a_sign1 = 4'd9; a_sign2 = 4'd16; a_sign3 = 4'd4;
b_sign0 = 4'd10; b_sign1 = 4'd1; b_sign2 = 4'd14; b_sign3 = 4'd7;
@(posedge clk_i);
a_mant0 = 8'd186; a_mant1 = 8'd148; a_mant2 = 8'd55; a_mant3 = 8'd251;
b_mant0 = 8'd151; b_mant1 = 8'd97; b_mant2 = 8'd185; b_mant3 = 8'd174;
a_exp0 = 10'd578; a_exp1 = 10'd491; a_exp2 = 10'd274; a_exp3 = 10'd52;
b_exp0 = 10'd589; b_exp1 = 10'd901; b_exp2 = 10'd799; b_exp3 = 10'd1023;
a_sign0 = 4'd7; a_sign1 = 4'd11; a_sign2 = 4'd1; a_sign3 = 4'd16;
b_sign0 = 4'd2; b_sign1 = 4'd12; b_sign2 = 4'd4; b_sign3 = 4'd10;
@(posedge clk_i);
a_mant0 = 8'd55; a_mant1 = 8'd252; a_mant2 = 8'd60; a_mant3 = 8'd71;
b_mant0 = 8'd78; b_mant1 = 8'd156; b_mant2 = 8'd173; b_mant3 = 8'd101;
a_exp0 = 10'd401; a_exp1 = 10'd39; a_exp2 = 10'd894; a_exp3 = 10'd187;
b_exp0 = 10'd668; b_exp1 = 10'd820; b_exp2 = 10'd36; b_exp3 = 10'd406;
a_sign0 = 4'd9; a_sign1 = 4'd6; a_sign2 = 4'd5; a_sign3 = 4'd9;
b_sign0 = 4'd16; b_sign1 = 4'd10; b_sign2 = 4'd2; b_sign3 = 4'd0;
@(posedge clk_i);
a_mant0 = 8'd233; a_mant1 = 8'd219; a_mant2 = 8'd175; a_mant3 = 8'd104;
b_mant0 = 8'd4; b_mant1 = 8'd96; b_mant2 = 8'd95; b_mant3 = 8'd209;
a_exp0 = 10'd768; a_exp1 = 10'd714; a_exp2 = 10'd619; a_exp3 = 10'd855;
b_exp0 = 10'd96; b_exp1 = 10'd500; b_exp2 = 10'd849; b_exp3 = 10'd347;
a_sign0 = 4'd3; a_sign1 = 4'd15; a_sign2 = 4'd7; a_sign3 = 4'd9;
b_sign0 = 4'd2; b_sign1 = 4'd8; b_sign2 = 4'd14; b_sign3 = 4'd9;
@(posedge clk_i);
a_mant0 = 8'd157; a_mant1 = 8'd243; a_mant2 = 8'd75; a_mant3 = 8'd34;
b_mant0 = 8'd99; b_mant1 = 8'd7; b_mant2 = 8'd145; b_mant3 = 8'd170;
a_exp0 = 10'd366; a_exp1 = 10'd55; a_exp2 = 10'd910; a_exp3 = 10'd882;
b_exp0 = 10'd786; b_exp1 = 10'd327; b_exp2 = 10'd814; b_exp3 = 10'd58;
a_sign0 = 4'd13; a_sign1 = 4'd10; a_sign2 = 4'd1; a_sign3 = 4'd12;
b_sign0 = 4'd3; b_sign1 = 4'd9; b_sign2 = 4'd5; b_sign3 = 4'd6;
@(posedge clk_i);
shared_exps0 = 8'd132;
shared_exps1 = 8'd129;
a_mant0 = 8'd54; a_mant1 = 8'd137; a_mant2 = 8'd48; a_mant3 = 8'd142;
b_mant0 = 8'd62; b_mant1 = 8'd84; b_mant2 = 8'd96; b_mant3 = 8'd231;
a_exp0 = 10'd435; a_exp1 = 10'd911; a_exp2 = 10'd329; a_exp3 = 10'd330;
b_exp0 = 10'd717; b_exp1 = 10'd366; b_exp2 = 10'd329; b_exp3 = 10'd760;
a_sign0 = 4'd7; a_sign1 = 4'd0; a_sign2 = 4'd9; a_sign3 = 4'd0;
b_sign0 = 4'd2; b_sign1 = 4'd8; b_sign2 = 4'd16; b_sign3 = 4'd1;
@(posedge clk_i);
a_mant0 = 8'd90; a_mant1 = 8'd138; a_mant2 = 8'd212; a_mant3 = 8'd128;
b_mant0 = 8'd112; b_mant1 = 8'd195; b_mant2 = 8'd0; b_mant3 = 8'd220;
a_exp0 = 10'd679; a_exp1 = 10'd365; a_exp2 = 10'd411; a_exp3 = 10'd531;
b_exp0 = 10'd106; b_exp1 = 10'd612; b_exp2 = 10'd1001; b_exp3 = 10'd178;
a_sign0 = 4'd4; a_sign1 = 4'd4; a_sign2 = 4'd4; a_sign3 = 4'd6;
b_sign0 = 4'd2; b_sign1 = 4'd1; b_sign2 = 4'd12; b_sign3 = 4'd10;
@(posedge clk_i);
a_mant0 = 8'd81; a_mant1 = 8'd177; a_mant2 = 8'd40; a_mant3 = 8'd84;
b_mant0 = 8'd186; b_mant1 = 8'd164; b_mant2 = 8'd132; b_mant3 = 8'd10;
a_exp0 = 10'd932; a_exp1 = 10'd589; a_exp2 = 10'd783; a_exp3 = 10'd225;
b_exp0 = 10'd157; b_exp1 = 10'd327; b_exp2 = 10'd195; b_exp3 = 10'd416;
a_sign0 = 4'd3; a_sign1 = 4'd10; a_sign2 = 4'd10; a_sign3 = 4'd3;
b_sign0 = 4'd3; b_sign1 = 4'd6; b_sign2 = 4'd8; b_sign3 = 4'd2;
@(posedge clk_i);
a_mant0 = 8'd115; a_mant1 = 8'd176; a_mant2 = 8'd216; a_mant3 = 8'd170;
b_mant0 = 8'd50; b_mant1 = 8'd121; b_mant2 = 8'd109; b_mant3 = 8'd46;
a_exp0 = 10'd88; a_exp1 = 10'd245; a_exp2 = 10'd721; a_exp3 = 10'd511;
b_exp0 = 10'd86; b_exp1 = 10'd977; b_exp2 = 10'd600; b_exp3 = 10'd996;
a_sign0 = 4'd5; a_sign1 = 4'd2; a_sign2 = 4'd6; a_sign3 = 4'd12;
b_sign0 = 4'd9; b_sign1 = 4'd0; b_sign2 = 4'd2; b_sign3 = 4'd6;
@(posedge clk_i);
a_mant0 = 8'd140; a_mant1 = 8'd136; a_mant2 = 8'd170; a_mant3 = 8'd178;
b_mant0 = 8'd54; b_mant1 = 8'd56; b_mant2 = 8'd143; b_mant3 = 8'd70;
a_exp0 = 10'd462; a_exp1 = 10'd337; a_exp2 = 10'd64; a_exp3 = 10'd86;
b_exp0 = 10'd563; b_exp1 = 10'd84; b_exp2 = 10'd236; b_exp3 = 10'd795;
a_sign0 = 4'd1; a_sign1 = 4'd14; a_sign2 = 4'd0; a_sign3 = 4'd1;
b_sign0 = 4'd13; b_sign1 = 4'd1; b_sign2 = 4'd3; b_sign3 = 4'd6;
@(posedge clk_i);
a_mant0 = 8'd237; a_mant1 = 8'd178; a_mant2 = 8'd228; a_mant3 = 8'd32;
b_mant0 = 8'd250; b_mant1 = 8'd165; b_mant2 = 8'd244; b_mant3 = 8'd106;
a_exp0 = 10'd341; a_exp1 = 10'd667; a_exp2 = 10'd307; a_exp3 = 10'd59;
b_exp0 = 10'd181; b_exp1 = 10'd844; b_exp2 = 10'd376; b_exp3 = 10'd374;
a_sign0 = 4'd14; a_sign1 = 4'd13; a_sign2 = 4'd10; a_sign3 = 4'd5;
b_sign0 = 4'd13; b_sign1 = 4'd12; b_sign2 = 4'd0; b_sign3 = 4'd3;
@(posedge clk_i);
a_mant0 = 8'd70; a_mant1 = 8'd16; a_mant2 = 8'd103; a_mant3 = 8'd58;
b_mant0 = 8'd120; b_mant1 = 8'd156; b_mant2 = 8'd129; b_mant3 = 8'd3;
a_exp0 = 10'd928; a_exp1 = 10'd258; a_exp2 = 10'd712; a_exp3 = 10'd694;
b_exp0 = 10'd830; b_exp1 = 10'd635; b_exp2 = 10'd346; b_exp3 = 10'd610;
a_sign0 = 4'd15; a_sign1 = 4'd11; a_sign2 = 4'd2; a_sign3 = 4'd16;
b_sign0 = 4'd5; b_sign1 = 4'd9; b_sign2 = 4'd7; b_sign3 = 4'd11;
@(posedge clk_i);
a_mant0 = 8'd34; a_mant1 = 8'd190; a_mant2 = 8'd96; a_mant3 = 8'd246;
b_mant0 = 8'd98; b_mant1 = 8'd9; b_mant2 = 8'd95; b_mant3 = 8'd252;
a_exp0 = 10'd314; a_exp1 = 10'd476; a_exp2 = 10'd998; a_exp3 = 10'd806;
b_exp0 = 10'd487; b_exp1 = 10'd809; b_exp2 = 10'd496; b_exp3 = 10'd23;
a_sign0 = 4'd4; a_sign1 = 4'd11; a_sign2 = 4'd5; a_sign3 = 4'd12;
b_sign0 = 4'd13; b_sign1 = 4'd6; b_sign2 = 4'd2; b_sign3 = 4'd12;
@(posedge clk_i);
shared_exps0 = 8'd143;
shared_exps1 = 8'd131;
a_mant0 = 8'd165; a_mant1 = 8'd99; a_mant2 = 8'd72; a_mant3 = 8'd161;
b_mant0 = 8'd72; b_mant1 = 8'd211; b_mant2 = 8'd65; b_mant3 = 8'd5;
a_exp0 = 10'd555; a_exp1 = 10'd548; a_exp2 = 10'd727; a_exp3 = 10'd736;
b_exp0 = 10'd791; b_exp1 = 10'd258; b_exp2 = 10'd997; b_exp3 = 10'd140;
a_sign0 = 4'd3; a_sign1 = 4'd13; a_sign2 = 4'd4; a_sign3 = 4'd10;
b_sign0 = 4'd8; b_sign1 = 4'd5; b_sign2 = 4'd3; b_sign3 = 4'd16;
@(posedge clk_i);
a_mant0 = 8'd8; a_mant1 = 8'd138; a_mant2 = 8'd19; a_mant3 = 8'd191;
b_mant0 = 8'd226; b_mant1 = 8'd132; b_mant2 = 8'd25; b_mant3 = 8'd236;
a_exp0 = 10'd165; a_exp1 = 10'd582; a_exp2 = 10'd765; a_exp3 = 10'd361;
b_exp0 = 10'd103; b_exp1 = 10'd603; b_exp2 = 10'd756; b_exp3 = 10'd224;
a_sign0 = 4'd13; a_sign1 = 4'd8; a_sign2 = 4'd1; a_sign3 = 4'd16;
b_sign0 = 4'd6; b_sign1 = 4'd3; b_sign2 = 4'd6; b_sign3 = 4'd8;
@(posedge clk_i);
a_mant0 = 8'd22; a_mant1 = 8'd223; a_mant2 = 8'd16; a_mant3 = 8'd238;
b_mant0 = 8'd213; b_mant1 = 8'd83; b_mant2 = 8'd185; b_mant3 = 8'd149;
a_exp0 = 10'd853; a_exp1 = 10'd694; a_exp2 = 10'd219; a_exp3 = 10'd617;
b_exp0 = 10'd829; b_exp1 = 10'd316; b_exp2 = 10'd536; b_exp3 = 10'd869;
a_sign0 = 4'd13; a_sign1 = 4'd8; a_sign2 = 4'd5; a_sign3 = 4'd2;
b_sign0 = 4'd3; b_sign1 = 4'd15; b_sign2 = 4'd5; b_sign3 = 4'd4;
@(posedge clk_i);
a_mant0 = 8'd86; a_mant1 = 8'd7; a_mant2 = 8'd111; a_mant3 = 8'd76;
b_mant0 = 8'd191; b_mant1 = 8'd6; b_mant2 = 8'd226; b_mant3 = 8'd59;
a_exp0 = 10'd621; a_exp1 = 10'd839; a_exp2 = 10'd327; a_exp3 = 10'd265;
b_exp0 = 10'd617; b_exp1 = 10'd697; b_exp2 = 10'd292; b_exp3 = 10'd992;
a_sign0 = 4'd5; a_sign1 = 4'd3; a_sign2 = 4'd12; a_sign3 = 4'd1;
b_sign0 = 4'd10; b_sign1 = 4'd16; b_sign2 = 4'd10; b_sign3 = 4'd10;
@(posedge clk_i);
a_mant0 = 8'd54; a_mant1 = 8'd51; a_mant2 = 8'd179; a_mant3 = 8'd223;
b_mant0 = 8'd243; b_mant1 = 8'd17; b_mant2 = 8'd5; b_mant3 = 8'd39;
a_exp0 = 10'd486; a_exp1 = 10'd1000; a_exp2 = 10'd392; a_exp3 = 10'd488;
b_exp0 = 10'd952; b_exp1 = 10'd477; b_exp2 = 10'd920; b_exp3 = 10'd289;
a_sign0 = 4'd2; a_sign1 = 4'd0; a_sign2 = 4'd13; a_sign3 = 4'd13;
b_sign0 = 4'd1; b_sign1 = 4'd1; b_sign2 = 4'd4; b_sign3 = 4'd12;
@(posedge clk_i);
a_mant0 = 8'd99; a_mant1 = 8'd169; a_mant2 = 8'd248; a_mant3 = 8'd70;
b_mant0 = 8'd34; b_mant1 = 8'd27; b_mant2 = 8'd86; b_mant3 = 8'd175;
a_exp0 = 10'd1009; a_exp1 = 10'd493; a_exp2 = 10'd481; a_exp3 = 10'd362;
b_exp0 = 10'd825; b_exp1 = 10'd345; b_exp2 = 10'd474; b_exp3 = 10'd643;
a_sign0 = 4'd11; a_sign1 = 4'd1; a_sign2 = 4'd14; a_sign3 = 4'd9;
b_sign0 = 4'd12; b_sign1 = 4'd10; b_sign2 = 4'd7; b_sign3 = 4'd16;
@(posedge clk_i);
a_mant0 = 8'd26; a_mant1 = 8'd140; a_mant2 = 8'd53; a_mant3 = 8'd2;
b_mant0 = 8'd169; b_mant1 = 8'd112; b_mant2 = 8'd197; b_mant3 = 8'd5;
a_exp0 = 10'd731; a_exp1 = 10'd351; a_exp2 = 10'd287; a_exp3 = 10'd993;
b_exp0 = 10'd719; b_exp1 = 10'd408; b_exp2 = 10'd701; b_exp3 = 10'd431;
a_sign0 = 4'd8; a_sign1 = 4'd0; a_sign2 = 4'd5; a_sign3 = 4'd14;
b_sign0 = 4'd13; b_sign1 = 4'd7; b_sign2 = 4'd13; b_sign3 = 4'd15;
@(posedge clk_i);
a_mant0 = 8'd224; a_mant1 = 8'd93; a_mant2 = 8'd209; a_mant3 = 8'd204;
b_mant0 = 8'd95; b_mant1 = 8'd203; b_mant2 = 8'd192; b_mant3 = 8'd54;
a_exp0 = 10'd990; a_exp1 = 10'd866; a_exp2 = 10'd217; a_exp3 = 10'd818;
b_exp0 = 10'd588; b_exp1 = 10'd266; b_exp2 = 10'd432; b_exp3 = 10'd823;
a_sign0 = 4'd15; a_sign1 = 4'd6; a_sign2 = 4'd16; a_sign3 = 4'd15;
b_sign0 = 4'd3; b_sign1 = 4'd2; b_sign2 = 4'd16; b_sign3 = 4'd13;
@(posedge clk_i);
shared_exps0 = 8'd110;
shared_exps1 = 8'd132;
a_mant0 = 8'd80; a_mant1 = 8'd137; a_mant2 = 8'd99; a_mant3 = 8'd21;
b_mant0 = 8'd206; b_mant1 = 8'd207; b_mant2 = 8'd84; b_mant3 = 8'd72;
a_exp0 = 10'd411; a_exp1 = 10'd967; a_exp2 = 10'd645; a_exp3 = 10'd285;
b_exp0 = 10'd676; b_exp1 = 10'd525; b_exp2 = 10'd581; b_exp3 = 10'd696;
a_sign0 = 4'd5; a_sign1 = 4'd7; a_sign2 = 4'd14; a_sign3 = 4'd9;
b_sign0 = 4'd8; b_sign1 = 4'd1; b_sign2 = 4'd13; b_sign3 = 4'd10;
@(posedge clk_i);
a_mant0 = 8'd183; a_mant1 = 8'd97; a_mant2 = 8'd247; a_mant3 = 8'd150;
b_mant0 = 8'd9; b_mant1 = 8'd89; b_mant2 = 8'd186; b_mant3 = 8'd252;
a_exp0 = 10'd160; a_exp1 = 10'd365; a_exp2 = 10'd380; a_exp3 = 10'd419;
b_exp0 = 10'd834; b_exp1 = 10'd337; b_exp2 = 10'd738; b_exp3 = 10'd309;
a_sign0 = 4'd12; a_sign1 = 4'd9; a_sign2 = 4'd13; a_sign3 = 4'd15;
b_sign0 = 4'd7; b_sign1 = 4'd10; b_sign2 = 4'd12; b_sign3 = 4'd14;
@(posedge clk_i);
a_mant0 = 8'd91; a_mant1 = 8'd110; a_mant2 = 8'd54; a_mant3 = 8'd147;
b_mant0 = 8'd151; b_mant1 = 8'd139; b_mant2 = 8'd166; b_mant3 = 8'd183;
a_exp0 = 10'd563; a_exp1 = 10'd723; a_exp2 = 10'd865; a_exp3 = 10'd924;
b_exp0 = 10'd1019; b_exp1 = 10'd168; b_exp2 = 10'd519; b_exp3 = 10'd649;
a_sign0 = 4'd3; a_sign1 = 4'd13; a_sign2 = 4'd15; a_sign3 = 4'd13;
b_sign0 = 4'd13; b_sign1 = 4'd1; b_sign2 = 4'd9; b_sign3 = 4'd8;
@(posedge clk_i);
a_mant0 = 8'd23; a_mant1 = 8'd139; a_mant2 = 8'd14; a_mant3 = 8'd14;
b_mant0 = 8'd90; b_mant1 = 8'd84; b_mant2 = 8'd1; b_mant3 = 8'd125;
a_exp0 = 10'd955; a_exp1 = 10'd489; a_exp2 = 10'd236; a_exp3 = 10'd944;
b_exp0 = 10'd826; b_exp1 = 10'd659; b_exp2 = 10'd485; b_exp3 = 10'd648;
a_sign0 = 4'd4; a_sign1 = 4'd16; a_sign2 = 4'd13; a_sign3 = 4'd6;
b_sign0 = 4'd3; b_sign1 = 4'd12; b_sign2 = 4'd3; b_sign3 = 4'd13;
@(posedge clk_i);
a_mant0 = 8'd69; a_mant1 = 8'd96; a_mant2 = 8'd181; a_mant3 = 8'd214;
b_mant0 = 8'd73; b_mant1 = 8'd187; b_mant2 = 8'd138; b_mant3 = 8'd87;
a_exp0 = 10'd643; a_exp1 = 10'd916; a_exp2 = 10'd497; a_exp3 = 10'd834;
b_exp0 = 10'd1004; b_exp1 = 10'd978; b_exp2 = 10'd752; b_exp3 = 10'd487;
a_sign0 = 4'd7; a_sign1 = 4'd3; a_sign2 = 4'd13; a_sign3 = 4'd11;
b_sign0 = 4'd2; b_sign1 = 4'd2; b_sign2 = 4'd12; b_sign3 = 4'd4;
@(posedge clk_i);
a_mant0 = 8'd74; a_mant1 = 8'd184; a_mant2 = 8'd90; a_mant3 = 8'd15;
b_mant0 = 8'd250; b_mant1 = 8'd46; b_mant2 = 8'd149; b_mant3 = 8'd106;
a_exp0 = 10'd395; a_exp1 = 10'd572; a_exp2 = 10'd628; a_exp3 = 10'd132;
b_exp0 = 10'd132; b_exp1 = 10'd896; b_exp2 = 10'd521; b_exp3 = 10'd922;
a_sign0 = 4'd0; a_sign1 = 4'd7; a_sign2 = 4'd8; a_sign3 = 4'd12;
b_sign0 = 4'd16; b_sign1 = 4'd10; b_sign2 = 4'd3; b_sign3 = 4'd3;
@(posedge clk_i);
a_mant0 = 8'd196; a_mant1 = 8'd59; a_mant2 = 8'd10; a_mant3 = 8'd126;
b_mant0 = 8'd222; b_mant1 = 8'd41; b_mant2 = 8'd107; b_mant3 = 8'd122;
a_exp0 = 10'd884; a_exp1 = 10'd537; a_exp2 = 10'd694; a_exp3 = 10'd640;
b_exp0 = 10'd551; b_exp1 = 10'd363; b_exp2 = 10'd859; b_exp3 = 10'd117;
a_sign0 = 4'd10; a_sign1 = 4'd7; a_sign2 = 4'd16; a_sign3 = 4'd16;
b_sign0 = 4'd13; b_sign1 = 4'd5; b_sign2 = 4'd11; b_sign3 = 4'd11;
@(posedge clk_i);
a_mant0 = 8'd216; a_mant1 = 8'd90; a_mant2 = 8'd45; a_mant3 = 8'd235;
b_mant0 = 8'd103; b_mant1 = 8'd221; b_mant2 = 8'd7; b_mant3 = 8'd73;
a_exp0 = 10'd630; a_exp1 = 10'd621; a_exp2 = 10'd914; a_exp3 = 10'd452;
b_exp0 = 10'd598; b_exp1 = 10'd541; b_exp2 = 10'd52; b_exp3 = 10'd787;
a_sign0 = 4'd0; a_sign1 = 4'd9; a_sign2 = 4'd11; a_sign3 = 4'd9;
b_sign0 = 4'd13; b_sign1 = 4'd5; b_sign2 = 4'd5; b_sign3 = 4'd2;
@(posedge clk_i);
shared_exps0 = 8'd152;
shared_exps1 = 8'd141;
rstn = 0;
@(posedge clk_i);
rstn = 1;
a_mant0 = 8'd254; a_mant1 = 8'd8; a_mant2 = 8'd203; a_mant3 = 8'd139;
b_mant0 = 8'd83; b_mant1 = 8'd238; b_mant2 = 8'd80; b_mant3 = 8'd52;
a_exp0 = 10'd740; a_exp1 = 10'd781; a_exp2 = 10'd468; a_exp3 = 10'd186;
b_exp0 = 10'd927; b_exp1 = 10'd512; b_exp2 = 10'd147; b_exp3 = 10'd400;
a_sign0 = 4'd10; a_sign1 = 4'd14; a_sign2 = 4'd14; a_sign3 = 4'd1;
b_sign0 = 4'd6; b_sign1 = 4'd10; b_sign2 = 4'd10; b_sign3 = 4'd3;
@(posedge clk_i);
a_mant0 = 8'd36; a_mant1 = 8'd14; a_mant2 = 8'd52; a_mant3 = 8'd170;
b_mant0 = 8'd143; b_mant1 = 8'd34; b_mant2 = 8'd182; b_mant3 = 8'd56;
a_exp0 = 10'd67; a_exp1 = 10'd70; a_exp2 = 10'd203; a_exp3 = 10'd251;
b_exp0 = 10'd182; b_exp1 = 10'd244; b_exp2 = 10'd135; b_exp3 = 10'd580;
a_sign0 = 4'd11; a_sign1 = 4'd4; a_sign2 = 4'd0; a_sign3 = 4'd16;
b_sign0 = 4'd9; b_sign1 = 4'd10; b_sign2 = 4'd9; b_sign3 = 4'd14;
@(posedge clk_i);
a_mant0 = 8'd194; a_mant1 = 8'd199; a_mant2 = 8'd239; a_mant3 = 8'd108;
b_mant0 = 8'd196; b_mant1 = 8'd181; b_mant2 = 8'd121; b_mant3 = 8'd238;
a_exp0 = 10'd558; a_exp1 = 10'd106; a_exp2 = 10'd646; a_exp3 = 10'd972;
b_exp0 = 10'd748; b_exp1 = 10'd332; b_exp2 = 10'd881; b_exp3 = 10'd76;
a_sign0 = 4'd8; a_sign1 = 4'd3; a_sign2 = 4'd11; a_sign3 = 4'd10;
b_sign0 = 4'd14; b_sign1 = 4'd16; b_sign2 = 4'd12; b_sign3 = 4'd0;
@(posedge clk_i);
a_mant0 = 8'd220; a_mant1 = 8'd164; a_mant2 = 8'd181; a_mant3 = 8'd40;
b_mant0 = 8'd122; b_mant1 = 8'd61; b_mant2 = 8'd191; b_mant3 = 8'd196;
a_exp0 = 10'd363; a_exp1 = 10'd190; a_exp2 = 10'd629; a_exp3 = 10'd978;
b_exp0 = 10'd260; b_exp1 = 10'd269; b_exp2 = 10'd125; b_exp3 = 10'd874;
a_sign0 = 4'd5; a_sign1 = 4'd9; a_sign2 = 4'd0; a_sign3 = 4'd5;
b_sign0 = 4'd5; b_sign1 = 4'd14; b_sign2 = 4'd13; b_sign3 = 4'd4;
@(posedge clk_i);
a_mant0 = 8'd189; a_mant1 = 8'd86; a_mant2 = 8'd33; a_mant3 = 8'd67;
b_mant0 = 8'd215; b_mant1 = 8'd235; b_mant2 = 8'd48; b_mant3 = 8'd31;
a_exp0 = 10'd382; a_exp1 = 10'd265; a_exp2 = 10'd610; a_exp3 = 10'd203;
b_exp0 = 10'd15; b_exp1 = 10'd796; b_exp2 = 10'd724; b_exp3 = 10'd984;
a_sign0 = 4'd10; a_sign1 = 4'd16; a_sign2 = 4'd11; a_sign3 = 4'd13;
b_sign0 = 4'd9; b_sign1 = 4'd13; b_sign2 = 4'd0; b_sign3 = 4'd9;
@(posedge clk_i);
a_mant0 = 8'd127; a_mant1 = 8'd186; a_mant2 = 8'd97; a_mant3 = 8'd112;
b_mant0 = 8'd155; b_mant1 = 8'd165; b_mant2 = 8'd22; b_mant3 = 8'd147;
a_exp0 = 10'd549; a_exp1 = 10'd1018; a_exp2 = 10'd477; a_exp3 = 10'd496;
b_exp0 = 10'd513; b_exp1 = 10'd252; b_exp2 = 10'd90; b_exp3 = 10'd192;
a_sign0 = 4'd13; a_sign1 = 4'd6; a_sign2 = 4'd2; a_sign3 = 4'd3;
b_sign0 = 4'd14; b_sign1 = 4'd14; b_sign2 = 4'd14; b_sign3 = 4'd1;
@(posedge clk_i);
a_mant0 = 8'd39; a_mant1 = 8'd135; a_mant2 = 8'd220; a_mant3 = 8'd147;
b_mant0 = 8'd205; b_mant1 = 8'd254; b_mant2 = 8'd164; b_mant3 = 8'd219;
a_exp0 = 10'd137; a_exp1 = 10'd626; a_exp2 = 10'd303; a_exp3 = 10'd764;
b_exp0 = 10'd791; b_exp1 = 10'd33; b_exp2 = 10'd371; b_exp3 = 10'd484;
a_sign0 = 4'd14; a_sign1 = 4'd13; a_sign2 = 4'd5; a_sign3 = 4'd16;
b_sign0 = 4'd4; b_sign1 = 4'd13; b_sign2 = 4'd8; b_sign3 = 4'd14;
@(posedge clk_i);
shared_exps0 = 8'd125;
shared_exps1 = 8'd147;
a_mant0 = 8'd109; a_mant1 = 8'd234; a_mant2 = 8'd236; a_mant3 = 8'd49;
b_mant0 = 8'd201; b_mant1 = 8'd160; b_mant2 = 8'd108; b_mant3 = 8'd202;
a_exp0 = 10'd90; a_exp1 = 10'd707; a_exp2 = 10'd929; a_exp3 = 10'd419;
b_exp0 = 10'd82; b_exp1 = 10'd959; b_exp2 = 10'd906; b_exp3 = 10'd309;
a_sign0 = 4'd6; a_sign1 = 4'd9; a_sign2 = 4'd5; a_sign3 = 4'd14;
b_sign0 = 4'd3; b_sign1 = 4'd8; b_sign2 = 4'd14; b_sign3 = 4'd14;
@(posedge clk_i);
a_mant0 = 8'd233; a_mant1 = 8'd48; a_mant2 = 8'd135; a_mant3 = 8'd230;
b_mant0 = 8'd115; b_mant1 = 8'd153; b_mant2 = 8'd179; b_mant3 = 8'd191;
a_exp0 = 10'd419; a_exp1 = 10'd46; a_exp2 = 10'd48; a_exp3 = 10'd740;
b_exp0 = 10'd349; b_exp1 = 10'd162; b_exp2 = 10'd996; b_exp3 = 10'd282;
a_sign0 = 4'd6; a_sign1 = 4'd5; a_sign2 = 4'd3; a_sign3 = 4'd8;
b_sign0 = 4'd9; b_sign1 = 4'd12; b_sign2 = 4'd5; b_sign3 = 4'd15;
@(posedge clk_i);
a_mant0 = 8'd119; a_mant1 = 8'd244; a_mant2 = 8'd120; a_mant3 = 8'd157;
b_mant0 = 8'd144; b_mant1 = 8'd129; b_mant2 = 8'd16; b_mant3 = 8'd29;
a_exp0 = 10'd995; a_exp1 = 10'd214; a_exp2 = 10'd163; a_exp3 = 10'd807;
b_exp0 = 10'd456; b_exp1 = 10'd469; b_exp2 = 10'd466; b_exp3 = 10'd999;
a_sign0 = 4'd7; a_sign1 = 4'd8; a_sign2 = 4'd8; a_sign3 = 4'd5;
b_sign0 = 4'd11; b_sign1 = 4'd8; b_sign2 = 4'd10; b_sign3 = 4'd1;
@(posedge clk_i);
a_mant0 = 8'd106; a_mant1 = 8'd227; a_mant2 = 8'd137; a_mant3 = 8'd218;
b_mant0 = 8'd121; b_mant1 = 8'd29; b_mant2 = 8'd216; b_mant3 = 8'd190;
a_exp0 = 10'd713; a_exp1 = 10'd299; a_exp2 = 10'd147; a_exp3 = 10'd805;
b_exp0 = 10'd266; b_exp1 = 10'd669; b_exp2 = 10'd999; b_exp3 = 10'd102;
a_sign0 = 4'd6; a_sign1 = 4'd0; a_sign2 = 4'd11; a_sign3 = 4'd4;
b_sign0 = 4'd7; b_sign1 = 4'd8; b_sign2 = 4'd16; b_sign3 = 4'd10;
@(posedge clk_i);
a_mant0 = 8'd68; a_mant1 = 8'd91; a_mant2 = 8'd175; a_mant3 = 8'd160;
b_mant0 = 8'd178; b_mant1 = 8'd21; b_mant2 = 8'd152; b_mant3 = 8'd59;
a_exp0 = 10'd38; a_exp1 = 10'd188; a_exp2 = 10'd517; a_exp3 = 10'd363;
b_exp0 = 10'd237; b_exp1 = 10'd144; b_exp2 = 10'd991; b_exp3 = 10'd192;
a_sign0 = 4'd16; a_sign1 = 4'd3; a_sign2 = 4'd12; a_sign3 = 4'd11;
b_sign0 = 4'd9; b_sign1 = 4'd8; b_sign2 = 4'd7; b_sign3 = 4'd16;
@(posedge clk_i);
a_mant0 = 8'd74; a_mant1 = 8'd220; a_mant2 = 8'd202; a_mant3 = 8'd99;
b_mant0 = 8'd139; b_mant1 = 8'd113; b_mant2 = 8'd125; b_mant3 = 8'd117;
a_exp0 = 10'd48; a_exp1 = 10'd613; a_exp2 = 10'd292; a_exp3 = 10'd797;
b_exp0 = 10'd625; b_exp1 = 10'd59; b_exp2 = 10'd142; b_exp3 = 10'd981;
a_sign0 = 4'd12; a_sign1 = 4'd4; a_sign2 = 4'd12; a_sign3 = 4'd12;
b_sign0 = 4'd1; b_sign1 = 4'd14; b_sign2 = 4'd11; b_sign3 = 4'd2;
@(posedge clk_i);
a_mant0 = 8'd242; a_mant1 = 8'd157; a_mant2 = 8'd121; a_mant3 = 8'd148;
b_mant0 = 8'd24; b_mant1 = 8'd45; b_mant2 = 8'd183; b_mant3 = 8'd105;
a_exp0 = 10'd529; a_exp1 = 10'd152; a_exp2 = 10'd564; a_exp3 = 10'd312;
b_exp0 = 10'd317; b_exp1 = 10'd844; b_exp2 = 10'd456; b_exp3 = 10'd739;
a_sign0 = 4'd2; a_sign1 = 4'd15; a_sign2 = 4'd0; a_sign3 = 4'd3;
b_sign0 = 4'd7; b_sign1 = 4'd7; b_sign2 = 4'd3; b_sign3 = 4'd13;
@(posedge clk_i);
a_mant0 = 8'd169; a_mant1 = 8'd244; a_mant2 = 8'd130; a_mant3 = 8'd44;
b_mant0 = 8'd228; b_mant1 = 8'd65; b_mant2 = 8'd115; b_mant3 = 8'd44;
a_exp0 = 10'd103; a_exp1 = 10'd754; a_exp2 = 10'd212; a_exp3 = 10'd716;
b_exp0 = 10'd523; b_exp1 = 10'd597; b_exp2 = 10'd994; b_exp3 = 10'd888;
a_sign0 = 4'd15; a_sign1 = 4'd2; a_sign2 = 4'd8; a_sign3 = 4'd13;
b_sign0 = 4'd9; b_sign1 = 4'd13; b_sign2 = 4'd6; b_sign3 = 4'd0;
@(posedge clk_i);
shared_exps0 = 8'd133;
shared_exps1 = 8'd123;
a_mant0 = 8'd59; a_mant1 = 8'd96; a_mant2 = 8'd82; a_mant3 = 8'd192;
b_mant0 = 8'd97; b_mant1 = 8'd182; b_mant2 = 8'd226; b_mant3 = 8'd89;
a_exp0 = 10'd27; a_exp1 = 10'd28; a_exp2 = 10'd1008; a_exp3 = 10'd161;
b_exp0 = 10'd210; b_exp1 = 10'd398; b_exp2 = 10'd800; b_exp3 = 10'd816;
a_sign0 = 4'd6; a_sign1 = 4'd16; a_sign2 = 4'd0; a_sign3 = 4'd2;
b_sign0 = 4'd16; b_sign1 = 4'd14; b_sign2 = 4'd3; b_sign3 = 4'd5;
@(posedge clk_i);
a_mant0 = 8'd196; a_mant1 = 8'd1; a_mant2 = 8'd207; a_mant3 = 8'd87;
b_mant0 = 8'd198; b_mant1 = 8'd159; b_mant2 = 8'd31; b_mant3 = 8'd80;
a_exp0 = 10'd1012; a_exp1 = 10'd469; a_exp2 = 10'd942; a_exp3 = 10'd886;
b_exp0 = 10'd908; b_exp1 = 10'd804; b_exp2 = 10'd896; b_exp3 = 10'd916;
a_sign0 = 4'd1; a_sign1 = 4'd4; a_sign2 = 4'd14; a_sign3 = 4'd12;
b_sign0 = 4'd12; b_sign1 = 4'd8; b_sign2 = 4'd8; b_sign3 = 4'd8;
@(posedge clk_i);
a_mant0 = 8'd165; a_mant1 = 8'd14; a_mant2 = 8'd119; a_mant3 = 8'd106;
b_mant0 = 8'd15; b_mant1 = 8'd143; b_mant2 = 8'd141; b_mant3 = 8'd39;
a_exp0 = 10'd881; a_exp1 = 10'd124; a_exp2 = 10'd205; a_exp3 = 10'd221;
b_exp0 = 10'd790; b_exp1 = 10'd702; b_exp2 = 10'd256; b_exp3 = 10'd719;
a_sign0 = 4'd4; a_sign1 = 4'd0; a_sign2 = 4'd0; a_sign3 = 4'd10;
b_sign0 = 4'd5; b_sign1 = 4'd9; b_sign2 = 4'd12; b_sign3 = 4'd10;
@(posedge clk_i);
a_mant0 = 8'd62; a_mant1 = 8'd172; a_mant2 = 8'd33; a_mant3 = 8'd218;
b_mant0 = 8'd18; b_mant1 = 8'd67; b_mant2 = 8'd159; b_mant3 = 8'd118;
a_exp0 = 10'd581; a_exp1 = 10'd100; a_exp2 = 10'd333; a_exp3 = 10'd86;
b_exp0 = 10'd79; b_exp1 = 10'd276; b_exp2 = 10'd818; b_exp3 = 10'd785;
a_sign0 = 4'd1; a_sign1 = 4'd14; a_sign2 = 4'd7; a_sign3 = 4'd5;
b_sign0 = 4'd13; b_sign1 = 4'd3; b_sign2 = 4'd4; b_sign3 = 4'd8;
@(posedge clk_i);
a_mant0 = 8'd103; a_mant1 = 8'd148; a_mant2 = 8'd94; a_mant3 = 8'd168;
b_mant0 = 8'd245; b_mant1 = 8'd128; b_mant2 = 8'd174; b_mant3 = 8'd235;
a_exp0 = 10'd522; a_exp1 = 10'd837; a_exp2 = 10'd949; a_exp3 = 10'd391;
b_exp0 = 10'd270; b_exp1 = 10'd34; b_exp2 = 10'd788; b_exp3 = 10'd948;
a_sign0 = 4'd14; a_sign1 = 4'd4; a_sign2 = 4'd16; a_sign3 = 4'd8;
b_sign0 = 4'd9; b_sign1 = 4'd14; b_sign2 = 4'd16; b_sign3 = 4'd0;
@(posedge clk_i);
a_mant0 = 8'd42; a_mant1 = 8'd95; a_mant2 = 8'd2; a_mant3 = 8'd169;
b_mant0 = 8'd16; b_mant1 = 8'd76; b_mant2 = 8'd19; b_mant3 = 8'd86;
a_exp0 = 10'd374; a_exp1 = 10'd140; a_exp2 = 10'd521; a_exp3 = 10'd390;
b_exp0 = 10'd814; b_exp1 = 10'd310; b_exp2 = 10'd144; b_exp3 = 10'd999;
a_sign0 = 4'd4; a_sign1 = 4'd7; a_sign2 = 4'd14; a_sign3 = 4'd6;
b_sign0 = 4'd9; b_sign1 = 4'd16; b_sign2 = 4'd10; b_sign3 = 4'd6;
@(posedge clk_i);
a_mant0 = 8'd19; a_mant1 = 8'd64; a_mant2 = 8'd178; a_mant3 = 8'd122;
b_mant0 = 8'd69; b_mant1 = 8'd129; b_mant2 = 8'd75; b_mant3 = 8'd18;
a_exp0 = 10'd245; a_exp1 = 10'd861; a_exp2 = 10'd205; a_exp3 = 10'd406;
b_exp0 = 10'd384; b_exp1 = 10'd772; b_exp2 = 10'd131; b_exp3 = 10'd3;
a_sign0 = 4'd16; a_sign1 = 4'd7; a_sign2 = 4'd4; a_sign3 = 4'd5;
b_sign0 = 4'd6; b_sign1 = 4'd16; b_sign2 = 4'd11; b_sign3 = 4'd14;
@(posedge clk_i);
a_mant0 = 8'd104; a_mant1 = 8'd46; a_mant2 = 8'd112; a_mant3 = 8'd145;
b_mant0 = 8'd238; b_mant1 = 8'd169; b_mant2 = 8'd130; b_mant3 = 8'd20;
a_exp0 = 10'd899; a_exp1 = 10'd307; a_exp2 = 10'd655; a_exp3 = 10'd432;
b_exp0 = 10'd321; b_exp1 = 10'd287; b_exp2 = 10'd636; b_exp3 = 10'd675;
a_sign0 = 4'd6; a_sign1 = 4'd2; a_sign2 = 4'd3; a_sign3 = 4'd8;
b_sign0 = 4'd11; b_sign1 = 4'd15; b_sign2 = 4'd4; b_sign3 = 4'd4;
@(posedge clk_i);
shared_exps0 = 8'd104;
shared_exps1 = 8'd143;
a_mant0 = 8'd113; a_mant1 = 8'd120; a_mant2 = 8'd69; a_mant3 = 8'd54;
b_mant0 = 8'd131; b_mant1 = 8'd38; b_mant2 = 8'd190; b_mant3 = 8'd12;
a_exp0 = 10'd528; a_exp1 = 10'd863; a_exp2 = 10'd649; a_exp3 = 10'd472;
b_exp0 = 10'd741; b_exp1 = 10'd1021; b_exp2 = 10'd852; b_exp3 = 10'd0;
a_sign0 = 4'd4; a_sign1 = 4'd7; a_sign2 = 4'd15; a_sign3 = 4'd5;
b_sign0 = 4'd15; b_sign1 = 4'd11; b_sign2 = 4'd0; b_sign3 = 4'd16;
@(posedge clk_i);
a_mant0 = 8'd10; a_mant1 = 8'd202; a_mant2 = 8'd184; a_mant3 = 8'd104;
b_mant0 = 8'd203; b_mant1 = 8'd182; b_mant2 = 8'd90; b_mant3 = 8'd24;
a_exp0 = 10'd347; a_exp1 = 10'd523; a_exp2 = 10'd482; a_exp3 = 10'd324;
b_exp0 = 10'd710; b_exp1 = 10'd4; b_exp2 = 10'd58; b_exp3 = 10'd486;
a_sign0 = 4'd12; a_sign1 = 4'd8; a_sign2 = 4'd9; a_sign3 = 4'd2;
b_sign0 = 4'd15; b_sign1 = 4'd3; b_sign2 = 4'd10; b_sign3 = 4'd16;
@(posedge clk_i);
a_mant0 = 8'd236; a_mant1 = 8'd13; a_mant2 = 8'd85; a_mant3 = 8'd93;
b_mant0 = 8'd230; b_mant1 = 8'd35; b_mant2 = 8'd248; b_mant3 = 8'd92;
a_exp0 = 10'd977; a_exp1 = 10'd325; a_exp2 = 10'd899; a_exp3 = 10'd118;
b_exp0 = 10'd589; b_exp1 = 10'd498; b_exp2 = 10'd128; b_exp3 = 10'd542;
a_sign0 = 4'd15; a_sign1 = 4'd7; a_sign2 = 4'd1; a_sign3 = 4'd4;
b_sign0 = 4'd9; b_sign1 = 4'd13; b_sign2 = 4'd14; b_sign3 = 4'd6;
@(posedge clk_i);
a_mant0 = 8'd90; a_mant1 = 8'd29; a_mant2 = 8'd97; a_mant3 = 8'd34;
b_mant0 = 8'd74; b_mant1 = 8'd168; b_mant2 = 8'd13; b_mant3 = 8'd153;
a_exp0 = 10'd993; a_exp1 = 10'd706; a_exp2 = 10'd703; a_exp3 = 10'd611;
b_exp0 = 10'd312; b_exp1 = 10'd572; b_exp2 = 10'd68; b_exp3 = 10'd97;
a_sign0 = 4'd3; a_sign1 = 4'd2; a_sign2 = 4'd1; a_sign3 = 4'd10;
b_sign0 = 4'd16; b_sign1 = 4'd15; b_sign2 = 4'd10; b_sign3 = 4'd4;
@(posedge clk_i);
a_mant0 = 8'd31; a_mant1 = 8'd44; a_mant2 = 8'd116; a_mant3 = 8'd205;
b_mant0 = 8'd80; b_mant1 = 8'd86; b_mant2 = 8'd87; b_mant3 = 8'd147;
a_exp0 = 10'd566; a_exp1 = 10'd741; a_exp2 = 10'd148; a_exp3 = 10'd219;
b_exp0 = 10'd960; b_exp1 = 10'd639; b_exp2 = 10'd781; b_exp3 = 10'd1010;
a_sign0 = 4'd10; a_sign1 = 4'd9; a_sign2 = 4'd8; a_sign3 = 4'd1;
b_sign0 = 4'd4; b_sign1 = 4'd8; b_sign2 = 4'd11; b_sign3 = 4'd9;
@(posedge clk_i);
a_mant0 = 8'd16; a_mant1 = 8'd95; a_mant2 = 8'd101; a_mant3 = 8'd107;
b_mant0 = 8'd108; b_mant1 = 8'd99; b_mant2 = 8'd180; b_mant3 = 8'd127;
a_exp0 = 10'd724; a_exp1 = 10'd493; a_exp2 = 10'd67; a_exp3 = 10'd943;
b_exp0 = 10'd757; b_exp1 = 10'd651; b_exp2 = 10'd247; b_exp3 = 10'd47;
a_sign0 = 4'd3; a_sign1 = 4'd12; a_sign2 = 4'd9; a_sign3 = 4'd14;
b_sign0 = 4'd2; b_sign1 = 4'd9; b_sign2 = 4'd4; b_sign3 = 4'd3;
@(posedge clk_i);
a_mant0 = 8'd18; a_mant1 = 8'd17; a_mant2 = 8'd32; a_mant3 = 8'd227;
b_mant0 = 8'd254; b_mant1 = 8'd240; b_mant2 = 8'd88; b_mant3 = 8'd166;
a_exp0 = 10'd738; a_exp1 = 10'd291; a_exp2 = 10'd105; a_exp3 = 10'd71;
b_exp0 = 10'd28; b_exp1 = 10'd970; b_exp2 = 10'd61; b_exp3 = 10'd69;
a_sign0 = 4'd0; a_sign1 = 4'd2; a_sign2 = 4'd9; a_sign3 = 4'd2;
b_sign0 = 4'd0; b_sign1 = 4'd15; b_sign2 = 4'd11; b_sign3 = 4'd13;
@(posedge clk_i);
a_mant0 = 8'd56; a_mant1 = 8'd236; a_mant2 = 8'd75; a_mant3 = 8'd89;
b_mant0 = 8'd220; b_mant1 = 8'd173; b_mant2 = 8'd118; b_mant3 = 8'd252;
a_exp0 = 10'd936; a_exp1 = 10'd907; a_exp2 = 10'd362; a_exp3 = 10'd0;
b_exp0 = 10'd344; b_exp1 = 10'd736; b_exp2 = 10'd691; b_exp3 = 10'd843;
a_sign0 = 4'd0; a_sign1 = 4'd10; a_sign2 = 4'd9; a_sign3 = 4'd0;
b_sign0 = 4'd5; b_sign1 = 4'd10; b_sign2 = 4'd13; b_sign3 = 4'd6;
@(posedge clk_i);
shared_exps0 = 8'd114;
shared_exps1 = 8'd134;
rstn = 0;
@(posedge clk_i);
rstn = 1;
a_mant0 = 8'd173; a_mant1 = 8'd103; a_mant2 = 8'd65; a_mant3 = 8'd252;
b_mant0 = 8'd51; b_mant1 = 8'd191; b_mant2 = 8'd253; b_mant3 = 8'd123;
a_exp0 = 10'd264; a_exp1 = 10'd452; a_exp2 = 10'd245; a_exp3 = 10'd954;
b_exp0 = 10'd880; b_exp1 = 10'd241; b_exp2 = 10'd343; b_exp3 = 10'd640;
a_sign0 = 4'd1; a_sign1 = 4'd5; a_sign2 = 4'd6; a_sign3 = 4'd4;
b_sign0 = 4'd2; b_sign1 = 4'd7; b_sign2 = 4'd4; b_sign3 = 4'd15;
@(posedge clk_i);
a_mant0 = 8'd71; a_mant1 = 8'd23; a_mant2 = 8'd38; a_mant3 = 8'd61;
b_mant0 = 8'd199; b_mant1 = 8'd84; b_mant2 = 8'd198; b_mant3 = 8'd138;
a_exp0 = 10'd846; a_exp1 = 10'd538; a_exp2 = 10'd81; a_exp3 = 10'd717;
b_exp0 = 10'd937; b_exp1 = 10'd710; b_exp2 = 10'd253; b_exp3 = 10'd912;
a_sign0 = 4'd2; a_sign1 = 4'd16; a_sign2 = 4'd12; a_sign3 = 4'd6;
b_sign0 = 4'd9; b_sign1 = 4'd6; b_sign2 = 4'd4; b_sign3 = 4'd12;
@(posedge clk_i);
a_mant0 = 8'd184; a_mant1 = 8'd117; a_mant2 = 8'd168; a_mant3 = 8'd189;
b_mant0 = 8'd74; b_mant1 = 8'd127; b_mant2 = 8'd80; b_mant3 = 8'd38;
a_exp0 = 10'd888; a_exp1 = 10'd839; a_exp2 = 10'd30; a_exp3 = 10'd263;
b_exp0 = 10'd752; b_exp1 = 10'd63; b_exp2 = 10'd449; b_exp3 = 10'd879;
a_sign0 = 4'd2; a_sign1 = 4'd7; a_sign2 = 4'd16; a_sign3 = 4'd15;
b_sign0 = 4'd12; b_sign1 = 4'd12; b_sign2 = 4'd3; b_sign3 = 4'd1;
@(posedge clk_i);
a_mant0 = 8'd121; a_mant1 = 8'd18; a_mant2 = 8'd57; a_mant3 = 8'd234;
b_mant0 = 8'd182; b_mant1 = 8'd117; b_mant2 = 8'd196; b_mant3 = 8'd132;
a_exp0 = 10'd973; a_exp1 = 10'd597; a_exp2 = 10'd457; a_exp3 = 10'd470;
b_exp0 = 10'd573; b_exp1 = 10'd325; b_exp2 = 10'd919; b_exp3 = 10'd169;
a_sign0 = 4'd2; a_sign1 = 4'd13; a_sign2 = 4'd1; a_sign3 = 4'd1;
b_sign0 = 4'd14; b_sign1 = 4'd10; b_sign2 = 4'd5; b_sign3 = 4'd9;
@(posedge clk_i);
a_mant0 = 8'd240; a_mant1 = 8'd118; a_mant2 = 8'd214; a_mant3 = 8'd98;
b_mant0 = 8'd16; b_mant1 = 8'd188; b_mant2 = 8'd244; b_mant3 = 8'd210;
a_exp0 = 10'd112; a_exp1 = 10'd206; a_exp2 = 10'd503; a_exp3 = 10'd855;
b_exp0 = 10'd569; b_exp1 = 10'd225; b_exp2 = 10'd885; b_exp3 = 10'd953;
a_sign0 = 4'd1; a_sign1 = 4'd8; a_sign2 = 4'd12; a_sign3 = 4'd0;
b_sign0 = 4'd2; b_sign1 = 4'd16; b_sign2 = 4'd1; b_sign3 = 4'd12;
@(posedge clk_i);
a_mant0 = 8'd254; a_mant1 = 8'd66; a_mant2 = 8'd196; a_mant3 = 8'd152;
b_mant0 = 8'd187; b_mant1 = 8'd80; b_mant2 = 8'd74; b_mant3 = 8'd233;
a_exp0 = 10'd696; a_exp1 = 10'd648; a_exp2 = 10'd928; a_exp3 = 10'd669;
b_exp0 = 10'd397; b_exp1 = 10'd870; b_exp2 = 10'd922; b_exp3 = 10'd23;
a_sign0 = 4'd1; a_sign1 = 4'd7; a_sign2 = 4'd15; a_sign3 = 4'd15;
b_sign0 = 4'd5; b_sign1 = 4'd3; b_sign2 = 4'd8; b_sign3 = 4'd6;
@(posedge clk_i);
a_mant0 = 8'd143; a_mant1 = 8'd147; a_mant2 = 8'd170; a_mant3 = 8'd238;
b_mant0 = 8'd169; b_mant1 = 8'd106; b_mant2 = 8'd116; b_mant3 = 8'd65;
a_exp0 = 10'd750; a_exp1 = 10'd816; a_exp2 = 10'd295; a_exp3 = 10'd611;
b_exp0 = 10'd41; b_exp1 = 10'd113; b_exp2 = 10'd122; b_exp3 = 10'd989;
a_sign0 = 4'd11; a_sign1 = 4'd4; a_sign2 = 4'd15; a_sign3 = 4'd4;
b_sign0 = 4'd3; b_sign1 = 4'd0; b_sign2 = 4'd0; b_sign3 = 4'd8;
@(posedge clk_i);
shared_exps0 = 8'd146;
shared_exps1 = 8'd137;
a_mant0 = 8'd181; a_mant1 = 8'd54; a_mant2 = 8'd90; a_mant3 = 8'd166;
b_mant0 = 8'd158; b_mant1 = 8'd64; b_mant2 = 8'd244; b_mant3 = 8'd199;
a_exp0 = 10'd243; a_exp1 = 10'd863; a_exp2 = 10'd35; a_exp3 = 10'd899;
b_exp0 = 10'd573; b_exp1 = 10'd601; b_exp2 = 10'd317; b_exp3 = 10'd995;
a_sign0 = 4'd11; a_sign1 = 4'd3; a_sign2 = 4'd9; a_sign3 = 4'd14;
b_sign0 = 4'd10; b_sign1 = 4'd10; b_sign2 = 4'd6; b_sign3 = 4'd2;
@(posedge clk_i);
a_mant0 = 8'd236; a_mant1 = 8'd208; a_mant2 = 8'd60; a_mant3 = 8'd122;
b_mant0 = 8'd182; b_mant1 = 8'd90; b_mant2 = 8'd81; b_mant3 = 8'd69;
a_exp0 = 10'd797; a_exp1 = 10'd108; a_exp2 = 10'd159; a_exp3 = 10'd379;
b_exp0 = 10'd705; b_exp1 = 10'd175; b_exp2 = 10'd929; b_exp3 = 10'd580;
a_sign0 = 4'd11; a_sign1 = 4'd10; a_sign2 = 4'd14; a_sign3 = 4'd4;
b_sign0 = 4'd15; b_sign1 = 4'd11; b_sign2 = 4'd9; b_sign3 = 4'd11;
@(posedge clk_i);
a_mant0 = 8'd88; a_mant1 = 8'd232; a_mant2 = 8'd251; a_mant3 = 8'd195;
b_mant0 = 8'd247; b_mant1 = 8'd31; b_mant2 = 8'd240; b_mant3 = 8'd60;
a_exp0 = 10'd686; a_exp1 = 10'd240; a_exp2 = 10'd304; a_exp3 = 10'd801;
b_exp0 = 10'd853; b_exp1 = 10'd294; b_exp2 = 10'd437; b_exp3 = 10'd1;
a_sign0 = 4'd14; a_sign1 = 4'd1; a_sign2 = 4'd9; a_sign3 = 4'd6;
b_sign0 = 4'd0; b_sign1 = 4'd11; b_sign2 = 4'd1; b_sign3 = 4'd4;
@(posedge clk_i);
a_mant0 = 8'd115; a_mant1 = 8'd56; a_mant2 = 8'd122; a_mant3 = 8'd15;
b_mant0 = 8'd211; b_mant1 = 8'd154; b_mant2 = 8'd80; b_mant3 = 8'd11;
a_exp0 = 10'd149; a_exp1 = 10'd801; a_exp2 = 10'd766; a_exp3 = 10'd438;
b_exp0 = 10'd446; b_exp1 = 10'd749; b_exp2 = 10'd746; b_exp3 = 10'd680;
a_sign0 = 4'd14; a_sign1 = 4'd8; a_sign2 = 4'd4; a_sign3 = 4'd2;
b_sign0 = 4'd8; b_sign1 = 4'd5; b_sign2 = 4'd5; b_sign3 = 4'd14;
@(posedge clk_i);
a_mant0 = 8'd228; a_mant1 = 8'd27; a_mant2 = 8'd73; a_mant3 = 8'd15;
b_mant0 = 8'd151; b_mant1 = 8'd110; b_mant2 = 8'd147; b_mant3 = 8'd173;
a_exp0 = 10'd24; a_exp1 = 10'd192; a_exp2 = 10'd941; a_exp3 = 10'd830;
b_exp0 = 10'd588; b_exp1 = 10'd300; b_exp2 = 10'd592; b_exp3 = 10'd509;
a_sign0 = 4'd10; a_sign1 = 4'd15; a_sign2 = 4'd7; a_sign3 = 4'd13;
b_sign0 = 4'd16; b_sign1 = 4'd12; b_sign2 = 4'd7; b_sign3 = 4'd12;
@(posedge clk_i);
a_mant0 = 8'd35; a_mant1 = 8'd185; a_mant2 = 8'd111; a_mant3 = 8'd104;
b_mant0 = 8'd176; b_mant1 = 8'd36; b_mant2 = 8'd167; b_mant3 = 8'd162;
a_exp0 = 10'd334; a_exp1 = 10'd26; a_exp2 = 10'd167; a_exp3 = 10'd194;
b_exp0 = 10'd90; b_exp1 = 10'd444; b_exp2 = 10'd636; b_exp3 = 10'd409;
a_sign0 = 4'd15; a_sign1 = 4'd8; a_sign2 = 4'd11; a_sign3 = 4'd0;
b_sign0 = 4'd9; b_sign1 = 4'd12; b_sign2 = 4'd16; b_sign3 = 4'd12;
@(posedge clk_i);
a_mant0 = 8'd43; a_mant1 = 8'd224; a_mant2 = 8'd64; a_mant3 = 8'd143;
b_mant0 = 8'd38; b_mant1 = 8'd75; b_mant2 = 8'd21; b_mant3 = 8'd15;
a_exp0 = 10'd608; a_exp1 = 10'd591; a_exp2 = 10'd254; a_exp3 = 10'd634;
b_exp0 = 10'd413; b_exp1 = 10'd427; b_exp2 = 10'd357; b_exp3 = 10'd577;
a_sign0 = 4'd11; a_sign1 = 4'd3; a_sign2 = 4'd7; a_sign3 = 4'd10;
b_sign0 = 4'd14; b_sign1 = 4'd2; b_sign2 = 4'd0; b_sign3 = 4'd13;
@(posedge clk_i);
a_mant0 = 8'd235; a_mant1 = 8'd0; a_mant2 = 8'd198; a_mant3 = 8'd241;
b_mant0 = 8'd59; b_mant1 = 8'd75; b_mant2 = 8'd38; b_mant3 = 8'd120;
a_exp0 = 10'd351; a_exp1 = 10'd659; a_exp2 = 10'd206; a_exp3 = 10'd58;
b_exp0 = 10'd152; b_exp1 = 10'd991; b_exp2 = 10'd21; b_exp3 = 10'd425;
a_sign0 = 4'd4; a_sign1 = 4'd4; a_sign2 = 4'd7; a_sign3 = 4'd11;
b_sign0 = 4'd7; b_sign1 = 4'd9; b_sign2 = 4'd4; b_sign3 = 4'd2;
@(posedge clk_i);
shared_exps0 = 8'd131;
shared_exps1 = 8'd133;
a_mant0 = 8'd176; a_mant1 = 8'd9; a_mant2 = 8'd174; a_mant3 = 8'd177;
b_mant0 = 8'd79; b_mant1 = 8'd148; b_mant2 = 8'd119; b_mant3 = 8'd156;
a_exp0 = 10'd437; a_exp1 = 10'd24; a_exp2 = 10'd829; a_exp3 = 10'd202;
b_exp0 = 10'd500; b_exp1 = 10'd107; b_exp2 = 10'd505; b_exp3 = 10'd610;
a_sign0 = 4'd10; a_sign1 = 4'd8; a_sign2 = 4'd2; a_sign3 = 4'd2;
b_sign0 = 4'd9; b_sign1 = 4'd16; b_sign2 = 4'd7; b_sign3 = 4'd15;
@(posedge clk_i);
a_mant0 = 8'd230; a_mant1 = 8'd146; a_mant2 = 8'd113; a_mant3 = 8'd203;
b_mant0 = 8'd22; b_mant1 = 8'd49; b_mant2 = 8'd240; b_mant3 = 8'd112;
a_exp0 = 10'd381; a_exp1 = 10'd866; a_exp2 = 10'd238; a_exp3 = 10'd655;
b_exp0 = 10'd966; b_exp1 = 10'd625; b_exp2 = 10'd4; b_exp3 = 10'd174;
a_sign0 = 4'd16; a_sign1 = 4'd7; a_sign2 = 4'd9; a_sign3 = 4'd5;
b_sign0 = 4'd13; b_sign1 = 4'd10; b_sign2 = 4'd9; b_sign3 = 4'd5;
@(posedge clk_i);
a_mant0 = 8'd168; a_mant1 = 8'd106; a_mant2 = 8'd6; a_mant3 = 8'd191;
b_mant0 = 8'd68; b_mant1 = 8'd146; b_mant2 = 8'd124; b_mant3 = 8'd225;
a_exp0 = 10'd880; a_exp1 = 10'd728; a_exp2 = 10'd591; a_exp3 = 10'd481;
b_exp0 = 10'd340; b_exp1 = 10'd63; b_exp2 = 10'd787; b_exp3 = 10'd701;
a_sign0 = 4'd10; a_sign1 = 4'd16; a_sign2 = 4'd2; a_sign3 = 4'd16;
b_sign0 = 4'd10; b_sign1 = 4'd5; b_sign2 = 4'd13; b_sign3 = 4'd5;
@(posedge clk_i);
a_mant0 = 8'd172; a_mant1 = 8'd192; a_mant2 = 8'd76; a_mant3 = 8'd65;
b_mant0 = 8'd215; b_mant1 = 8'd158; b_mant2 = 8'd150; b_mant3 = 8'd253;
a_exp0 = 10'd662; a_exp1 = 10'd841; a_exp2 = 10'd985; a_exp3 = 10'd374;
b_exp0 = 10'd692; b_exp1 = 10'd944; b_exp2 = 10'd941; b_exp3 = 10'd395;
a_sign0 = 4'd9; a_sign1 = 4'd13; a_sign2 = 4'd16; a_sign3 = 4'd6;
b_sign0 = 4'd11; b_sign1 = 4'd4; b_sign2 = 4'd3; b_sign3 = 4'd2;
@(posedge clk_i);
a_mant0 = 8'd112; a_mant1 = 8'd210; a_mant2 = 8'd110; a_mant3 = 8'd9;
b_mant0 = 8'd249; b_mant1 = 8'd205; b_mant2 = 8'd186; b_mant3 = 8'd21;
a_exp0 = 10'd502; a_exp1 = 10'd98; a_exp2 = 10'd345; a_exp3 = 10'd502;
b_exp0 = 10'd976; b_exp1 = 10'd639; b_exp2 = 10'd329; b_exp3 = 10'd555;
a_sign0 = 4'd5; a_sign1 = 4'd8; a_sign2 = 4'd12; a_sign3 = 4'd8;
b_sign0 = 4'd7; b_sign1 = 4'd12; b_sign2 = 4'd8; b_sign3 = 4'd16;
@(posedge clk_i);
a_mant0 = 8'd200; a_mant1 = 8'd70; a_mant2 = 8'd9; a_mant3 = 8'd53;
b_mant0 = 8'd212; b_mant1 = 8'd167; b_mant2 = 8'd68; b_mant3 = 8'd70;
a_exp0 = 10'd830; a_exp1 = 10'd896; a_exp2 = 10'd279; a_exp3 = 10'd958;
b_exp0 = 10'd336; b_exp1 = 10'd170; b_exp2 = 10'd432; b_exp3 = 10'd436;
a_sign0 = 4'd6; a_sign1 = 4'd8; a_sign2 = 4'd1; a_sign3 = 4'd16;
b_sign0 = 4'd7; b_sign1 = 4'd4; b_sign2 = 4'd2; b_sign3 = 4'd0;
@(posedge clk_i);
a_mant0 = 8'd249; a_mant1 = 8'd4; a_mant2 = 8'd196; a_mant3 = 8'd34;
b_mant0 = 8'd81; b_mant1 = 8'd90; b_mant2 = 8'd86; b_mant3 = 8'd164;
a_exp0 = 10'd470; a_exp1 = 10'd445; a_exp2 = 10'd283; a_exp3 = 10'd583;
b_exp0 = 10'd607; b_exp1 = 10'd205; b_exp2 = 10'd459; b_exp3 = 10'd624;
a_sign0 = 4'd8; a_sign1 = 4'd3; a_sign2 = 4'd12; a_sign3 = 4'd14;
b_sign0 = 4'd9; b_sign1 = 4'd3; b_sign2 = 4'd15; b_sign3 = 4'd10;
@(posedge clk_i);
a_mant0 = 8'd61; a_mant1 = 8'd116; a_mant2 = 8'd204; a_mant3 = 8'd164;
b_mant0 = 8'd4; b_mant1 = 8'd179; b_mant2 = 8'd193; b_mant3 = 8'd47;
a_exp0 = 10'd50; a_exp1 = 10'd777; a_exp2 = 10'd686; a_exp3 = 10'd746;
b_exp0 = 10'd431; b_exp1 = 10'd693; b_exp2 = 10'd582; b_exp3 = 10'd560;
a_sign0 = 4'd0; a_sign1 = 4'd6; a_sign2 = 4'd5; a_sign3 = 4'd7;
b_sign0 = 4'd3; b_sign1 = 4'd12; b_sign2 = 4'd14; b_sign3 = 4'd15;
@(posedge clk_i);
shared_exps0 = 8'd114;
shared_exps1 = 8'd112;
a_mant0 = 8'd85; a_mant1 = 8'd222; a_mant2 = 8'd241; a_mant3 = 8'd192;
b_mant0 = 8'd140; b_mant1 = 8'd163; b_mant2 = 8'd250; b_mant3 = 8'd104;
a_exp0 = 10'd763; a_exp1 = 10'd936; a_exp2 = 10'd370; a_exp3 = 10'd815;
b_exp0 = 10'd464; b_exp1 = 10'd945; b_exp2 = 10'd212; b_exp3 = 10'd131;
a_sign0 = 4'd6; a_sign1 = 4'd6; a_sign2 = 4'd0; a_sign3 = 4'd15;
b_sign0 = 4'd14; b_sign1 = 4'd8; b_sign2 = 4'd3; b_sign3 = 4'd14;
@(posedge clk_i);
a_mant0 = 8'd212; a_mant1 = 8'd60; a_mant2 = 8'd64; a_mant3 = 8'd250;
b_mant0 = 8'd152; b_mant1 = 8'd203; b_mant2 = 8'd26; b_mant3 = 8'd6;
a_exp0 = 10'd944; a_exp1 = 10'd578; a_exp2 = 10'd676; a_exp3 = 10'd576;
b_exp0 = 10'd207; b_exp1 = 10'd789; b_exp2 = 10'd10; b_exp3 = 10'd969;
a_sign0 = 4'd6; a_sign1 = 4'd2; a_sign2 = 4'd4; a_sign3 = 4'd2;
b_sign0 = 4'd3; b_sign1 = 4'd8; b_sign2 = 4'd15; b_sign3 = 4'd14;
@(posedge clk_i);
a_mant0 = 8'd94; a_mant1 = 8'd123; a_mant2 = 8'd2; a_mant3 = 8'd26;
b_mant0 = 8'd91; b_mant1 = 8'd137; b_mant2 = 8'd236; b_mant3 = 8'd120;
a_exp0 = 10'd243; a_exp1 = 10'd973; a_exp2 = 10'd606; a_exp3 = 10'd529;
b_exp0 = 10'd993; b_exp1 = 10'd235; b_exp2 = 10'd418; b_exp3 = 10'd288;
a_sign0 = 4'd3; a_sign1 = 4'd3; a_sign2 = 4'd16; a_sign3 = 4'd13;
b_sign0 = 4'd1; b_sign1 = 4'd1; b_sign2 = 4'd5; b_sign3 = 4'd0;
@(posedge clk_i);
a_mant0 = 8'd75; a_mant1 = 8'd233; a_mant2 = 8'd27; a_mant3 = 8'd41;
b_mant0 = 8'd83; b_mant1 = 8'd121; b_mant2 = 8'd153; b_mant3 = 8'd42;
a_exp0 = 10'd1004; a_exp1 = 10'd224; a_exp2 = 10'd878; a_exp3 = 10'd840;
b_exp0 = 10'd871; b_exp1 = 10'd203; b_exp2 = 10'd420; b_exp3 = 10'd17;
a_sign0 = 4'd11; a_sign1 = 4'd4; a_sign2 = 4'd4; a_sign3 = 4'd3;
b_sign0 = 4'd7; b_sign1 = 4'd5; b_sign2 = 4'd13; b_sign3 = 4'd8;
@(posedge clk_i);
a_mant0 = 8'd37; a_mant1 = 8'd233; a_mant2 = 8'd9; a_mant3 = 8'd49;
b_mant0 = 8'd166; b_mant1 = 8'd28; b_mant2 = 8'd216; b_mant3 = 8'd178;
a_exp0 = 10'd476; a_exp1 = 10'd96; a_exp2 = 10'd236; a_exp3 = 10'd341;
b_exp0 = 10'd42; b_exp1 = 10'd245; b_exp2 = 10'd189; b_exp3 = 10'd55;
a_sign0 = 4'd10; a_sign1 = 4'd14; a_sign2 = 4'd14; a_sign3 = 4'd3;
b_sign0 = 4'd15; b_sign1 = 4'd7; b_sign2 = 4'd1; b_sign3 = 4'd11;
@(posedge clk_i);
a_mant0 = 8'd199; a_mant1 = 8'd136; a_mant2 = 8'd131; a_mant3 = 8'd200;
b_mant0 = 8'd118; b_mant1 = 8'd29; b_mant2 = 8'd78; b_mant3 = 8'd72;
a_exp0 = 10'd785; a_exp1 = 10'd679; a_exp2 = 10'd831; a_exp3 = 10'd217;
b_exp0 = 10'd666; b_exp1 = 10'd30; b_exp2 = 10'd91; b_exp3 = 10'd905;
a_sign0 = 4'd13; a_sign1 = 4'd9; a_sign2 = 4'd4; a_sign3 = 4'd4;
b_sign0 = 4'd7; b_sign1 = 4'd8; b_sign2 = 4'd7; b_sign3 = 4'd9;
@(posedge clk_i);
a_mant0 = 8'd149; a_mant1 = 8'd95; a_mant2 = 8'd148; a_mant3 = 8'd112;
b_mant0 = 8'd242; b_mant1 = 8'd76; b_mant2 = 8'd41; b_mant3 = 8'd14;
a_exp0 = 10'd963; a_exp1 = 10'd718; a_exp2 = 10'd342; a_exp3 = 10'd329;
b_exp0 = 10'd627; b_exp1 = 10'd731; b_exp2 = 10'd28; b_exp3 = 10'd963;
a_sign0 = 4'd10; a_sign1 = 4'd13; a_sign2 = 4'd10; a_sign3 = 4'd12;
b_sign0 = 4'd9; b_sign1 = 4'd11; b_sign2 = 4'd10; b_sign3 = 4'd1;
@(posedge clk_i);
a_mant0 = 8'd109; a_mant1 = 8'd143; a_mant2 = 8'd141; a_mant3 = 8'd165;
b_mant0 = 8'd200; b_mant1 = 8'd195; b_mant2 = 8'd199; b_mant3 = 8'd148;
a_exp0 = 10'd270; a_exp1 = 10'd588; a_exp2 = 10'd687; a_exp3 = 10'd80;
b_exp0 = 10'd893; b_exp1 = 10'd799; b_exp2 = 10'd390; b_exp3 = 10'd919;
a_sign0 = 4'd10; a_sign1 = 4'd0; a_sign2 = 4'd1; a_sign3 = 4'd14;
b_sign0 = 4'd5; b_sign1 = 4'd11; b_sign2 = 4'd9; b_sign3 = 4'd10;
@(posedge clk_i);
shared_exps0 = 8'd129;
shared_exps1 = 8'd122;
rstn = 0;
@(posedge clk_i);
rstn = 1;
a_mant0 = 8'd1; a_mant1 = 8'd11; a_mant2 = 8'd229; a_mant3 = 8'd104;
b_mant0 = 8'd235; b_mant1 = 8'd248; b_mant2 = 8'd192; b_mant3 = 8'd238;
a_exp0 = 10'd568; a_exp1 = 10'd946; a_exp2 = 10'd403; a_exp3 = 10'd639;
b_exp0 = 10'd992; b_exp1 = 10'd744; b_exp2 = 10'd62; b_exp3 = 10'd487;
a_sign0 = 4'd1; a_sign1 = 4'd12; a_sign2 = 4'd5; a_sign3 = 4'd4;
b_sign0 = 4'd10; b_sign1 = 4'd8; b_sign2 = 4'd4; b_sign3 = 4'd2;
@(posedge clk_i);
a_mant0 = 8'd80; a_mant1 = 8'd150; a_mant2 = 8'd101; a_mant3 = 8'd215;
b_mant0 = 8'd140; b_mant1 = 8'd173; b_mant2 = 8'd130; b_mant3 = 8'd207;
a_exp0 = 10'd719; a_exp1 = 10'd199; a_exp2 = 10'd401; a_exp3 = 10'd212;
b_exp0 = 10'd794; b_exp1 = 10'd348; b_exp2 = 10'd942; b_exp3 = 10'd117;
a_sign0 = 4'd6; a_sign1 = 4'd8; a_sign2 = 4'd10; a_sign3 = 4'd9;
b_sign0 = 4'd2; b_sign1 = 4'd14; b_sign2 = 4'd13; b_sign3 = 4'd13;
@(posedge clk_i);
a_mant0 = 8'd181; a_mant1 = 8'd33; a_mant2 = 8'd221; a_mant3 = 8'd88;
b_mant0 = 8'd82; b_mant1 = 8'd198; b_mant2 = 8'd14; b_mant3 = 8'd54;
a_exp0 = 10'd779; a_exp1 = 10'd336; a_exp2 = 10'd732; a_exp3 = 10'd952;
b_exp0 = 10'd303; b_exp1 = 10'd414; b_exp2 = 10'd846; b_exp3 = 10'd851;
a_sign0 = 4'd6; a_sign1 = 4'd3; a_sign2 = 4'd10; a_sign3 = 4'd7;
b_sign0 = 4'd2; b_sign1 = 4'd10; b_sign2 = 4'd5; b_sign3 = 4'd7;
@(posedge clk_i);
a_mant0 = 8'd34; a_mant1 = 8'd236; a_mant2 = 8'd214; a_mant3 = 8'd171;
b_mant0 = 8'd26; b_mant1 = 8'd219; b_mant2 = 8'd46; b_mant3 = 8'd175;
a_exp0 = 10'd552; a_exp1 = 10'd864; a_exp2 = 10'd946; a_exp3 = 10'd869;
b_exp0 = 10'd849; b_exp1 = 10'd260; b_exp2 = 10'd594; b_exp3 = 10'd171;
a_sign0 = 4'd1; a_sign1 = 4'd6; a_sign2 = 4'd5; a_sign3 = 4'd15;
b_sign0 = 4'd1; b_sign1 = 4'd7; b_sign2 = 4'd0; b_sign3 = 4'd1;
@(posedge clk_i);
a_mant0 = 8'd232; a_mant1 = 8'd66; a_mant2 = 8'd118; a_mant3 = 8'd13;
b_mant0 = 8'd221; b_mant1 = 8'd167; b_mant2 = 8'd241; b_mant3 = 8'd1;
a_exp0 = 10'd688; a_exp1 = 10'd220; a_exp2 = 10'd385; a_exp3 = 10'd807;
b_exp0 = 10'd208; b_exp1 = 10'd33; b_exp2 = 10'd439; b_exp3 = 10'd65;
a_sign0 = 4'd4; a_sign1 = 4'd10; a_sign2 = 4'd15; a_sign3 = 4'd1;
b_sign0 = 4'd8; b_sign1 = 4'd5; b_sign2 = 4'd0; b_sign3 = 4'd6;
@(posedge clk_i);
a_mant0 = 8'd99; a_mant1 = 8'd31; a_mant2 = 8'd249; a_mant3 = 8'd31;
b_mant0 = 8'd24; b_mant1 = 8'd171; b_mant2 = 8'd201; b_mant3 = 8'd227;
a_exp0 = 10'd80; a_exp1 = 10'd559; a_exp2 = 10'd845; a_exp3 = 10'd46;
b_exp0 = 10'd53; b_exp1 = 10'd746; b_exp2 = 10'd354; b_exp3 = 10'd760;
a_sign0 = 4'd12; a_sign1 = 4'd8; a_sign2 = 4'd2; a_sign3 = 4'd10;
b_sign0 = 4'd10; b_sign1 = 4'd13; b_sign2 = 4'd6; b_sign3 = 4'd14;
@(posedge clk_i);
a_mant0 = 8'd250; a_mant1 = 8'd22; a_mant2 = 8'd233; a_mant3 = 8'd109;
b_mant0 = 8'd136; b_mant1 = 8'd136; b_mant2 = 8'd156; b_mant3 = 8'd183;
a_exp0 = 10'd359; a_exp1 = 10'd129; a_exp2 = 10'd261; a_exp3 = 10'd288;
b_exp0 = 10'd185; b_exp1 = 10'd181; b_exp2 = 10'd276; b_exp3 = 10'd232;
a_sign0 = 4'd5; a_sign1 = 4'd2; a_sign2 = 4'd1; a_sign3 = 4'd14;
b_sign0 = 4'd14; b_sign1 = 4'd8; b_sign2 = 4'd16; b_sign3 = 4'd1;
@(posedge clk_i);
shared_exps0 = 8'd134;
shared_exps1 = 8'd132;
a_mant0 = 8'd30; a_mant1 = 8'd48; a_mant2 = 8'd94; a_mant3 = 8'd188;
b_mant0 = 8'd225; b_mant1 = 8'd166; b_mant2 = 8'd223; b_mant3 = 8'd105;
a_exp0 = 10'd117; a_exp1 = 10'd328; a_exp2 = 10'd992; a_exp3 = 10'd83;
b_exp0 = 10'd109; b_exp1 = 10'd837; b_exp2 = 10'd570; b_exp3 = 10'd733;
a_sign0 = 4'd6; a_sign1 = 4'd15; a_sign2 = 4'd14; a_sign3 = 4'd4;
b_sign0 = 4'd3; b_sign1 = 4'd12; b_sign2 = 4'd0; b_sign3 = 4'd5;
@(posedge clk_i);
a_mant0 = 8'd209; a_mant1 = 8'd70; a_mant2 = 8'd183; a_mant3 = 8'd146;
b_mant0 = 8'd64; b_mant1 = 8'd80; b_mant2 = 8'd27; b_mant3 = 8'd234;
a_exp0 = 10'd832; a_exp1 = 10'd578; a_exp2 = 10'd739; a_exp3 = 10'd901;
b_exp0 = 10'd89; b_exp1 = 10'd4; b_exp2 = 10'd12; b_exp3 = 10'd848;
a_sign0 = 4'd6; a_sign1 = 4'd4; a_sign2 = 4'd15; a_sign3 = 4'd13;
b_sign0 = 4'd6; b_sign1 = 4'd6; b_sign2 = 4'd16; b_sign3 = 4'd9;
@(posedge clk_i);
a_mant0 = 8'd95; a_mant1 = 8'd254; a_mant2 = 8'd135; a_mant3 = 8'd57;
b_mant0 = 8'd101; b_mant1 = 8'd44; b_mant2 = 8'd114; b_mant3 = 8'd174;
a_exp0 = 10'd261; a_exp1 = 10'd353; a_exp2 = 10'd279; a_exp3 = 10'd1018;
b_exp0 = 10'd426; b_exp1 = 10'd805; b_exp2 = 10'd190; b_exp3 = 10'd519;
a_sign0 = 4'd7; a_sign1 = 4'd5; a_sign2 = 4'd5; a_sign3 = 4'd5;
b_sign0 = 4'd2; b_sign1 = 4'd10; b_sign2 = 4'd14; b_sign3 = 4'd15;
@(posedge clk_i);
a_mant0 = 8'd102; a_mant1 = 8'd213; a_mant2 = 8'd37; a_mant3 = 8'd117;
b_mant0 = 8'd60; b_mant1 = 8'd155; b_mant2 = 8'd46; b_mant3 = 8'd183;
a_exp0 = 10'd796; a_exp1 = 10'd459; a_exp2 = 10'd28; a_exp3 = 10'd688;
b_exp0 = 10'd302; b_exp1 = 10'd415; b_exp2 = 10'd997; b_exp3 = 10'd167;
a_sign0 = 4'd4; a_sign1 = 4'd7; a_sign2 = 4'd9; a_sign3 = 4'd4;
b_sign0 = 4'd0; b_sign1 = 4'd0; b_sign2 = 4'd14; b_sign3 = 4'd7;
@(posedge clk_i);
a_mant0 = 8'd85; a_mant1 = 8'd205; a_mant2 = 8'd192; a_mant3 = 8'd12;
b_mant0 = 8'd197; b_mant1 = 8'd132; b_mant2 = 8'd154; b_mant3 = 8'd150;
a_exp0 = 10'd905; a_exp1 = 10'd435; a_exp2 = 10'd741; a_exp3 = 10'd975;
b_exp0 = 10'd293; b_exp1 = 10'd273; b_exp2 = 10'd976; b_exp3 = 10'd236;
a_sign0 = 4'd12; a_sign1 = 4'd12; a_sign2 = 4'd6; a_sign3 = 4'd0;
b_sign0 = 4'd7; b_sign1 = 4'd13; b_sign2 = 4'd14; b_sign3 = 4'd9;
@(posedge clk_i);
a_mant0 = 8'd40; a_mant1 = 8'd234; a_mant2 = 8'd223; a_mant3 = 8'd21;
b_mant0 = 8'd96; b_mant1 = 8'd243; b_mant2 = 8'd193; b_mant3 = 8'd231;
a_exp0 = 10'd759; a_exp1 = 10'd786; a_exp2 = 10'd205; a_exp3 = 10'd613;
b_exp0 = 10'd566; b_exp1 = 10'd470; b_exp2 = 10'd768; b_exp3 = 10'd366;
a_sign0 = 4'd2; a_sign1 = 4'd6; a_sign2 = 4'd16; a_sign3 = 4'd8;
b_sign0 = 4'd8; b_sign1 = 4'd15; b_sign2 = 4'd15; b_sign3 = 4'd5;
@(posedge clk_i);
a_mant0 = 8'd170; a_mant1 = 8'd77; a_mant2 = 8'd216; a_mant3 = 8'd55;
b_mant0 = 8'd1; b_mant1 = 8'd204; b_mant2 = 8'd105; b_mant3 = 8'd84;
a_exp0 = 10'd101; a_exp1 = 10'd95; a_exp2 = 10'd994; a_exp3 = 10'd1017;
b_exp0 = 10'd731; b_exp1 = 10'd128; b_exp2 = 10'd157; b_exp3 = 10'd979;
a_sign0 = 4'd5; a_sign1 = 4'd9; a_sign2 = 4'd13; a_sign3 = 4'd7;
b_sign0 = 4'd15; b_sign1 = 4'd12; b_sign2 = 4'd16; b_sign3 = 4'd3;
@(posedge clk_i);
a_mant0 = 8'd176; a_mant1 = 8'd138; a_mant2 = 8'd212; a_mant3 = 8'd237;
b_mant0 = 8'd209; b_mant1 = 8'd151; b_mant2 = 8'd67; b_mant3 = 8'd153;
a_exp0 = 10'd66; a_exp1 = 10'd976; a_exp2 = 10'd532; a_exp3 = 10'd384;
b_exp0 = 10'd39; b_exp1 = 10'd276; b_exp2 = 10'd284; b_exp3 = 10'd175;
a_sign0 = 4'd1; a_sign1 = 4'd16; a_sign2 = 4'd11; a_sign3 = 4'd16;
b_sign0 = 4'd8; b_sign1 = 4'd3; b_sign2 = 4'd5; b_sign3 = 4'd11;
@(posedge clk_i);
shared_exps0 = 8'd128;
shared_exps1 = 8'd145;
a_mant0 = 8'd36; a_mant1 = 8'd60; a_mant2 = 8'd43; a_mant3 = 8'd173;
b_mant0 = 8'd34; b_mant1 = 8'd211; b_mant2 = 8'd109; b_mant3 = 8'd174;
a_exp0 = 10'd214; a_exp1 = 10'd550; a_exp2 = 10'd32; a_exp3 = 10'd769;
b_exp0 = 10'd162; b_exp1 = 10'd262; b_exp2 = 10'd669; b_exp3 = 10'd311;
a_sign0 = 4'd3; a_sign1 = 4'd8; a_sign2 = 4'd0; a_sign3 = 4'd7;
b_sign0 = 4'd14; b_sign1 = 4'd13; b_sign2 = 4'd8; b_sign3 = 4'd13;
@(posedge clk_i);
a_mant0 = 8'd17; a_mant1 = 8'd204; a_mant2 = 8'd182; a_mant3 = 8'd142;
b_mant0 = 8'd44; b_mant1 = 8'd63; b_mant2 = 8'd213; b_mant3 = 8'd128;
a_exp0 = 10'd525; a_exp1 = 10'd58; a_exp2 = 10'd999; a_exp3 = 10'd22;
b_exp0 = 10'd150; b_exp1 = 10'd776; b_exp2 = 10'd415; b_exp3 = 10'd100;
a_sign0 = 4'd0; a_sign1 = 4'd4; a_sign2 = 4'd16; a_sign3 = 4'd13;
b_sign0 = 4'd15; b_sign1 = 4'd5; b_sign2 = 4'd8; b_sign3 = 4'd5;
@(posedge clk_i);
a_mant0 = 8'd154; a_mant1 = 8'd225; a_mant2 = 8'd35; a_mant3 = 8'd186;
b_mant0 = 8'd212; b_mant1 = 8'd118; b_mant2 = 8'd35; b_mant3 = 8'd70;
a_exp0 = 10'd883; a_exp1 = 10'd77; a_exp2 = 10'd739; a_exp3 = 10'd543;
b_exp0 = 10'd185; b_exp1 = 10'd538; b_exp2 = 10'd14; b_exp3 = 10'd9;
a_sign0 = 4'd15; a_sign1 = 4'd9; a_sign2 = 4'd0; a_sign3 = 4'd11;
b_sign0 = 4'd12; b_sign1 = 4'd5; b_sign2 = 4'd12; b_sign3 = 4'd4;
@(posedge clk_i);
a_mant0 = 8'd246; a_mant1 = 8'd188; a_mant2 = 8'd148; a_mant3 = 8'd126;
b_mant0 = 8'd44; b_mant1 = 8'd213; b_mant2 = 8'd49; b_mant3 = 8'd107;
a_exp0 = 10'd438; a_exp1 = 10'd743; a_exp2 = 10'd193; a_exp3 = 10'd289;
b_exp0 = 10'd775; b_exp1 = 10'd83; b_exp2 = 10'd17; b_exp3 = 10'd515;
a_sign0 = 4'd9; a_sign1 = 4'd7; a_sign2 = 4'd5; a_sign3 = 4'd16;
b_sign0 = 4'd10; b_sign1 = 4'd0; b_sign2 = 4'd5; b_sign3 = 4'd2;
@(posedge clk_i);
a_mant0 = 8'd229; a_mant1 = 8'd235; a_mant2 = 8'd4; a_mant3 = 8'd196;
b_mant0 = 8'd204; b_mant1 = 8'd11; b_mant2 = 8'd138; b_mant3 = 8'd63;
a_exp0 = 10'd236; a_exp1 = 10'd338; a_exp2 = 10'd667; a_exp3 = 10'd166;
b_exp0 = 10'd427; b_exp1 = 10'd531; b_exp2 = 10'd157; b_exp3 = 10'd951;
a_sign0 = 4'd7; a_sign1 = 4'd14; a_sign2 = 4'd6; a_sign3 = 4'd16;
b_sign0 = 4'd3; b_sign1 = 4'd7; b_sign2 = 4'd6; b_sign3 = 4'd4;
@(posedge clk_i);
a_mant0 = 8'd173; a_mant1 = 8'd64; a_mant2 = 8'd49; a_mant3 = 8'd73;
b_mant0 = 8'd33; b_mant1 = 8'd241; b_mant2 = 8'd158; b_mant3 = 8'd103;
a_exp0 = 10'd694; a_exp1 = 10'd275; a_exp2 = 10'd242; a_exp3 = 10'd623;
b_exp0 = 10'd386; b_exp1 = 10'd866; b_exp2 = 10'd291; b_exp3 = 10'd151;
a_sign0 = 4'd4; a_sign1 = 4'd16; a_sign2 = 4'd1; a_sign3 = 4'd5;
b_sign0 = 4'd0; b_sign1 = 4'd15; b_sign2 = 4'd11; b_sign3 = 4'd7;
@(posedge clk_i);
a_mant0 = 8'd210; a_mant1 = 8'd168; a_mant2 = 8'd154; a_mant3 = 8'd14;
b_mant0 = 8'd206; b_mant1 = 8'd48; b_mant2 = 8'd187; b_mant3 = 8'd189;
a_exp0 = 10'd926; a_exp1 = 10'd669; a_exp2 = 10'd571; a_exp3 = 10'd25;
b_exp0 = 10'd386; b_exp1 = 10'd396; b_exp2 = 10'd117; b_exp3 = 10'd140;
a_sign0 = 4'd12; a_sign1 = 4'd13; a_sign2 = 4'd5; a_sign3 = 4'd13;
b_sign0 = 4'd16; b_sign1 = 4'd3; b_sign2 = 4'd4; b_sign3 = 4'd3;
@(posedge clk_i);
a_mant0 = 8'd170; a_mant1 = 8'd126; a_mant2 = 8'd12; a_mant3 = 8'd225;
b_mant0 = 8'd97; b_mant1 = 8'd57; b_mant2 = 8'd192; b_mant3 = 8'd234;
a_exp0 = 10'd70; a_exp1 = 10'd195; a_exp2 = 10'd508; a_exp3 = 10'd908;
b_exp0 = 10'd225; b_exp1 = 10'd642; b_exp2 = 10'd382; b_exp3 = 10'd143;
a_sign0 = 4'd10; a_sign1 = 4'd13; a_sign2 = 4'd14; a_sign3 = 4'd3;
b_sign0 = 4'd3; b_sign1 = 4'd15; b_sign2 = 4'd10; b_sign3 = 4'd1;
@(posedge clk_i);
shared_exps0 = 8'd130;
shared_exps1 = 8'd85;
a_mant0 = 8'd178; a_mant1 = 8'd187; a_mant2 = 8'd148; a_mant3 = 8'd97;
b_mant0 = 8'd196; b_mant1 = 8'd123; b_mant2 = 8'd255; b_mant3 = 8'd212;
a_exp0 = 10'd292; a_exp1 = 10'd882; a_exp2 = 10'd964; a_exp3 = 10'd272;
b_exp0 = 10'd16; b_exp1 = 10'd614; b_exp2 = 10'd240; b_exp3 = 10'd270;
a_sign0 = 4'd13; a_sign1 = 4'd14; a_sign2 = 4'd16; a_sign3 = 4'd2;
b_sign0 = 4'd6; b_sign1 = 4'd10; b_sign2 = 4'd12; b_sign3 = 4'd16;
@(posedge clk_i);
a_mant0 = 8'd165; a_mant1 = 8'd142; a_mant2 = 8'd165; a_mant3 = 8'd82;
b_mant0 = 8'd236; b_mant1 = 8'd115; b_mant2 = 8'd171; b_mant3 = 8'd3;
a_exp0 = 10'd996; a_exp1 = 10'd743; a_exp2 = 10'd616; a_exp3 = 10'd960;
b_exp0 = 10'd633; b_exp1 = 10'd785; b_exp2 = 10'd345; b_exp3 = 10'd789;
a_sign0 = 4'd8; a_sign1 = 4'd5; a_sign2 = 4'd9; a_sign3 = 4'd12;
b_sign0 = 4'd5; b_sign1 = 4'd10; b_sign2 = 4'd4; b_sign3 = 4'd8;
@(posedge clk_i);
a_mant0 = 8'd60; a_mant1 = 8'd70; a_mant2 = 8'd129; a_mant3 = 8'd98;
b_mant0 = 8'd83; b_mant1 = 8'd254; b_mant2 = 8'd167; b_mant3 = 8'd58;
a_exp0 = 10'd616; a_exp1 = 10'd617; a_exp2 = 10'd1008; a_exp3 = 10'd354;
b_exp0 = 10'd382; b_exp1 = 10'd955; b_exp2 = 10'd705; b_exp3 = 10'd489;
a_sign0 = 4'd1; a_sign1 = 4'd12; a_sign2 = 4'd5; a_sign3 = 4'd9;
b_sign0 = 4'd13; b_sign1 = 4'd15; b_sign2 = 4'd2; b_sign3 = 4'd4;
@(posedge clk_i);
a_mant0 = 8'd207; a_mant1 = 8'd18; a_mant2 = 8'd232; a_mant3 = 8'd170;
b_mant0 = 8'd160; b_mant1 = 8'd118; b_mant2 = 8'd67; b_mant3 = 8'd218;
a_exp0 = 10'd361; a_exp1 = 10'd207; a_exp2 = 10'd186; a_exp3 = 10'd411;
b_exp0 = 10'd380; b_exp1 = 10'd977; b_exp2 = 10'd237; b_exp3 = 10'd842;
a_sign0 = 4'd2; a_sign1 = 4'd16; a_sign2 = 4'd7; a_sign3 = 4'd2;
b_sign0 = 4'd13; b_sign1 = 4'd13; b_sign2 = 4'd14; b_sign3 = 4'd2;
@(posedge clk_i);
a_mant0 = 8'd80; a_mant1 = 8'd70; a_mant2 = 8'd88; a_mant3 = 8'd7;
b_mant0 = 8'd117; b_mant1 = 8'd217; b_mant2 = 8'd218; b_mant3 = 8'd30;
a_exp0 = 10'd247; a_exp1 = 10'd924; a_exp2 = 10'd989; a_exp3 = 10'd981;
b_exp0 = 10'd620; b_exp1 = 10'd420; b_exp2 = 10'd199; b_exp3 = 10'd731;
a_sign0 = 4'd12; a_sign1 = 4'd15; a_sign2 = 4'd11; a_sign3 = 4'd7;
b_sign0 = 4'd5; b_sign1 = 4'd10; b_sign2 = 4'd10; b_sign3 = 4'd8;
@(posedge clk_i);
a_mant0 = 8'd183; a_mant1 = 8'd151; a_mant2 = 8'd140; a_mant3 = 8'd228;
b_mant0 = 8'd80; b_mant1 = 8'd217; b_mant2 = 8'd122; b_mant3 = 8'd235;
a_exp0 = 10'd923; a_exp1 = 10'd44; a_exp2 = 10'd120; a_exp3 = 10'd696;
b_exp0 = 10'd43; b_exp1 = 10'd388; b_exp2 = 10'd244; b_exp3 = 10'd581;
a_sign0 = 4'd10; a_sign1 = 4'd2; a_sign2 = 4'd9; a_sign3 = 4'd11;
b_sign0 = 4'd3; b_sign1 = 4'd14; b_sign2 = 4'd6; b_sign3 = 4'd16;
@(posedge clk_i);
a_mant0 = 8'd245; a_mant1 = 8'd69; a_mant2 = 8'd96; a_mant3 = 8'd181;
b_mant0 = 8'd147; b_mant1 = 8'd194; b_mant2 = 8'd215; b_mant3 = 8'd185;
a_exp0 = 10'd873; a_exp1 = 10'd940; a_exp2 = 10'd301; a_exp3 = 10'd648;
b_exp0 = 10'd458; b_exp1 = 10'd923; b_exp2 = 10'd912; b_exp3 = 10'd636;
a_sign0 = 4'd9; a_sign1 = 4'd8; a_sign2 = 4'd4; a_sign3 = 4'd10;
b_sign0 = 4'd4; b_sign1 = 4'd8; b_sign2 = 4'd6; b_sign3 = 4'd2;
@(posedge clk_i);
a_mant0 = 8'd74; a_mant1 = 8'd221; a_mant2 = 8'd23; a_mant3 = 8'd223;
b_mant0 = 8'd165; b_mant1 = 8'd180; b_mant2 = 8'd185; b_mant3 = 8'd200;
a_exp0 = 10'd964; a_exp1 = 10'd189; a_exp2 = 10'd747; a_exp3 = 10'd1000;
b_exp0 = 10'd23; b_exp1 = 10'd310; b_exp2 = 10'd411; b_exp3 = 10'd846;
a_sign0 = 4'd16; a_sign1 = 4'd10; a_sign2 = 4'd3; a_sign3 = 4'd1;
b_sign0 = 4'd1; b_sign1 = 4'd13; b_sign2 = 4'd4; b_sign3 = 4'd2;
@(posedge clk_i);
shared_exps0 = 8'd157;
shared_exps1 = 8'd136;
rstn = 0;
@(posedge clk_i);
rstn = 1;
a_mant0 = 8'd219; a_mant1 = 8'd52; a_mant2 = 8'd151; a_mant3 = 8'd151;
b_mant0 = 8'd28; b_mant1 = 8'd106; b_mant2 = 8'd103; b_mant3 = 8'd199;
a_exp0 = 10'd38; a_exp1 = 10'd904; a_exp2 = 10'd182; a_exp3 = 10'd514;
b_exp0 = 10'd904; b_exp1 = 10'd908; b_exp2 = 10'd960; b_exp3 = 10'd506;
a_sign0 = 4'd4; a_sign1 = 4'd13; a_sign2 = 4'd3; a_sign3 = 4'd16;
b_sign0 = 4'd2; b_sign1 = 4'd2; b_sign2 = 4'd10; b_sign3 = 4'd16;
@(posedge clk_i);
a_mant0 = 8'd114; a_mant1 = 8'd220; a_mant2 = 8'd49; a_mant3 = 8'd25;
b_mant0 = 8'd108; b_mant1 = 8'd17; b_mant2 = 8'd100; b_mant3 = 8'd96;
a_exp0 = 10'd418; a_exp1 = 10'd86; a_exp2 = 10'd1013; a_exp3 = 10'd562;
b_exp0 = 10'd700; b_exp1 = 10'd748; b_exp2 = 10'd842; b_exp3 = 10'd402;
a_sign0 = 4'd4; a_sign1 = 4'd16; a_sign2 = 4'd12; a_sign3 = 4'd10;
b_sign0 = 4'd7; b_sign1 = 4'd10; b_sign2 = 4'd16; b_sign3 = 4'd5;
@(posedge clk_i);
a_mant0 = 8'd167; a_mant1 = 8'd222; a_mant2 = 8'd11; a_mant3 = 8'd154;
b_mant0 = 8'd1; b_mant1 = 8'd253; b_mant2 = 8'd113; b_mant3 = 8'd191;
a_exp0 = 10'd395; a_exp1 = 10'd40; a_exp2 = 10'd62; a_exp3 = 10'd838;
b_exp0 = 10'd1002; b_exp1 = 10'd53; b_exp2 = 10'd313; b_exp3 = 10'd44;
a_sign0 = 4'd6; a_sign1 = 4'd3; a_sign2 = 4'd16; a_sign3 = 4'd11;
b_sign0 = 4'd7; b_sign1 = 4'd14; b_sign2 = 4'd11; b_sign3 = 4'd8;
@(posedge clk_i);
a_mant0 = 8'd58; a_mant1 = 8'd163; a_mant2 = 8'd131; a_mant3 = 8'd85;
b_mant0 = 8'd228; b_mant1 = 8'd251; b_mant2 = 8'd30; b_mant3 = 8'd88;
a_exp0 = 10'd732; a_exp1 = 10'd548; a_exp2 = 10'd67; a_exp3 = 10'd899;
b_exp0 = 10'd119; b_exp1 = 10'd329; b_exp2 = 10'd378; b_exp3 = 10'd584;
a_sign0 = 4'd0; a_sign1 = 4'd14; a_sign2 = 4'd5; a_sign3 = 4'd7;
b_sign0 = 4'd6; b_sign1 = 4'd16; b_sign2 = 4'd11; b_sign3 = 4'd5;
@(posedge clk_i);
a_mant0 = 8'd151; a_mant1 = 8'd244; a_mant2 = 8'd92; a_mant3 = 8'd36;
b_mant0 = 8'd254; b_mant1 = 8'd40; b_mant2 = 8'd211; b_mant3 = 8'd92;
a_exp0 = 10'd130; a_exp1 = 10'd84; a_exp2 = 10'd281; a_exp3 = 10'd181;
b_exp0 = 10'd39; b_exp1 = 10'd8; b_exp2 = 10'd978; b_exp3 = 10'd636;
a_sign0 = 4'd1; a_sign1 = 4'd14; a_sign2 = 4'd10; a_sign3 = 4'd16;
b_sign0 = 4'd1; b_sign1 = 4'd8; b_sign2 = 4'd1; b_sign3 = 4'd11;
@(posedge clk_i);
a_mant0 = 8'd138; a_mant1 = 8'd57; a_mant2 = 8'd133; a_mant3 = 8'd24;
b_mant0 = 8'd7; b_mant1 = 8'd59; b_mant2 = 8'd237; b_mant3 = 8'd141;
a_exp0 = 10'd875; a_exp1 = 10'd526; a_exp2 = 10'd68; a_exp3 = 10'd555;
b_exp0 = 10'd990; b_exp1 = 10'd953; b_exp2 = 10'd238; b_exp3 = 10'd152;
a_sign0 = 4'd7; a_sign1 = 4'd3; a_sign2 = 4'd4; a_sign3 = 4'd10;
b_sign0 = 4'd0; b_sign1 = 4'd8; b_sign2 = 4'd0; b_sign3 = 4'd7;
@(posedge clk_i);
a_mant0 = 8'd168; a_mant1 = 8'd68; a_mant2 = 8'd56; a_mant3 = 8'd232;
b_mant0 = 8'd168; b_mant1 = 8'd236; b_mant2 = 8'd177; b_mant3 = 8'd204;
a_exp0 = 10'd333; a_exp1 = 10'd656; a_exp2 = 10'd671; a_exp3 = 10'd754;
b_exp0 = 10'd61; b_exp1 = 10'd444; b_exp2 = 10'd871; b_exp3 = 10'd89;
a_sign0 = 4'd13; a_sign1 = 4'd7; a_sign2 = 4'd3; a_sign3 = 4'd9;
b_sign0 = 4'd12; b_sign1 = 4'd12; b_sign2 = 4'd2; b_sign3 = 4'd11;
@(posedge clk_i);
shared_exps0 = 8'd121;
shared_exps1 = 8'd107;
a_mant0 = 8'd104; a_mant1 = 8'd61; a_mant2 = 8'd199; a_mant3 = 8'd114;
b_mant0 = 8'd52; b_mant1 = 8'd36; b_mant2 = 8'd226; b_mant3 = 8'd114;
a_exp0 = 10'd97; a_exp1 = 10'd1017; a_exp2 = 10'd652; a_exp3 = 10'd779;
b_exp0 = 10'd328; b_exp1 = 10'd930; b_exp2 = 10'd359; b_exp3 = 10'd67;
a_sign0 = 4'd4; a_sign1 = 4'd13; a_sign2 = 4'd10; a_sign3 = 4'd2;
b_sign0 = 4'd7; b_sign1 = 4'd10; b_sign2 = 4'd0; b_sign3 = 4'd1;
@(posedge clk_i);
a_mant0 = 8'd215; a_mant1 = 8'd3; a_mant2 = 8'd183; a_mant3 = 8'd152;
b_mant0 = 8'd80; b_mant1 = 8'd69; b_mant2 = 8'd178; b_mant3 = 8'd168;
a_exp0 = 10'd718; a_exp1 = 10'd676; a_exp2 = 10'd328; a_exp3 = 10'd123;
b_exp0 = 10'd899; b_exp1 = 10'd248; b_exp2 = 10'd281; b_exp3 = 10'd90;
a_sign0 = 4'd11; a_sign1 = 4'd16; a_sign2 = 4'd14; a_sign3 = 4'd1;
b_sign0 = 4'd4; b_sign1 = 4'd5; b_sign2 = 4'd6; b_sign3 = 4'd16;
@(posedge clk_i);
a_mant0 = 8'd20; a_mant1 = 8'd54; a_mant2 = 8'd174; a_mant3 = 8'd155;
b_mant0 = 8'd180; b_mant1 = 8'd218; b_mant2 = 8'd119; b_mant3 = 8'd247;
a_exp0 = 10'd101; a_exp1 = 10'd144; a_exp2 = 10'd20; a_exp3 = 10'd12;
b_exp0 = 10'd695; b_exp1 = 10'd259; b_exp2 = 10'd400; b_exp3 = 10'd78;
a_sign0 = 4'd15; a_sign1 = 4'd4; a_sign2 = 4'd0; a_sign3 = 4'd3;
b_sign0 = 4'd12; b_sign1 = 4'd16; b_sign2 = 4'd15; b_sign3 = 4'd2;
@(posedge clk_i);
a_mant0 = 8'd159; a_mant1 = 8'd67; a_mant2 = 8'd27; a_mant3 = 8'd0;
b_mant0 = 8'd20; b_mant1 = 8'd221; b_mant2 = 8'd206; b_mant3 = 8'd82;
a_exp0 = 10'd844; a_exp1 = 10'd1009; a_exp2 = 10'd811; a_exp3 = 10'd620;
b_exp0 = 10'd705; b_exp1 = 10'd45; b_exp2 = 10'd835; b_exp3 = 10'd50;
a_sign0 = 4'd0; a_sign1 = 4'd15; a_sign2 = 4'd12; a_sign3 = 4'd6;
b_sign0 = 4'd16; b_sign1 = 4'd7; b_sign2 = 4'd11; b_sign3 = 4'd14;
@(posedge clk_i);
a_mant0 = 8'd110; a_mant1 = 8'd148; a_mant2 = 8'd240; a_mant3 = 8'd224;
b_mant0 = 8'd193; b_mant1 = 8'd107; b_mant2 = 8'd202; b_mant3 = 8'd247;
a_exp0 = 10'd188; a_exp1 = 10'd123; a_exp2 = 10'd141; a_exp3 = 10'd34;
b_exp0 = 10'd89; b_exp1 = 10'd935; b_exp2 = 10'd236; b_exp3 = 10'd579;
a_sign0 = 4'd11; a_sign1 = 4'd7; a_sign2 = 4'd10; a_sign3 = 4'd10;
b_sign0 = 4'd8; b_sign1 = 4'd2; b_sign2 = 4'd9; b_sign3 = 4'd13;
@(posedge clk_i);
a_mant0 = 8'd164; a_mant1 = 8'd94; a_mant2 = 8'd21; a_mant3 = 8'd133;
b_mant0 = 8'd3; b_mant1 = 8'd198; b_mant2 = 8'd174; b_mant3 = 8'd103;
a_exp0 = 10'd14; a_exp1 = 10'd656; a_exp2 = 10'd119; a_exp3 = 10'd565;
b_exp0 = 10'd961; b_exp1 = 10'd463; b_exp2 = 10'd648; b_exp3 = 10'd318;
a_sign0 = 4'd16; a_sign1 = 4'd8; a_sign2 = 4'd6; a_sign3 = 4'd9;
b_sign0 = 4'd14; b_sign1 = 4'd15; b_sign2 = 4'd13; b_sign3 = 4'd15;
@(posedge clk_i);
a_mant0 = 8'd15; a_mant1 = 8'd187; a_mant2 = 8'd163; a_mant3 = 8'd86;
b_mant0 = 8'd153; b_mant1 = 8'd193; b_mant2 = 8'd143; b_mant3 = 8'd73;
a_exp0 = 10'd772; a_exp1 = 10'd482; a_exp2 = 10'd24; a_exp3 = 10'd936;
b_exp0 = 10'd329; b_exp1 = 10'd84; b_exp2 = 10'd325; b_exp3 = 10'd452;
a_sign0 = 4'd4; a_sign1 = 4'd10; a_sign2 = 4'd13; a_sign3 = 4'd16;
b_sign0 = 4'd9; b_sign1 = 4'd16; b_sign2 = 4'd3; b_sign3 = 4'd9;
@(posedge clk_i);
a_mant0 = 8'd206; a_mant1 = 8'd75; a_mant2 = 8'd122; a_mant3 = 8'd157;
b_mant0 = 8'd191; b_mant1 = 8'd60; b_mant2 = 8'd125; b_mant3 = 8'd252;
a_exp0 = 10'd83; a_exp1 = 10'd624; a_exp2 = 10'd880; a_exp3 = 10'd268;
b_exp0 = 10'd947; b_exp1 = 10'd164; b_exp2 = 10'd287; b_exp3 = 10'd474;
a_sign0 = 4'd8; a_sign1 = 4'd7; a_sign2 = 4'd7; a_sign3 = 4'd12;
b_sign0 = 4'd11; b_sign1 = 4'd15; b_sign2 = 4'd9; b_sign3 = 4'd3;
@(posedge clk_i);
shared_exps0 = 8'd110;
shared_exps1 = 8'd143;
a_mant0 = 8'd3; a_mant1 = 8'd180; a_mant2 = 8'd168; a_mant3 = 8'd250;
b_mant0 = 8'd211; b_mant1 = 8'd167; b_mant2 = 8'd3; b_mant3 = 8'd63;
a_exp0 = 10'd67; a_exp1 = 10'd197; a_exp2 = 10'd941; a_exp3 = 10'd352;
b_exp0 = 10'd387; b_exp1 = 10'd682; b_exp2 = 10'd158; b_exp3 = 10'd493;
a_sign0 = 4'd13; a_sign1 = 4'd8; a_sign2 = 4'd15; a_sign3 = 4'd6;
b_sign0 = 4'd9; b_sign1 = 4'd16; b_sign2 = 4'd13; b_sign3 = 4'd0;
@(posedge clk_i);
a_mant0 = 8'd75; a_mant1 = 8'd180; a_mant2 = 8'd214; a_mant3 = 8'd89;
b_mant0 = 8'd88; b_mant1 = 8'd204; b_mant2 = 8'd58; b_mant3 = 8'd171;
a_exp0 = 10'd186; a_exp1 = 10'd842; a_exp2 = 10'd630; a_exp3 = 10'd205;
b_exp0 = 10'd395; b_exp1 = 10'd376; b_exp2 = 10'd774; b_exp3 = 10'd895;
a_sign0 = 4'd16; a_sign1 = 4'd16; a_sign2 = 4'd5; a_sign3 = 4'd7;
b_sign0 = 4'd4; b_sign1 = 4'd3; b_sign2 = 4'd6; b_sign3 = 4'd16;
@(posedge clk_i);
a_mant0 = 8'd177; a_mant1 = 8'd199; a_mant2 = 8'd186; a_mant3 = 8'd233;
b_mant0 = 8'd1; b_mant1 = 8'd242; b_mant2 = 8'd166; b_mant3 = 8'd51;
a_exp0 = 10'd308; a_exp1 = 10'd191; a_exp2 = 10'd430; a_exp3 = 10'd817;
b_exp0 = 10'd987; b_exp1 = 10'd350; b_exp2 = 10'd1008; b_exp3 = 10'd975;
a_sign0 = 4'd11; a_sign1 = 4'd8; a_sign2 = 4'd6; a_sign3 = 4'd3;
b_sign0 = 4'd0; b_sign1 = 4'd7; b_sign2 = 4'd9; b_sign3 = 4'd8;
@(posedge clk_i);
a_mant0 = 8'd227; a_mant1 = 8'd149; a_mant2 = 8'd195; a_mant3 = 8'd222;
b_mant0 = 8'd64; b_mant1 = 8'd183; b_mant2 = 8'd109; b_mant3 = 8'd134;
a_exp0 = 10'd843; a_exp1 = 10'd436; a_exp2 = 10'd297; a_exp3 = 10'd658;
b_exp0 = 10'd1005; b_exp1 = 10'd918; b_exp2 = 10'd387; b_exp3 = 10'd346;
a_sign0 = 4'd14; a_sign1 = 4'd12; a_sign2 = 4'd5; a_sign3 = 4'd15;
b_sign0 = 4'd1; b_sign1 = 4'd8; b_sign2 = 4'd14; b_sign3 = 4'd10;
@(posedge clk_i);
a_mant0 = 8'd133; a_mant1 = 8'd181; a_mant2 = 8'd227; a_mant3 = 8'd153;
b_mant0 = 8'd192; b_mant1 = 8'd139; b_mant2 = 8'd236; b_mant3 = 8'd117;
a_exp0 = 10'd884; a_exp1 = 10'd57; a_exp2 = 10'd789; a_exp3 = 10'd1004;
b_exp0 = 10'd129; b_exp1 = 10'd811; b_exp2 = 10'd201; b_exp3 = 10'd1;
a_sign0 = 4'd7; a_sign1 = 4'd1; a_sign2 = 4'd2; a_sign3 = 4'd9;
b_sign0 = 4'd1; b_sign1 = 4'd7; b_sign2 = 4'd10; b_sign3 = 4'd10;
@(posedge clk_i);
a_mant0 = 8'd18; a_mant1 = 8'd23; a_mant2 = 8'd34; a_mant3 = 8'd22;
b_mant0 = 8'd79; b_mant1 = 8'd247; b_mant2 = 8'd142; b_mant3 = 8'd95;
a_exp0 = 10'd888; a_exp1 = 10'd311; a_exp2 = 10'd801; a_exp3 = 10'd199;
b_exp0 = 10'd704; b_exp1 = 10'd810; b_exp2 = 10'd687; b_exp3 = 10'd835;
a_sign0 = 4'd7; a_sign1 = 4'd16; a_sign2 = 4'd7; a_sign3 = 4'd6;
b_sign0 = 4'd6; b_sign1 = 4'd15; b_sign2 = 4'd3; b_sign3 = 4'd1;
@(posedge clk_i);
a_mant0 = 8'd239; a_mant1 = 8'd67; a_mant2 = 8'd190; a_mant3 = 8'd48;
b_mant0 = 8'd226; b_mant1 = 8'd121; b_mant2 = 8'd103; b_mant3 = 8'd27;
a_exp0 = 10'd455; a_exp1 = 10'd944; a_exp2 = 10'd259; a_exp3 = 10'd700;
b_exp0 = 10'd328; b_exp1 = 10'd607; b_exp2 = 10'd887; b_exp3 = 10'd581;
a_sign0 = 4'd3; a_sign1 = 4'd9; a_sign2 = 4'd0; a_sign3 = 4'd9;
b_sign0 = 4'd1; b_sign1 = 4'd11; b_sign2 = 4'd3; b_sign3 = 4'd0;
@(posedge clk_i);
a_mant0 = 8'd212; a_mant1 = 8'd186; a_mant2 = 8'd48; a_mant3 = 8'd51;
b_mant0 = 8'd170; b_mant1 = 8'd212; b_mant2 = 8'd253; b_mant3 = 8'd249;
a_exp0 = 10'd358; a_exp1 = 10'd271; a_exp2 = 10'd965; a_exp3 = 10'd37;
b_exp0 = 10'd583; b_exp1 = 10'd1016; b_exp2 = 10'd895; b_exp3 = 10'd405;
a_sign0 = 4'd12; a_sign1 = 4'd8; a_sign2 = 4'd13; a_sign3 = 4'd1;
b_sign0 = 4'd4; b_sign1 = 4'd5; b_sign2 = 4'd8; b_sign3 = 4'd12;
@(posedge clk_i);
shared_exps0 = 8'd103;
shared_exps1 = 8'd134;
a_mant0 = 8'd7; a_mant1 = 8'd117; a_mant2 = 8'd138; a_mant3 = 8'd61;
b_mant0 = 8'd165; b_mant1 = 8'd13; b_mant2 = 8'd172; b_mant3 = 8'd172;
a_exp0 = 10'd52; a_exp1 = 10'd63; a_exp2 = 10'd251; a_exp3 = 10'd554;
b_exp0 = 10'd886; b_exp1 = 10'd112; b_exp2 = 10'd985; b_exp3 = 10'd529;
a_sign0 = 4'd13; a_sign1 = 4'd15; a_sign2 = 4'd3; a_sign3 = 4'd11;
b_sign0 = 4'd12; b_sign1 = 4'd14; b_sign2 = 4'd7; b_sign3 = 4'd5;
@(posedge clk_i);
a_mant0 = 8'd21; a_mant1 = 8'd155; a_mant2 = 8'd6; a_mant3 = 8'd31;
b_mant0 = 8'd102; b_mant1 = 8'd191; b_mant2 = 8'd64; b_mant3 = 8'd29;
a_exp0 = 10'd683; a_exp1 = 10'd413; a_exp2 = 10'd789; a_exp3 = 10'd684;
b_exp0 = 10'd409; b_exp1 = 10'd599; b_exp2 = 10'd450; b_exp3 = 10'd926;
a_sign0 = 4'd2; a_sign1 = 4'd11; a_sign2 = 4'd10; a_sign3 = 4'd3;
b_sign0 = 4'd12; b_sign1 = 4'd10; b_sign2 = 4'd8; b_sign3 = 4'd9;
@(posedge clk_i);
a_mant0 = 8'd153; a_mant1 = 8'd151; a_mant2 = 8'd231; a_mant3 = 8'd206;
b_mant0 = 8'd34; b_mant1 = 8'd143; b_mant2 = 8'd52; b_mant3 = 8'd111;
a_exp0 = 10'd419; a_exp1 = 10'd997; a_exp2 = 10'd660; a_exp3 = 10'd748;
b_exp0 = 10'd58; b_exp1 = 10'd839; b_exp2 = 10'd247; b_exp3 = 10'd291;
a_sign0 = 4'd9; a_sign1 = 4'd16; a_sign2 = 4'd4; a_sign3 = 4'd2;
b_sign0 = 4'd0; b_sign1 = 4'd15; b_sign2 = 4'd7; b_sign3 = 4'd6;
@(posedge clk_i);
a_mant0 = 8'd180; a_mant1 = 8'd82; a_mant2 = 8'd100; a_mant3 = 8'd158;
b_mant0 = 8'd241; b_mant1 = 8'd56; b_mant2 = 8'd24; b_mant3 = 8'd208;
a_exp0 = 10'd155; a_exp1 = 10'd780; a_exp2 = 10'd896; a_exp3 = 10'd987;
b_exp0 = 10'd397; b_exp1 = 10'd326; b_exp2 = 10'd664; b_exp3 = 10'd302;
a_sign0 = 4'd8; a_sign1 = 4'd15; a_sign2 = 4'd13; a_sign3 = 4'd16;
b_sign0 = 4'd10; b_sign1 = 4'd14; b_sign2 = 4'd7; b_sign3 = 4'd1;
@(posedge clk_i);
a_mant0 = 8'd157; a_mant1 = 8'd253; a_mant2 = 8'd75; a_mant3 = 8'd168;
b_mant0 = 8'd206; b_mant1 = 8'd30; b_mant2 = 8'd144; b_mant3 = 8'd147;
a_exp0 = 10'd871; a_exp1 = 10'd329; a_exp2 = 10'd874; a_exp3 = 10'd954;
b_exp0 = 10'd795; b_exp1 = 10'd30; b_exp2 = 10'd879; b_exp3 = 10'd325;
a_sign0 = 4'd8; a_sign1 = 4'd5; a_sign2 = 4'd2; a_sign3 = 4'd0;
b_sign0 = 4'd3; b_sign1 = 4'd5; b_sign2 = 4'd1; b_sign3 = 4'd1;
@(posedge clk_i);
a_mant0 = 8'd180; a_mant1 = 8'd76; a_mant2 = 8'd21; a_mant3 = 8'd188;
b_mant0 = 8'd160; b_mant1 = 8'd249; b_mant2 = 8'd158; b_mant3 = 8'd143;
a_exp0 = 10'd830; a_exp1 = 10'd898; a_exp2 = 10'd601; a_exp3 = 10'd256;
b_exp0 = 10'd298; b_exp1 = 10'd4; b_exp2 = 10'd151; b_exp3 = 10'd970;
a_sign0 = 4'd6; a_sign1 = 4'd9; a_sign2 = 4'd2; a_sign3 = 4'd15;
b_sign0 = 4'd7; b_sign1 = 4'd12; b_sign2 = 4'd11; b_sign3 = 4'd1;
@(posedge clk_i);
a_mant0 = 8'd242; a_mant1 = 8'd51; a_mant2 = 8'd200; a_mant3 = 8'd122;
b_mant0 = 8'd85; b_mant1 = 8'd50; b_mant2 = 8'd11; b_mant3 = 8'd65;
a_exp0 = 10'd122; a_exp1 = 10'd291; a_exp2 = 10'd5; a_exp3 = 10'd675;
b_exp0 = 10'd593; b_exp1 = 10'd709; b_exp2 = 10'd108; b_exp3 = 10'd980;
a_sign0 = 4'd14; a_sign1 = 4'd1; a_sign2 = 4'd7; a_sign3 = 4'd2;
b_sign0 = 4'd11; b_sign1 = 4'd3; b_sign2 = 4'd1; b_sign3 = 4'd7;
@(posedge clk_i);
a_mant0 = 8'd87; a_mant1 = 8'd198; a_mant2 = 8'd172; a_mant3 = 8'd44;
b_mant0 = 8'd13; b_mant1 = 8'd153; b_mant2 = 8'd48; b_mant3 = 8'd29;
a_exp0 = 10'd462; a_exp1 = 10'd816; a_exp2 = 10'd78; a_exp3 = 10'd546;
b_exp0 = 10'd932; b_exp1 = 10'd925; b_exp2 = 10'd741; b_exp3 = 10'd688;
a_sign0 = 4'd1; a_sign1 = 4'd13; a_sign2 = 4'd0; a_sign3 = 4'd3;
b_sign0 = 4'd7; b_sign1 = 4'd16; b_sign2 = 4'd2; b_sign3 = 4'd13;
@(posedge clk_i);
shared_exps0 = 8'd93;
shared_exps1 = 8'd160;
rstn = 0;
@(posedge clk_i);
rstn = 1;
a_mant0 = 8'd100; a_mant1 = 8'd215; a_mant2 = 8'd233; a_mant3 = 8'd189;
b_mant0 = 8'd183; b_mant1 = 8'd251; b_mant2 = 8'd133; b_mant3 = 8'd171;
a_exp0 = 10'd650; a_exp1 = 10'd557; a_exp2 = 10'd959; a_exp3 = 10'd885;
b_exp0 = 10'd642; b_exp1 = 10'd200; b_exp2 = 10'd321; b_exp3 = 10'd599;
a_sign0 = 4'd1; a_sign1 = 4'd8; a_sign2 = 4'd6; a_sign3 = 4'd3;
b_sign0 = 4'd3; b_sign1 = 4'd2; b_sign2 = 4'd4; b_sign3 = 4'd11;
@(posedge clk_i);
a_mant0 = 8'd193; a_mant1 = 8'd12; a_mant2 = 8'd2; a_mant3 = 8'd206;
b_mant0 = 8'd26; b_mant1 = 8'd73; b_mant2 = 8'd254; b_mant3 = 8'd250;
a_exp0 = 10'd988; a_exp1 = 10'd422; a_exp2 = 10'd354; a_exp3 = 10'd981;
b_exp0 = 10'd14; b_exp1 = 10'd898; b_exp2 = 10'd902; b_exp3 = 10'd994;
a_sign0 = 4'd16; a_sign1 = 4'd13; a_sign2 = 4'd12; a_sign3 = 4'd3;
b_sign0 = 4'd15; b_sign1 = 4'd13; b_sign2 = 4'd2; b_sign3 = 4'd16;
@(posedge clk_i);
a_mant0 = 8'd234; a_mant1 = 8'd89; a_mant2 = 8'd228; a_mant3 = 8'd68;
b_mant0 = 8'd227; b_mant1 = 8'd194; b_mant2 = 8'd6; b_mant3 = 8'd7;
a_exp0 = 10'd355; a_exp1 = 10'd439; a_exp2 = 10'd268; a_exp3 = 10'd550;
b_exp0 = 10'd1008; b_exp1 = 10'd502; b_exp2 = 10'd777; b_exp3 = 10'd492;
a_sign0 = 4'd10; a_sign1 = 4'd8; a_sign2 = 4'd6; a_sign3 = 4'd14;
b_sign0 = 4'd16; b_sign1 = 4'd13; b_sign2 = 4'd1; b_sign3 = 4'd12;
@(posedge clk_i);
a_mant0 = 8'd138; a_mant1 = 8'd151; a_mant2 = 8'd236; a_mant3 = 8'd41;
b_mant0 = 8'd166; b_mant1 = 8'd179; b_mant2 = 8'd37; b_mant3 = 8'd17;
a_exp0 = 10'd728; a_exp1 = 10'd492; a_exp2 = 10'd965; a_exp3 = 10'd784;
b_exp0 = 10'd732; b_exp1 = 10'd177; b_exp2 = 10'd675; b_exp3 = 10'd68;
a_sign0 = 4'd14; a_sign1 = 4'd9; a_sign2 = 4'd13; a_sign3 = 4'd16;
b_sign0 = 4'd15; b_sign1 = 4'd8; b_sign2 = 4'd16; b_sign3 = 4'd3;
@(posedge clk_i);
a_mant0 = 8'd76; a_mant1 = 8'd159; a_mant2 = 8'd114; a_mant3 = 8'd117;
b_mant0 = 8'd96; b_mant1 = 8'd75; b_mant2 = 8'd51; b_mant3 = 8'd150;
a_exp0 = 10'd280; a_exp1 = 10'd926; a_exp2 = 10'd80; a_exp3 = 10'd589;
b_exp0 = 10'd946; b_exp1 = 10'd877; b_exp2 = 10'd323; b_exp3 = 10'd530;
a_sign0 = 4'd0; a_sign1 = 4'd4; a_sign2 = 4'd14; a_sign3 = 4'd13;
b_sign0 = 4'd13; b_sign1 = 4'd5; b_sign2 = 4'd1; b_sign3 = 4'd14;
@(posedge clk_i);
a_mant0 = 8'd123; a_mant1 = 8'd77; a_mant2 = 8'd79; a_mant3 = 8'd45;
b_mant0 = 8'd112; b_mant1 = 8'd113; b_mant2 = 8'd193; b_mant3 = 8'd190;
a_exp0 = 10'd60; a_exp1 = 10'd965; a_exp2 = 10'd335; a_exp3 = 10'd255;
b_exp0 = 10'd238; b_exp1 = 10'd817; b_exp2 = 10'd310; b_exp3 = 10'd34;
a_sign0 = 4'd15; a_sign1 = 4'd12; a_sign2 = 4'd0; a_sign3 = 4'd11;
b_sign0 = 4'd9; b_sign1 = 4'd0; b_sign2 = 4'd16; b_sign3 = 4'd13;
@(posedge clk_i);
a_mant0 = 8'd4; a_mant1 = 8'd246; a_mant2 = 8'd60; a_mant3 = 8'd212;
b_mant0 = 8'd26; b_mant1 = 8'd46; b_mant2 = 8'd186; b_mant3 = 8'd126;
a_exp0 = 10'd801; a_exp1 = 10'd697; a_exp2 = 10'd641; a_exp3 = 10'd538;
b_exp0 = 10'd1019; b_exp1 = 10'd6; b_exp2 = 10'd921; b_exp3 = 10'd698;
a_sign0 = 4'd9; a_sign1 = 4'd10; a_sign2 = 4'd8; a_sign3 = 4'd15;
b_sign0 = 4'd14; b_sign1 = 4'd12; b_sign2 = 4'd6; b_sign3 = 4'd7;
@(posedge clk_i);
shared_exps0 = 8'd123;
shared_exps1 = 8'd125;
a_mant0 = 8'd116; a_mant1 = 8'd222; a_mant2 = 8'd72; a_mant3 = 8'd203;
b_mant0 = 8'd119; b_mant1 = 8'd1; b_mant2 = 8'd156; b_mant3 = 8'd48;
a_exp0 = 10'd990; a_exp1 = 10'd661; a_exp2 = 10'd358; a_exp3 = 10'd804;
b_exp0 = 10'd946; b_exp1 = 10'd465; b_exp2 = 10'd60; b_exp3 = 10'd44;
a_sign0 = 4'd13; a_sign1 = 4'd15; a_sign2 = 4'd12; a_sign3 = 4'd1;
b_sign0 = 4'd6; b_sign1 = 4'd8; b_sign2 = 4'd14; b_sign3 = 4'd9;
@(posedge clk_i);
a_mant0 = 8'd113; a_mant1 = 8'd226; a_mant2 = 8'd43; a_mant3 = 8'd23;
b_mant0 = 8'd160; b_mant1 = 8'd72; b_mant2 = 8'd120; b_mant3 = 8'd97;
a_exp0 = 10'd557; a_exp1 = 10'd664; a_exp2 = 10'd748; a_exp3 = 10'd489;
b_exp0 = 10'd806; b_exp1 = 10'd260; b_exp2 = 10'd494; b_exp3 = 10'd849;
a_sign0 = 4'd10; a_sign1 = 4'd12; a_sign2 = 4'd10; a_sign3 = 4'd13;
b_sign0 = 4'd16; b_sign1 = 4'd16; b_sign2 = 4'd11; b_sign3 = 4'd5;
@(posedge clk_i);
a_mant0 = 8'd63; a_mant1 = 8'd63; a_mant2 = 8'd120; a_mant3 = 8'd130;
b_mant0 = 8'd228; b_mant1 = 8'd103; b_mant2 = 8'd196; b_mant3 = 8'd105;
a_exp0 = 10'd489; a_exp1 = 10'd113; a_exp2 = 10'd725; a_exp3 = 10'd47;
b_exp0 = 10'd834; b_exp1 = 10'd179; b_exp2 = 10'd168; b_exp3 = 10'd368;
a_sign0 = 4'd6; a_sign1 = 4'd4; a_sign2 = 4'd9; a_sign3 = 4'd15;
b_sign0 = 4'd5; b_sign1 = 4'd5; b_sign2 = 4'd12; b_sign3 = 4'd7;
@(posedge clk_i);
a_mant0 = 8'd220; a_mant1 = 8'd67; a_mant2 = 8'd152; a_mant3 = 8'd221;
b_mant0 = 8'd1; b_mant1 = 8'd17; b_mant2 = 8'd24; b_mant3 = 8'd86;
a_exp0 = 10'd1; a_exp1 = 10'd795; a_exp2 = 10'd997; a_exp3 = 10'd978;
b_exp0 = 10'd871; b_exp1 = 10'd393; b_exp2 = 10'd702; b_exp3 = 10'd590;
a_sign0 = 4'd7; a_sign1 = 4'd11; a_sign2 = 4'd5; a_sign3 = 4'd10;
b_sign0 = 4'd7; b_sign1 = 4'd9; b_sign2 = 4'd7; b_sign3 = 4'd5;
@(posedge clk_i);
a_mant0 = 8'd245; a_mant1 = 8'd247; a_mant2 = 8'd111; a_mant3 = 8'd3;
b_mant0 = 8'd229; b_mant1 = 8'd188; b_mant2 = 8'd243; b_mant3 = 8'd215;
a_exp0 = 10'd813; a_exp1 = 10'd414; a_exp2 = 10'd798; a_exp3 = 10'd788;
b_exp0 = 10'd909; b_exp1 = 10'd209; b_exp2 = 10'd874; b_exp3 = 10'd943;
a_sign0 = 4'd8; a_sign1 = 4'd10; a_sign2 = 4'd15; a_sign3 = 4'd12;
b_sign0 = 4'd2; b_sign1 = 4'd12; b_sign2 = 4'd8; b_sign3 = 4'd0;
@(posedge clk_i);
a_mant0 = 8'd4; a_mant1 = 8'd119; a_mant2 = 8'd174; a_mant3 = 8'd102;
b_mant0 = 8'd80; b_mant1 = 8'd23; b_mant2 = 8'd73; b_mant3 = 8'd149;
a_exp0 = 10'd818; a_exp1 = 10'd703; a_exp2 = 10'd2; a_exp3 = 10'd116;
b_exp0 = 10'd407; b_exp1 = 10'd908; b_exp2 = 10'd885; b_exp3 = 10'd116;
a_sign0 = 4'd6; a_sign1 = 4'd8; a_sign2 = 4'd11; a_sign3 = 4'd9;
b_sign0 = 4'd1; b_sign1 = 4'd4; b_sign2 = 4'd2; b_sign3 = 4'd11;
@(posedge clk_i);
a_mant0 = 8'd223; a_mant1 = 8'd138; a_mant2 = 8'd213; a_mant3 = 8'd143;
b_mant0 = 8'd76; b_mant1 = 8'd38; b_mant2 = 8'd145; b_mant3 = 8'd21;
a_exp0 = 10'd167; a_exp1 = 10'd812; a_exp2 = 10'd567; a_exp3 = 10'd713;
b_exp0 = 10'd315; b_exp1 = 10'd207; b_exp2 = 10'd307; b_exp3 = 10'd794;
a_sign0 = 4'd0; a_sign1 = 4'd4; a_sign2 = 4'd6; a_sign3 = 4'd10;
b_sign0 = 4'd0; b_sign1 = 4'd16; b_sign2 = 4'd16; b_sign3 = 4'd10;
@(posedge clk_i);
a_mant0 = 8'd166; a_mant1 = 8'd241; a_mant2 = 8'd5; a_mant3 = 8'd26;
b_mant0 = 8'd80; b_mant1 = 8'd155; b_mant2 = 8'd136; b_mant3 = 8'd170;
a_exp0 = 10'd620; a_exp1 = 10'd785; a_exp2 = 10'd860; a_exp3 = 10'd846;
b_exp0 = 10'd810; b_exp1 = 10'd274; b_exp2 = 10'd874; b_exp3 = 10'd817;
a_sign0 = 4'd5; a_sign1 = 4'd15; a_sign2 = 4'd8; a_sign3 = 4'd0;
b_sign0 = 4'd0; b_sign1 = 4'd12; b_sign2 = 4'd7; b_sign3 = 4'd9;
@(posedge clk_i);
shared_exps0 = 8'd142;
shared_exps1 = 8'd115;
a_mant0 = 8'd38; a_mant1 = 8'd155; a_mant2 = 8'd52; a_mant3 = 8'd135;
b_mant0 = 8'd229; b_mant1 = 8'd105; b_mant2 = 8'd108; b_mant3 = 8'd76;
a_exp0 = 10'd163; a_exp1 = 10'd819; a_exp2 = 10'd211; a_exp3 = 10'd357;
b_exp0 = 10'd869; b_exp1 = 10'd688; b_exp2 = 10'd627; b_exp3 = 10'd326;
a_sign0 = 4'd11; a_sign1 = 4'd4; a_sign2 = 4'd16; a_sign3 = 4'd7;
b_sign0 = 4'd13; b_sign1 = 4'd5; b_sign2 = 4'd12; b_sign3 = 4'd11;
@(posedge clk_i);
a_mant0 = 8'd112; a_mant1 = 8'd69; a_mant2 = 8'd72; a_mant3 = 8'd97;
b_mant0 = 8'd98; b_mant1 = 8'd191; b_mant2 = 8'd2; b_mant3 = 8'd180;
a_exp0 = 10'd32; a_exp1 = 10'd930; a_exp2 = 10'd735; a_exp3 = 10'd598;
b_exp0 = 10'd216; b_exp1 = 10'd78; b_exp2 = 10'd254; b_exp3 = 10'd389;
a_sign0 = 4'd14; a_sign1 = 4'd9; a_sign2 = 4'd16; a_sign3 = 4'd13;
b_sign0 = 4'd13; b_sign1 = 4'd5; b_sign2 = 4'd6; b_sign3 = 4'd7;
@(posedge clk_i);
a_mant0 = 8'd44; a_mant1 = 8'd74; a_mant2 = 8'd11; a_mant3 = 8'd232;
b_mant0 = 8'd53; b_mant1 = 8'd133; b_mant2 = 8'd0; b_mant3 = 8'd251;
a_exp0 = 10'd222; a_exp1 = 10'd693; a_exp2 = 10'd467; a_exp3 = 10'd912;
b_exp0 = 10'd651; b_exp1 = 10'd912; b_exp2 = 10'd553; b_exp3 = 10'd540;
a_sign0 = 4'd5; a_sign1 = 4'd15; a_sign2 = 4'd7; a_sign3 = 4'd12;
b_sign0 = 4'd11; b_sign1 = 4'd0; b_sign2 = 4'd3; b_sign3 = 4'd4;
@(posedge clk_i);
a_mant0 = 8'd82; a_mant1 = 8'd147; a_mant2 = 8'd22; a_mant3 = 8'd86;
b_mant0 = 8'd153; b_mant1 = 8'd75; b_mant2 = 8'd57; b_mant3 = 8'd22;
a_exp0 = 10'd246; a_exp1 = 10'd326; a_exp2 = 10'd265; a_exp3 = 10'd914;
b_exp0 = 10'd23; b_exp1 = 10'd156; b_exp2 = 10'd574; b_exp3 = 10'd37;
a_sign0 = 4'd15; a_sign1 = 4'd8; a_sign2 = 4'd2; a_sign3 = 4'd15;
b_sign0 = 4'd16; b_sign1 = 4'd16; b_sign2 = 4'd0; b_sign3 = 4'd6;
@(posedge clk_i);
a_mant0 = 8'd191; a_mant1 = 8'd167; a_mant2 = 8'd41; a_mant3 = 8'd159;
b_mant0 = 8'd190; b_mant1 = 8'd245; b_mant2 = 8'd51; b_mant3 = 8'd140;
a_exp0 = 10'd246; a_exp1 = 10'd201; a_exp2 = 10'd732; a_exp3 = 10'd64;
b_exp0 = 10'd547; b_exp1 = 10'd13; b_exp2 = 10'd653; b_exp3 = 10'd742;
a_sign0 = 4'd14; a_sign1 = 4'd4; a_sign2 = 4'd9; a_sign3 = 4'd11;
b_sign0 = 4'd3; b_sign1 = 4'd0; b_sign2 = 4'd9; b_sign3 = 4'd12;
@(posedge clk_i);
a_mant0 = 8'd143; a_mant1 = 8'd104; a_mant2 = 8'd131; a_mant3 = 8'd188;
b_mant0 = 8'd164; b_mant1 = 8'd67; b_mant2 = 8'd201; b_mant3 = 8'd63;
a_exp0 = 10'd455; a_exp1 = 10'd686; a_exp2 = 10'd322; a_exp3 = 10'd663;
b_exp0 = 10'd111; b_exp1 = 10'd136; b_exp2 = 10'd551; b_exp3 = 10'd992;
a_sign0 = 4'd2; a_sign1 = 4'd7; a_sign2 = 4'd13; a_sign3 = 4'd1;
b_sign0 = 4'd14; b_sign1 = 4'd5; b_sign2 = 4'd6; b_sign3 = 4'd7;
@(posedge clk_i);
a_mant0 = 8'd46; a_mant1 = 8'd124; a_mant2 = 8'd62; a_mant3 = 8'd63;
b_mant0 = 8'd78; b_mant1 = 8'd123; b_mant2 = 8'd163; b_mant3 = 8'd144;
a_exp0 = 10'd199; a_exp1 = 10'd983; a_exp2 = 10'd225; a_exp3 = 10'd638;
b_exp0 = 10'd947; b_exp1 = 10'd695; b_exp2 = 10'd273; b_exp3 = 10'd101;
a_sign0 = 4'd10; a_sign1 = 4'd12; a_sign2 = 4'd10; a_sign3 = 4'd2;
b_sign0 = 4'd1; b_sign1 = 4'd4; b_sign2 = 4'd3; b_sign3 = 4'd8;
@(posedge clk_i);
a_mant0 = 8'd112; a_mant1 = 8'd35; a_mant2 = 8'd222; a_mant3 = 8'd92;
b_mant0 = 8'd38; b_mant1 = 8'd119; b_mant2 = 8'd135; b_mant3 = 8'd182;
a_exp0 = 10'd315; a_exp1 = 10'd539; a_exp2 = 10'd869; a_exp3 = 10'd963;
b_exp0 = 10'd506; b_exp1 = 10'd358; b_exp2 = 10'd487; b_exp3 = 10'd764;
a_sign0 = 4'd9; a_sign1 = 4'd2; a_sign2 = 4'd14; a_sign3 = 4'd1;
b_sign0 = 4'd15; b_sign1 = 4'd1; b_sign2 = 4'd2; b_sign3 = 4'd14;
@(posedge clk_i);
shared_exps0 = 8'd131;
shared_exps1 = 8'd129;
a_mant0 = 8'd101; a_mant1 = 8'd173; a_mant2 = 8'd197; a_mant3 = 8'd171;
b_mant0 = 8'd52; b_mant1 = 8'd183; b_mant2 = 8'd254; b_mant3 = 8'd145;
a_exp0 = 10'd582; a_exp1 = 10'd1001; a_exp2 = 10'd864; a_exp3 = 10'd791;
b_exp0 = 10'd701; b_exp1 = 10'd412; b_exp2 = 10'd882; b_exp3 = 10'd439;
a_sign0 = 4'd6; a_sign1 = 4'd16; a_sign2 = 4'd10; a_sign3 = 4'd8;
b_sign0 = 4'd8; b_sign1 = 4'd0; b_sign2 = 4'd7; b_sign3 = 4'd2;
@(posedge clk_i);
a_mant0 = 8'd32; a_mant1 = 8'd51; a_mant2 = 8'd21; a_mant3 = 8'd99;
b_mant0 = 8'd78; b_mant1 = 8'd20; b_mant2 = 8'd26; b_mant3 = 8'd215;
a_exp0 = 10'd754; a_exp1 = 10'd567; a_exp2 = 10'd692; a_exp3 = 10'd998;
b_exp0 = 10'd509; b_exp1 = 10'd389; b_exp2 = 10'd680; b_exp3 = 10'd344;
a_sign0 = 4'd8; a_sign1 = 4'd1; a_sign2 = 4'd4; a_sign3 = 4'd16;
b_sign0 = 4'd2; b_sign1 = 4'd7; b_sign2 = 4'd0; b_sign3 = 4'd16;
@(posedge clk_i);
a_mant0 = 8'd150; a_mant1 = 8'd112; a_mant2 = 8'd201; a_mant3 = 8'd251;
b_mant0 = 8'd37; b_mant1 = 8'd63; b_mant2 = 8'd208; b_mant3 = 8'd52;
a_exp0 = 10'd981; a_exp1 = 10'd273; a_exp2 = 10'd592; a_exp3 = 10'd497;
b_exp0 = 10'd603; b_exp1 = 10'd447; b_exp2 = 10'd1017; b_exp3 = 10'd418;
a_sign0 = 4'd3; a_sign1 = 4'd16; a_sign2 = 4'd9; a_sign3 = 4'd14;
b_sign0 = 4'd0; b_sign1 = 4'd14; b_sign2 = 4'd0; b_sign3 = 4'd12;
@(posedge clk_i);
a_mant0 = 8'd149; a_mant1 = 8'd10; a_mant2 = 8'd116; a_mant3 = 8'd117;
b_mant0 = 8'd111; b_mant1 = 8'd233; b_mant2 = 8'd159; b_mant3 = 8'd97;
a_exp0 = 10'd415; a_exp1 = 10'd679; a_exp2 = 10'd552; a_exp3 = 10'd750;
b_exp0 = 10'd458; b_exp1 = 10'd596; b_exp2 = 10'd623; b_exp3 = 10'd0;
a_sign0 = 4'd14; a_sign1 = 4'd8; a_sign2 = 4'd6; a_sign3 = 4'd9;
b_sign0 = 4'd15; b_sign1 = 4'd14; b_sign2 = 4'd4; b_sign3 = 4'd16;
@(posedge clk_i);
a_mant0 = 8'd191; a_mant1 = 8'd205; a_mant2 = 8'd176; a_mant3 = 8'd102;
b_mant0 = 8'd254; b_mant1 = 8'd67; b_mant2 = 8'd191; b_mant3 = 8'd249;
a_exp0 = 10'd938; a_exp1 = 10'd239; a_exp2 = 10'd420; a_exp3 = 10'd921;
b_exp0 = 10'd1002; b_exp1 = 10'd758; b_exp2 = 10'd231; b_exp3 = 10'd399;
a_sign0 = 4'd4; a_sign1 = 4'd15; a_sign2 = 4'd4; a_sign3 = 4'd7;
b_sign0 = 4'd16; b_sign1 = 4'd13; b_sign2 = 4'd15; b_sign3 = 4'd8;
@(posedge clk_i);
a_mant0 = 8'd196; a_mant1 = 8'd172; a_mant2 = 8'd250; a_mant3 = 8'd93;
b_mant0 = 8'd67; b_mant1 = 8'd229; b_mant2 = 8'd232; b_mant3 = 8'd210;
a_exp0 = 10'd184; a_exp1 = 10'd572; a_exp2 = 10'd544; a_exp3 = 10'd237;
b_exp0 = 10'd556; b_exp1 = 10'd775; b_exp2 = 10'd628; b_exp3 = 10'd387;
a_sign0 = 4'd16; a_sign1 = 4'd15; a_sign2 = 4'd13; a_sign3 = 4'd15;
b_sign0 = 4'd13; b_sign1 = 4'd9; b_sign2 = 4'd6; b_sign3 = 4'd15;
@(posedge clk_i);
a_mant0 = 8'd137; a_mant1 = 8'd107; a_mant2 = 8'd133; a_mant3 = 8'd237;
b_mant0 = 8'd244; b_mant1 = 8'd7; b_mant2 = 8'd207; b_mant3 = 8'd28;
a_exp0 = 10'd797; a_exp1 = 10'd185; a_exp2 = 10'd279; a_exp3 = 10'd130;
b_exp0 = 10'd436; b_exp1 = 10'd1009; b_exp2 = 10'd397; b_exp3 = 10'd172;
a_sign0 = 4'd1; a_sign1 = 4'd10; a_sign2 = 4'd5; a_sign3 = 4'd11;
b_sign0 = 4'd1; b_sign1 = 4'd0; b_sign2 = 4'd13; b_sign3 = 4'd12;
@(posedge clk_i);
a_mant0 = 8'd33; a_mant1 = 8'd92; a_mant2 = 8'd15; a_mant3 = 8'd245;
b_mant0 = 8'd252; b_mant1 = 8'd104; b_mant2 = 8'd222; b_mant3 = 8'd12;
a_exp0 = 10'd494; a_exp1 = 10'd947; a_exp2 = 10'd885; a_exp3 = 10'd996;
b_exp0 = 10'd341; b_exp1 = 10'd70; b_exp2 = 10'd192; b_exp3 = 10'd740;
a_sign0 = 4'd4; a_sign1 = 4'd7; a_sign2 = 4'd16; a_sign3 = 4'd1;
b_sign0 = 4'd8; b_sign1 = 4'd0; b_sign2 = 4'd10; b_sign3 = 4'd14;
@(posedge clk_i);
shared_exps0 = 8'd125;
shared_exps1 = 8'd131;
rstn = 0;
@(posedge clk_i);
rstn = 1;
a_mant0 = 8'd61; a_mant1 = 8'd4; a_mant2 = 8'd63; a_mant3 = 8'd65;
b_mant0 = 8'd109; b_mant1 = 8'd231; b_mant2 = 8'd43; b_mant3 = 8'd157;
a_exp0 = 10'd366; a_exp1 = 10'd391; a_exp2 = 10'd28; a_exp3 = 10'd955;
b_exp0 = 10'd179; b_exp1 = 10'd446; b_exp2 = 10'd88; b_exp3 = 10'd410;
a_sign0 = 4'd6; a_sign1 = 4'd4; a_sign2 = 4'd6; a_sign3 = 4'd8;
b_sign0 = 4'd14; b_sign1 = 4'd3; b_sign2 = 4'd5; b_sign3 = 4'd5;
@(posedge clk_i);
a_mant0 = 8'd208; a_mant1 = 8'd98; a_mant2 = 8'd203; a_mant3 = 8'd65;
b_mant0 = 8'd52; b_mant1 = 8'd228; b_mant2 = 8'd73; b_mant3 = 8'd110;
a_exp0 = 10'd912; a_exp1 = 10'd492; a_exp2 = 10'd866; a_exp3 = 10'd169;
b_exp0 = 10'd781; b_exp1 = 10'd62; b_exp2 = 10'd208; b_exp3 = 10'd927;
a_sign0 = 4'd7; a_sign1 = 4'd11; a_sign2 = 4'd9; a_sign3 = 4'd16;
b_sign0 = 4'd3; b_sign1 = 4'd8; b_sign2 = 4'd1; b_sign3 = 4'd8;
@(posedge clk_i);
a_mant0 = 8'd222; a_mant1 = 8'd241; a_mant2 = 8'd49; a_mant3 = 8'd103;
b_mant0 = 8'd66; b_mant1 = 8'd147; b_mant2 = 8'd240; b_mant3 = 8'd73;
a_exp0 = 10'd457; a_exp1 = 10'd234; a_exp2 = 10'd466; a_exp3 = 10'd195;
b_exp0 = 10'd265; b_exp1 = 10'd739; b_exp2 = 10'd608; b_exp3 = 10'd301;
a_sign0 = 4'd3; a_sign1 = 4'd7; a_sign2 = 4'd1; a_sign3 = 4'd10;
b_sign0 = 4'd9; b_sign1 = 4'd2; b_sign2 = 4'd3; b_sign3 = 4'd0;
@(posedge clk_i);
a_mant0 = 8'd131; a_mant1 = 8'd204; a_mant2 = 8'd44; a_mant3 = 8'd44;
b_mant0 = 8'd27; b_mant1 = 8'd3; b_mant2 = 8'd143; b_mant3 = 8'd53;
a_exp0 = 10'd311; a_exp1 = 10'd453; a_exp2 = 10'd568; a_exp3 = 10'd96;
b_exp0 = 10'd204; b_exp1 = 10'd539; b_exp2 = 10'd708; b_exp3 = 10'd1017;
a_sign0 = 4'd13; a_sign1 = 4'd6; a_sign2 = 4'd14; a_sign3 = 4'd6;
b_sign0 = 4'd0; b_sign1 = 4'd0; b_sign2 = 4'd12; b_sign3 = 4'd10;
@(posedge clk_i);
a_mant0 = 8'd8; a_mant1 = 8'd144; a_mant2 = 8'd103; a_mant3 = 8'd212;
b_mant0 = 8'd25; b_mant1 = 8'd102; b_mant2 = 8'd1; b_mant3 = 8'd242;
a_exp0 = 10'd27; a_exp1 = 10'd695; a_exp2 = 10'd353; a_exp3 = 10'd418;
b_exp0 = 10'd330; b_exp1 = 10'd636; b_exp2 = 10'd389; b_exp3 = 10'd771;
a_sign0 = 4'd6; a_sign1 = 4'd8; a_sign2 = 4'd3; a_sign3 = 4'd6;
b_sign0 = 4'd13; b_sign1 = 4'd2; b_sign2 = 4'd9; b_sign3 = 4'd0;
@(posedge clk_i);
a_mant0 = 8'd38; a_mant1 = 8'd53; a_mant2 = 8'd239; a_mant3 = 8'd166;
b_mant0 = 8'd142; b_mant1 = 8'd50; b_mant2 = 8'd43; b_mant3 = 8'd32;
a_exp0 = 10'd902; a_exp1 = 10'd809; a_exp2 = 10'd417; a_exp3 = 10'd598;
b_exp0 = 10'd923; b_exp1 = 10'd540; b_exp2 = 10'd721; b_exp3 = 10'd672;
a_sign0 = 4'd5; a_sign1 = 4'd3; a_sign2 = 4'd5; a_sign3 = 4'd10;
b_sign0 = 4'd9; b_sign1 = 4'd12; b_sign2 = 4'd9; b_sign3 = 4'd11;
@(posedge clk_i);
a_mant0 = 8'd162; a_mant1 = 8'd167; a_mant2 = 8'd45; a_mant3 = 8'd175;
b_mant0 = 8'd124; b_mant1 = 8'd141; b_mant2 = 8'd59; b_mant3 = 8'd229;
a_exp0 = 10'd731; a_exp1 = 10'd826; a_exp2 = 10'd809; a_exp3 = 10'd999;
b_exp0 = 10'd622; b_exp1 = 10'd626; b_exp2 = 10'd866; b_exp3 = 10'd283;
a_sign0 = 4'd13; a_sign1 = 4'd1; a_sign2 = 4'd2; a_sign3 = 4'd5;
b_sign0 = 4'd12; b_sign1 = 4'd6; b_sign2 = 4'd9; b_sign3 = 4'd5;
@(posedge clk_i);
shared_exps0 = 8'd149;
shared_exps1 = 8'd108;
a_mant0 = 8'd96; a_mant1 = 8'd133; a_mant2 = 8'd217; a_mant3 = 8'd232;
b_mant0 = 8'd179; b_mant1 = 8'd162; b_mant2 = 8'd21; b_mant3 = 8'd41;
a_exp0 = 10'd460; a_exp1 = 10'd1007; a_exp2 = 10'd213; a_exp3 = 10'd998;
b_exp0 = 10'd567; b_exp1 = 10'd93; b_exp2 = 10'd106; b_exp3 = 10'd151;
a_sign0 = 4'd3; a_sign1 = 4'd2; a_sign2 = 4'd6; a_sign3 = 4'd15;
b_sign0 = 4'd4; b_sign1 = 4'd10; b_sign2 = 4'd6; b_sign3 = 4'd4;
@(posedge clk_i);
a_mant0 = 8'd255; a_mant1 = 8'd146; a_mant2 = 8'd43; a_mant3 = 8'd153;
b_mant0 = 8'd100; b_mant1 = 8'd252; b_mant2 = 8'd183; b_mant3 = 8'd10;
a_exp0 = 10'd959; a_exp1 = 10'd755; a_exp2 = 10'd74; a_exp3 = 10'd196;
b_exp0 = 10'd450; b_exp1 = 10'd767; b_exp2 = 10'd214; b_exp3 = 10'd978;
a_sign0 = 4'd14; a_sign1 = 4'd11; a_sign2 = 4'd4; a_sign3 = 4'd7;
b_sign0 = 4'd5; b_sign1 = 4'd13; b_sign2 = 4'd11; b_sign3 = 4'd8;
@(posedge clk_i);
a_mant0 = 8'd16; a_mant1 = 8'd47; a_mant2 = 8'd17; a_mant3 = 8'd184;
b_mant0 = 8'd125; b_mant1 = 8'd0; b_mant2 = 8'd241; b_mant3 = 8'd125;
a_exp0 = 10'd87; a_exp1 = 10'd353; a_exp2 = 10'd735; a_exp3 = 10'd612;
b_exp0 = 10'd789; b_exp1 = 10'd682; b_exp2 = 10'd510; b_exp3 = 10'd861;
a_sign0 = 4'd7; a_sign1 = 4'd15; a_sign2 = 4'd9; a_sign3 = 4'd4;
b_sign0 = 4'd6; b_sign1 = 4'd8; b_sign2 = 4'd14; b_sign3 = 4'd14;
@(posedge clk_i);
a_mant0 = 8'd114; a_mant1 = 8'd89; a_mant2 = 8'd133; a_mant3 = 8'd175;
b_mant0 = 8'd210; b_mant1 = 8'd134; b_mant2 = 8'd152; b_mant3 = 8'd145;
a_exp0 = 10'd868; a_exp1 = 10'd748; a_exp2 = 10'd736; a_exp3 = 10'd300;
b_exp0 = 10'd933; b_exp1 = 10'd648; b_exp2 = 10'd293; b_exp3 = 10'd919;
a_sign0 = 4'd10; a_sign1 = 4'd9; a_sign2 = 4'd6; a_sign3 = 4'd9;
b_sign0 = 4'd7; b_sign1 = 4'd9; b_sign2 = 4'd15; b_sign3 = 4'd12;
@(posedge clk_i);
a_mant0 = 8'd128; a_mant1 = 8'd27; a_mant2 = 8'd76; a_mant3 = 8'd35;
b_mant0 = 8'd122; b_mant1 = 8'd73; b_mant2 = 8'd58; b_mant3 = 8'd127;
a_exp0 = 10'd333; a_exp1 = 10'd740; a_exp2 = 10'd233; a_exp3 = 10'd210;
b_exp0 = 10'd462; b_exp1 = 10'd57; b_exp2 = 10'd988; b_exp3 = 10'd459;
a_sign0 = 4'd7; a_sign1 = 4'd11; a_sign2 = 4'd12; a_sign3 = 4'd1;
b_sign0 = 4'd15; b_sign1 = 4'd14; b_sign2 = 4'd5; b_sign3 = 4'd2;
@(posedge clk_i);
a_mant0 = 8'd32; a_mant1 = 8'd153; a_mant2 = 8'd147; a_mant3 = 8'd159;
b_mant0 = 8'd104; b_mant1 = 8'd116; b_mant2 = 8'd64; b_mant3 = 8'd2;
a_exp0 = 10'd754; a_exp1 = 10'd727; a_exp2 = 10'd880; a_exp3 = 10'd474;
b_exp0 = 10'd386; b_exp1 = 10'd302; b_exp2 = 10'd967; b_exp3 = 10'd868;
a_sign0 = 4'd3; a_sign1 = 4'd14; a_sign2 = 4'd12; a_sign3 = 4'd8;
b_sign0 = 4'd5; b_sign1 = 4'd7; b_sign2 = 4'd9; b_sign3 = 4'd5;
@(posedge clk_i);
a_mant0 = 8'd56; a_mant1 = 8'd118; a_mant2 = 8'd20; a_mant3 = 8'd145;
b_mant0 = 8'd180; b_mant1 = 8'd59; b_mant2 = 8'd147; b_mant3 = 8'd42;
a_exp0 = 10'd41; a_exp1 = 10'd20; a_exp2 = 10'd958; a_exp3 = 10'd229;
b_exp0 = 10'd167; b_exp1 = 10'd202; b_exp2 = 10'd95; b_exp3 = 10'd695;
a_sign0 = 4'd11; a_sign1 = 4'd9; a_sign2 = 4'd13; a_sign3 = 4'd7;
b_sign0 = 4'd4; b_sign1 = 4'd0; b_sign2 = 4'd7; b_sign3 = 4'd5;
@(posedge clk_i);
a_mant0 = 8'd97; a_mant1 = 8'd230; a_mant2 = 8'd133; a_mant3 = 8'd122;
b_mant0 = 8'd139; b_mant1 = 8'd254; b_mant2 = 8'd89; b_mant3 = 8'd87;
a_exp0 = 10'd56; a_exp1 = 10'd103; a_exp2 = 10'd618; a_exp3 = 10'd691;
b_exp0 = 10'd15; b_exp1 = 10'd856; b_exp2 = 10'd261; b_exp3 = 10'd614;
a_sign0 = 4'd4; a_sign1 = 4'd0; a_sign2 = 4'd15; a_sign3 = 4'd0;
b_sign0 = 4'd1; b_sign1 = 4'd14; b_sign2 = 4'd14; b_sign3 = 4'd11;
@(posedge clk_i);
shared_exps0 = 8'd156;
shared_exps1 = 8'd117;
a_mant0 = 8'd199; a_mant1 = 8'd107; a_mant2 = 8'd169; a_mant3 = 8'd115;
b_mant0 = 8'd170; b_mant1 = 8'd64; b_mant2 = 8'd247; b_mant3 = 8'd40;
a_exp0 = 10'd425; a_exp1 = 10'd23; a_exp2 = 10'd748; a_exp3 = 10'd646;
b_exp0 = 10'd12; b_exp1 = 10'd750; b_exp2 = 10'd784; b_exp3 = 10'd931;
a_sign0 = 4'd4; a_sign1 = 4'd12; a_sign2 = 4'd12; a_sign3 = 4'd0;
b_sign0 = 4'd14; b_sign1 = 4'd15; b_sign2 = 4'd4; b_sign3 = 4'd2;
@(posedge clk_i);
a_mant0 = 8'd214; a_mant1 = 8'd148; a_mant2 = 8'd234; a_mant3 = 8'd254;
b_mant0 = 8'd9; b_mant1 = 8'd18; b_mant2 = 8'd160; b_mant3 = 8'd159;
a_exp0 = 10'd124; a_exp1 = 10'd22; a_exp2 = 10'd474; a_exp3 = 10'd594;
b_exp0 = 10'd456; b_exp1 = 10'd776; b_exp2 = 10'd539; b_exp3 = 10'd294;
a_sign0 = 4'd5; a_sign1 = 4'd9; a_sign2 = 4'd4; a_sign3 = 4'd5;
b_sign0 = 4'd4; b_sign1 = 4'd15; b_sign2 = 4'd4; b_sign3 = 4'd8;
@(posedge clk_i);
a_mant0 = 8'd112; a_mant1 = 8'd67; a_mant2 = 8'd4; a_mant3 = 8'd241;
b_mant0 = 8'd226; b_mant1 = 8'd193; b_mant2 = 8'd7; b_mant3 = 8'd75;
a_exp0 = 10'd867; a_exp1 = 10'd457; a_exp2 = 10'd697; a_exp3 = 10'd326;
b_exp0 = 10'd172; b_exp1 = 10'd302; b_exp2 = 10'd212; b_exp3 = 10'd270;
a_sign0 = 4'd0; a_sign1 = 4'd16; a_sign2 = 4'd13; a_sign3 = 4'd4;
b_sign0 = 4'd8; b_sign1 = 4'd15; b_sign2 = 4'd3; b_sign3 = 4'd12;
@(posedge clk_i);
a_mant0 = 8'd13; a_mant1 = 8'd252; a_mant2 = 8'd2; a_mant3 = 8'd218;
b_mant0 = 8'd233; b_mant1 = 8'd158; b_mant2 = 8'd152; b_mant3 = 8'd15;
a_exp0 = 10'd185; a_exp1 = 10'd440; a_exp2 = 10'd107; a_exp3 = 10'd1015;
b_exp0 = 10'd682; b_exp1 = 10'd622; b_exp2 = 10'd183; b_exp3 = 10'd293;
a_sign0 = 4'd10; a_sign1 = 4'd4; a_sign2 = 4'd1; a_sign3 = 4'd11;
b_sign0 = 4'd6; b_sign1 = 4'd10; b_sign2 = 4'd3; b_sign3 = 4'd12;
@(posedge clk_i);
a_mant0 = 8'd243; a_mant1 = 8'd79; a_mant2 = 8'd90; a_mant3 = 8'd11;
b_mant0 = 8'd78; b_mant1 = 8'd103; b_mant2 = 8'd196; b_mant3 = 8'd225;
a_exp0 = 10'd599; a_exp1 = 10'd703; a_exp2 = 10'd479; a_exp3 = 10'd874;
b_exp0 = 10'd152; b_exp1 = 10'd701; b_exp2 = 10'd349; b_exp3 = 10'd566;
a_sign0 = 4'd5; a_sign1 = 4'd2; a_sign2 = 4'd2; a_sign3 = 4'd0;
b_sign0 = 4'd3; b_sign1 = 4'd10; b_sign2 = 4'd16; b_sign3 = 4'd6;
@(posedge clk_i);
a_mant0 = 8'd118; a_mant1 = 8'd50; a_mant2 = 8'd3; a_mant3 = 8'd16;
b_mant0 = 8'd184; b_mant1 = 8'd161; b_mant2 = 8'd194; b_mant3 = 8'd121;
a_exp0 = 10'd939; a_exp1 = 10'd811; a_exp2 = 10'd93; a_exp3 = 10'd567;
b_exp0 = 10'd913; b_exp1 = 10'd890; b_exp2 = 10'd775; b_exp3 = 10'd526;
a_sign0 = 4'd0; a_sign1 = 4'd15; a_sign2 = 4'd11; a_sign3 = 4'd5;
b_sign0 = 4'd7; b_sign1 = 4'd16; b_sign2 = 4'd5; b_sign3 = 4'd16;
@(posedge clk_i);
a_mant0 = 8'd70; a_mant1 = 8'd41; a_mant2 = 8'd74; a_mant3 = 8'd69;
b_mant0 = 8'd196; b_mant1 = 8'd176; b_mant2 = 8'd69; b_mant3 = 8'd67;
a_exp0 = 10'd871; a_exp1 = 10'd833; a_exp2 = 10'd808; a_exp3 = 10'd104;
b_exp0 = 10'd71; b_exp1 = 10'd62; b_exp2 = 10'd854; b_exp3 = 10'd279;
a_sign0 = 4'd14; a_sign1 = 4'd12; a_sign2 = 4'd16; a_sign3 = 4'd11;
b_sign0 = 4'd2; b_sign1 = 4'd6; b_sign2 = 4'd2; b_sign3 = 4'd5;
@(posedge clk_i);
a_mant0 = 8'd235; a_mant1 = 8'd60; a_mant2 = 8'd105; a_mant3 = 8'd151;
b_mant0 = 8'd182; b_mant1 = 8'd202; b_mant2 = 8'd245; b_mant3 = 8'd213;
a_exp0 = 10'd674; a_exp1 = 10'd526; a_exp2 = 10'd670; a_exp3 = 10'd184;
b_exp0 = 10'd939; b_exp1 = 10'd874; b_exp2 = 10'd87; b_exp3 = 10'd369;
a_sign0 = 4'd11; a_sign1 = 4'd6; a_sign2 = 4'd14; a_sign3 = 4'd2;
b_sign0 = 4'd1; b_sign1 = 4'd7; b_sign2 = 4'd3; b_sign3 = 4'd5;
@(posedge clk_i);
shared_exps0 = 8'd134;
shared_exps1 = 8'd109;
a_mant0 = 8'd206; a_mant1 = 8'd38; a_mant2 = 8'd110; a_mant3 = 8'd3;
b_mant0 = 8'd109; b_mant1 = 8'd112; b_mant2 = 8'd1; b_mant3 = 8'd48;
a_exp0 = 10'd243; a_exp1 = 10'd844; a_exp2 = 10'd780; a_exp3 = 10'd142;
b_exp0 = 10'd164; b_exp1 = 10'd626; b_exp2 = 10'd573; b_exp3 = 10'd694;
a_sign0 = 4'd6; a_sign1 = 4'd12; a_sign2 = 4'd16; a_sign3 = 4'd6;
b_sign0 = 4'd8; b_sign1 = 4'd12; b_sign2 = 4'd0; b_sign3 = 4'd8;
@(posedge clk_i);
a_mant0 = 8'd111; a_mant1 = 8'd44; a_mant2 = 8'd37; a_mant3 = 8'd85;
b_mant0 = 8'd25; b_mant1 = 8'd193; b_mant2 = 8'd115; b_mant3 = 8'd20;
a_exp0 = 10'd6; a_exp1 = 10'd499; a_exp2 = 10'd680; a_exp3 = 10'd322;
b_exp0 = 10'd374; b_exp1 = 10'd832; b_exp2 = 10'd267; b_exp3 = 10'd588;
a_sign0 = 4'd12; a_sign1 = 4'd9; a_sign2 = 4'd5; a_sign3 = 4'd9;
b_sign0 = 4'd9; b_sign1 = 4'd1; b_sign2 = 4'd14; b_sign3 = 4'd0;
@(posedge clk_i);
a_mant0 = 8'd13; a_mant1 = 8'd147; a_mant2 = 8'd139; a_mant3 = 8'd17;
b_mant0 = 8'd188; b_mant1 = 8'd43; b_mant2 = 8'd174; b_mant3 = 8'd46;
a_exp0 = 10'd63; a_exp1 = 10'd81; a_exp2 = 10'd679; a_exp3 = 10'd486;
b_exp0 = 10'd473; b_exp1 = 10'd161; b_exp2 = 10'd663; b_exp3 = 10'd623;
a_sign0 = 4'd16; a_sign1 = 4'd15; a_sign2 = 4'd12; a_sign3 = 4'd11;
b_sign0 = 4'd3; b_sign1 = 4'd5; b_sign2 = 4'd16; b_sign3 = 4'd8;
@(posedge clk_i);
a_mant0 = 8'd191; a_mant1 = 8'd6; a_mant2 = 8'd170; a_mant3 = 8'd91;
b_mant0 = 8'd205; b_mant1 = 8'd68; b_mant2 = 8'd178; b_mant3 = 8'd109;
a_exp0 = 10'd79; a_exp1 = 10'd119; a_exp2 = 10'd38; a_exp3 = 10'd876;
b_exp0 = 10'd1013; b_exp1 = 10'd1014; b_exp2 = 10'd955; b_exp3 = 10'd177;
a_sign0 = 4'd16; a_sign1 = 4'd11; a_sign2 = 4'd12; a_sign3 = 4'd10;
b_sign0 = 4'd8; b_sign1 = 4'd4; b_sign2 = 4'd11; b_sign3 = 4'd11;
@(posedge clk_i);
a_mant0 = 8'd60; a_mant1 = 8'd144; a_mant2 = 8'd72; a_mant3 = 8'd108;
b_mant0 = 8'd128; b_mant1 = 8'd147; b_mant2 = 8'd32; b_mant3 = 8'd238;
a_exp0 = 10'd984; a_exp1 = 10'd598; a_exp2 = 10'd460; a_exp3 = 10'd328;
b_exp0 = 10'd567; b_exp1 = 10'd991; b_exp2 = 10'd954; b_exp3 = 10'd762;
a_sign0 = 4'd13; a_sign1 = 4'd12; a_sign2 = 4'd2; a_sign3 = 4'd0;
b_sign0 = 4'd1; b_sign1 = 4'd7; b_sign2 = 4'd7; b_sign3 = 4'd5;
@(posedge clk_i);
a_mant0 = 8'd64; a_mant1 = 8'd241; a_mant2 = 8'd188; a_mant3 = 8'd167;
b_mant0 = 8'd128; b_mant1 = 8'd65; b_mant2 = 8'd205; b_mant3 = 8'd94;
a_exp0 = 10'd535; a_exp1 = 10'd521; a_exp2 = 10'd1020; a_exp3 = 10'd85;
b_exp0 = 10'd120; b_exp1 = 10'd7; b_exp2 = 10'd708; b_exp3 = 10'd872;
a_sign0 = 4'd6; a_sign1 = 4'd8; a_sign2 = 4'd0; a_sign3 = 4'd6;
b_sign0 = 4'd6; b_sign1 = 4'd0; b_sign2 = 4'd1; b_sign3 = 4'd9;
@(posedge clk_i);
a_mant0 = 8'd207; a_mant1 = 8'd236; a_mant2 = 8'd78; a_mant3 = 8'd134;
b_mant0 = 8'd107; b_mant1 = 8'd89; b_mant2 = 8'd134; b_mant3 = 8'd253;
a_exp0 = 10'd929; a_exp1 = 10'd670; a_exp2 = 10'd505; a_exp3 = 10'd543;
b_exp0 = 10'd1001; b_exp1 = 10'd774; b_exp2 = 10'd997; b_exp3 = 10'd845;
a_sign0 = 4'd3; a_sign1 = 4'd11; a_sign2 = 4'd14; a_sign3 = 4'd13;
b_sign0 = 4'd12; b_sign1 = 4'd14; b_sign2 = 4'd1; b_sign3 = 4'd16;
@(posedge clk_i);
a_mant0 = 8'd87; a_mant1 = 8'd187; a_mant2 = 8'd191; a_mant3 = 8'd162;
b_mant0 = 8'd35; b_mant1 = 8'd16; b_mant2 = 8'd236; b_mant3 = 8'd9;
a_exp0 = 10'd845; a_exp1 = 10'd815; a_exp2 = 10'd130; a_exp3 = 10'd180;
b_exp0 = 10'd182; b_exp1 = 10'd107; b_exp2 = 10'd1007; b_exp3 = 10'd657;
a_sign0 = 4'd8; a_sign1 = 4'd16; a_sign2 = 4'd3; a_sign3 = 4'd4;
b_sign0 = 4'd5; b_sign1 = 4'd8; b_sign2 = 4'd5; b_sign3 = 4'd2;
@(posedge clk_i);
shared_exps0 = 8'd135;
shared_exps1 = 8'd123;
rstn = 0;
@(posedge clk_i);
rstn = 1;
a_mant0 = 8'd144; a_mant1 = 8'd160; a_mant2 = 8'd114; a_mant3 = 8'd230;
b_mant0 = 8'd202; b_mant1 = 8'd167; b_mant2 = 8'd225; b_mant3 = 8'd64;
a_exp0 = 10'd932; a_exp1 = 10'd646; a_exp2 = 10'd294; a_exp3 = 10'd917;
b_exp0 = 10'd639; b_exp1 = 10'd884; b_exp2 = 10'd217; b_exp3 = 10'd626;
a_sign0 = 4'd8; a_sign1 = 4'd9; a_sign2 = 4'd5; a_sign3 = 4'd10;
b_sign0 = 4'd7; b_sign1 = 4'd5; b_sign2 = 4'd6; b_sign3 = 4'd13;
@(posedge clk_i);
a_mant0 = 8'd108; a_mant1 = 8'd132; a_mant2 = 8'd32; a_mant3 = 8'd180;
b_mant0 = 8'd43; b_mant1 = 8'd71; b_mant2 = 8'd178; b_mant3 = 8'd128;
a_exp0 = 10'd560; a_exp1 = 10'd496; a_exp2 = 10'd121; a_exp3 = 10'd486;
b_exp0 = 10'd952; b_exp1 = 10'd78; b_exp2 = 10'd610; b_exp3 = 10'd241;
a_sign0 = 4'd5; a_sign1 = 4'd15; a_sign2 = 4'd13; a_sign3 = 4'd3;
b_sign0 = 4'd8; b_sign1 = 4'd11; b_sign2 = 4'd12; b_sign3 = 4'd1;
@(posedge clk_i);
a_mant0 = 8'd240; a_mant1 = 8'd65; a_mant2 = 8'd239; a_mant3 = 8'd193;
b_mant0 = 8'd141; b_mant1 = 8'd243; b_mant2 = 8'd194; b_mant3 = 8'd82;
a_exp0 = 10'd699; a_exp1 = 10'd601; a_exp2 = 10'd762; a_exp3 = 10'd637;
b_exp0 = 10'd929; b_exp1 = 10'd385; b_exp2 = 10'd1011; b_exp3 = 10'd1009;
a_sign0 = 4'd3; a_sign1 = 4'd0; a_sign2 = 4'd13; a_sign3 = 4'd10;
b_sign0 = 4'd7; b_sign1 = 4'd15; b_sign2 = 4'd6; b_sign3 = 4'd2;
@(posedge clk_i);
a_mant0 = 8'd84; a_mant1 = 8'd82; a_mant2 = 8'd109; a_mant3 = 8'd81;
b_mant0 = 8'd210; b_mant1 = 8'd212; b_mant2 = 8'd213; b_mant3 = 8'd192;
a_exp0 = 10'd61; a_exp1 = 10'd757; a_exp2 = 10'd212; a_exp3 = 10'd452;
b_exp0 = 10'd817; b_exp1 = 10'd389; b_exp2 = 10'd818; b_exp3 = 10'd143;
a_sign0 = 4'd5; a_sign1 = 4'd0; a_sign2 = 4'd2; a_sign3 = 4'd7;
b_sign0 = 4'd9; b_sign1 = 4'd6; b_sign2 = 4'd7; b_sign3 = 4'd16;
@(posedge clk_i);
a_mant0 = 8'd232; a_mant1 = 8'd191; a_mant2 = 8'd162; a_mant3 = 8'd55;
b_mant0 = 8'd83; b_mant1 = 8'd156; b_mant2 = 8'd167; b_mant3 = 8'd119;
a_exp0 = 10'd649; a_exp1 = 10'd806; a_exp2 = 10'd261; a_exp3 = 10'd471;
b_exp0 = 10'd1016; b_exp1 = 10'd539; b_exp2 = 10'd821; b_exp3 = 10'd98;
a_sign0 = 4'd0; a_sign1 = 4'd4; a_sign2 = 4'd15; a_sign3 = 4'd1;
b_sign0 = 4'd4; b_sign1 = 4'd11; b_sign2 = 4'd2; b_sign3 = 4'd14;
@(posedge clk_i);
a_mant0 = 8'd123; a_mant1 = 8'd24; a_mant2 = 8'd57; a_mant3 = 8'd223;
b_mant0 = 8'd169; b_mant1 = 8'd240; b_mant2 = 8'd101; b_mant3 = 8'd166;
a_exp0 = 10'd987; a_exp1 = 10'd865; a_exp2 = 10'd94; a_exp3 = 10'd453;
b_exp0 = 10'd634; b_exp1 = 10'd683; b_exp2 = 10'd405; b_exp3 = 10'd684;
a_sign0 = 4'd1; a_sign1 = 4'd16; a_sign2 = 4'd6; a_sign3 = 4'd2;
b_sign0 = 4'd0; b_sign1 = 4'd10; b_sign2 = 4'd15; b_sign3 = 4'd5;
@(posedge clk_i);
a_mant0 = 8'd25; a_mant1 = 8'd97; a_mant2 = 8'd98; a_mant3 = 8'd63;
b_mant0 = 8'd241; b_mant1 = 8'd176; b_mant2 = 8'd37; b_mant3 = 8'd150;
a_exp0 = 10'd444; a_exp1 = 10'd221; a_exp2 = 10'd795; a_exp3 = 10'd18;
b_exp0 = 10'd743; b_exp1 = 10'd911; b_exp2 = 10'd383; b_exp3 = 10'd477;
a_sign0 = 4'd2; a_sign1 = 4'd2; a_sign2 = 4'd13; a_sign3 = 4'd3;
b_sign0 = 4'd6; b_sign1 = 4'd6; b_sign2 = 4'd15; b_sign3 = 4'd15;
@(posedge clk_i);
shared_exps0 = 8'd118;
shared_exps1 = 8'd128;
a_mant0 = 8'd122; a_mant1 = 8'd109; a_mant2 = 8'd198; a_mant3 = 8'd124;
b_mant0 = 8'd206; b_mant1 = 8'd79; b_mant2 = 8'd254; b_mant3 = 8'd203;
a_exp0 = 10'd683; a_exp1 = 10'd686; a_exp2 = 10'd510; a_exp3 = 10'd988;
b_exp0 = 10'd123; b_exp1 = 10'd434; b_exp2 = 10'd269; b_exp3 = 10'd1015;
a_sign0 = 4'd7; a_sign1 = 4'd5; a_sign2 = 4'd13; a_sign3 = 4'd8;
b_sign0 = 4'd13; b_sign1 = 4'd5; b_sign2 = 4'd1; b_sign3 = 4'd2;
@(posedge clk_i);
a_mant0 = 8'd95; a_mant1 = 8'd81; a_mant2 = 8'd122; a_mant3 = 8'd165;
b_mant0 = 8'd5; b_mant1 = 8'd33; b_mant2 = 8'd118; b_mant3 = 8'd142;
a_exp0 = 10'd102; a_exp1 = 10'd603; a_exp2 = 10'd387; a_exp3 = 10'd975;
b_exp0 = 10'd551; b_exp1 = 10'd99; b_exp2 = 10'd780; b_exp3 = 10'd911;
a_sign0 = 4'd10; a_sign1 = 4'd12; a_sign2 = 4'd9; a_sign3 = 4'd14;
b_sign0 = 4'd2; b_sign1 = 4'd3; b_sign2 = 4'd6; b_sign3 = 4'd13;
@(posedge clk_i);
a_mant0 = 8'd206; a_mant1 = 8'd19; a_mant2 = 8'd254; a_mant3 = 8'd235;
b_mant0 = 8'd133; b_mant1 = 8'd112; b_mant2 = 8'd164; b_mant3 = 8'd149;
a_exp0 = 10'd145; a_exp1 = 10'd587; a_exp2 = 10'd599; a_exp3 = 10'd701;
b_exp0 = 10'd648; b_exp1 = 10'd867; b_exp2 = 10'd808; b_exp3 = 10'd655;
a_sign0 = 4'd8; a_sign1 = 4'd4; a_sign2 = 4'd6; a_sign3 = 4'd0;
b_sign0 = 4'd11; b_sign1 = 4'd12; b_sign2 = 4'd6; b_sign3 = 4'd12;
@(posedge clk_i);
a_mant0 = 8'd22; a_mant1 = 8'd28; a_mant2 = 8'd2; a_mant3 = 8'd115;
b_mant0 = 8'd166; b_mant1 = 8'd61; b_mant2 = 8'd89; b_mant3 = 8'd19;
a_exp0 = 10'd363; a_exp1 = 10'd634; a_exp2 = 10'd532; a_exp3 = 10'd577;
b_exp0 = 10'd73; b_exp1 = 10'd748; b_exp2 = 10'd547; b_exp3 = 10'd413;
a_sign0 = 4'd6; a_sign1 = 4'd7; a_sign2 = 4'd0; a_sign3 = 4'd5;
b_sign0 = 4'd10; b_sign1 = 4'd2; b_sign2 = 4'd12; b_sign3 = 4'd1;
@(posedge clk_i);
a_mant0 = 8'd191; a_mant1 = 8'd129; a_mant2 = 8'd205; a_mant3 = 8'd111;
b_mant0 = 8'd144; b_mant1 = 8'd192; b_mant2 = 8'd184; b_mant3 = 8'd54;
a_exp0 = 10'd614; a_exp1 = 10'd682; a_exp2 = 10'd945; a_exp3 = 10'd66;
b_exp0 = 10'd718; b_exp1 = 10'd745; b_exp2 = 10'd388; b_exp3 = 10'd152;
a_sign0 = 4'd13; a_sign1 = 4'd3; a_sign2 = 4'd15; a_sign3 = 4'd9;
b_sign0 = 4'd15; b_sign1 = 4'd6; b_sign2 = 4'd7; b_sign3 = 4'd1;
@(posedge clk_i);
a_mant0 = 8'd159; a_mant1 = 8'd125; a_mant2 = 8'd61; a_mant3 = 8'd209;
b_mant0 = 8'd242; b_mant1 = 8'd107; b_mant2 = 8'd155; b_mant3 = 8'd162;
a_exp0 = 10'd676; a_exp1 = 10'd555; a_exp2 = 10'd864; a_exp3 = 10'd725;
b_exp0 = 10'd227; b_exp1 = 10'd637; b_exp2 = 10'd70; b_exp3 = 10'd977;
a_sign0 = 4'd14; a_sign1 = 4'd11; a_sign2 = 4'd5; a_sign3 = 4'd7;
b_sign0 = 4'd13; b_sign1 = 4'd1; b_sign2 = 4'd0; b_sign3 = 4'd6;
@(posedge clk_i);
a_mant0 = 8'd144; a_mant1 = 8'd162; a_mant2 = 8'd44; a_mant3 = 8'd59;
b_mant0 = 8'd54; b_mant1 = 8'd226; b_mant2 = 8'd216; b_mant3 = 8'd106;
a_exp0 = 10'd406; a_exp1 = 10'd339; a_exp2 = 10'd701; a_exp3 = 10'd367;
b_exp0 = 10'd594; b_exp1 = 10'd544; b_exp2 = 10'd419; b_exp3 = 10'd300;
a_sign0 = 4'd11; a_sign1 = 4'd9; a_sign2 = 4'd15; a_sign3 = 4'd14;
b_sign0 = 4'd11; b_sign1 = 4'd3; b_sign2 = 4'd2; b_sign3 = 4'd0;
@(posedge clk_i);
a_mant0 = 8'd232; a_mant1 = 8'd115; a_mant2 = 8'd7; a_mant3 = 8'd215;
b_mant0 = 8'd191; b_mant1 = 8'd163; b_mant2 = 8'd203; b_mant3 = 8'd107;
a_exp0 = 10'd712; a_exp1 = 10'd156; a_exp2 = 10'd95; a_exp3 = 10'd883;
b_exp0 = 10'd358; b_exp1 = 10'd764; b_exp2 = 10'd237; b_exp3 = 10'd494;
a_sign0 = 4'd15; a_sign1 = 4'd2; a_sign2 = 4'd1; a_sign3 = 4'd11;
b_sign0 = 4'd7; b_sign1 = 4'd11; b_sign2 = 4'd2; b_sign3 = 4'd16;
@(posedge clk_i);
shared_exps0 = 8'd108;
shared_exps1 = 8'd117;
a_mant0 = 8'd180; a_mant1 = 8'd138; a_mant2 = 8'd18; a_mant3 = 8'd221;
b_mant0 = 8'd112; b_mant1 = 8'd221; b_mant2 = 8'd65; b_mant3 = 8'd120;
a_exp0 = 10'd620; a_exp1 = 10'd980; a_exp2 = 10'd564; a_exp3 = 10'd622;
b_exp0 = 10'd385; b_exp1 = 10'd385; b_exp2 = 10'd41; b_exp3 = 10'd813;
a_sign0 = 4'd3; a_sign1 = 4'd1; a_sign2 = 4'd10; a_sign3 = 4'd14;
b_sign0 = 4'd2; b_sign1 = 4'd0; b_sign2 = 4'd8; b_sign3 = 4'd9;
@(posedge clk_i);
a_mant0 = 8'd15; a_mant1 = 8'd236; a_mant2 = 8'd220; a_mant3 = 8'd125;
b_mant0 = 8'd93; b_mant1 = 8'd217; b_mant2 = 8'd102; b_mant3 = 8'd59;
a_exp0 = 10'd723; a_exp1 = 10'd442; a_exp2 = 10'd472; a_exp3 = 10'd883;
b_exp0 = 10'd198; b_exp1 = 10'd62; b_exp2 = 10'd620; b_exp3 = 10'd557;
a_sign0 = 4'd13; a_sign1 = 4'd1; a_sign2 = 4'd15; a_sign3 = 4'd13;
b_sign0 = 4'd9; b_sign1 = 4'd0; b_sign2 = 4'd13; b_sign3 = 4'd13;
@(posedge clk_i);
a_mant0 = 8'd169; a_mant1 = 8'd82; a_mant2 = 8'd238; a_mant3 = 8'd58;
b_mant0 = 8'd158; b_mant1 = 8'd25; b_mant2 = 8'd248; b_mant3 = 8'd100;
a_exp0 = 10'd20; a_exp1 = 10'd76; a_exp2 = 10'd557; a_exp3 = 10'd303;
b_exp0 = 10'd66; b_exp1 = 10'd386; b_exp2 = 10'd540; b_exp3 = 10'd800;
a_sign0 = 4'd6; a_sign1 = 4'd3; a_sign2 = 4'd7; a_sign3 = 4'd0;
b_sign0 = 4'd13; b_sign1 = 4'd9; b_sign2 = 4'd0; b_sign3 = 4'd16;
@(posedge clk_i);
a_mant0 = 8'd231; a_mant1 = 8'd33; a_mant2 = 8'd228; a_mant3 = 8'd93;
b_mant0 = 8'd18; b_mant1 = 8'd97; b_mant2 = 8'd29; b_mant3 = 8'd118;
a_exp0 = 10'd471; a_exp1 = 10'd618; a_exp2 = 10'd183; a_exp3 = 10'd648;
b_exp0 = 10'd95; b_exp1 = 10'd443; b_exp2 = 10'd294; b_exp3 = 10'd817;
a_sign0 = 4'd1; a_sign1 = 4'd1; a_sign2 = 4'd3; a_sign3 = 4'd16;
b_sign0 = 4'd10; b_sign1 = 4'd13; b_sign2 = 4'd15; b_sign3 = 4'd10;
@(posedge clk_i);
a_mant0 = 8'd62; a_mant1 = 8'd156; a_mant2 = 8'd123; a_mant3 = 8'd177;
b_mant0 = 8'd187; b_mant1 = 8'd133; b_mant2 = 8'd254; b_mant3 = 8'd33;
a_exp0 = 10'd393; a_exp1 = 10'd151; a_exp2 = 10'd885; a_exp3 = 10'd640;
b_exp0 = 10'd815; b_exp1 = 10'd695; b_exp2 = 10'd226; b_exp3 = 10'd59;
a_sign0 = 4'd2; a_sign1 = 4'd12; a_sign2 = 4'd15; a_sign3 = 4'd11;
b_sign0 = 4'd7; b_sign1 = 4'd16; b_sign2 = 4'd8; b_sign3 = 4'd14;
@(posedge clk_i);
a_mant0 = 8'd239; a_mant1 = 8'd118; a_mant2 = 8'd12; a_mant3 = 8'd237;
b_mant0 = 8'd33; b_mant1 = 8'd9; b_mant2 = 8'd126; b_mant3 = 8'd253;
a_exp0 = 10'd447; a_exp1 = 10'd862; a_exp2 = 10'd962; a_exp3 = 10'd580;
b_exp0 = 10'd376; b_exp1 = 10'd910; b_exp2 = 10'd76; b_exp3 = 10'd1007;
a_sign0 = 4'd13; a_sign1 = 4'd5; a_sign2 = 4'd12; a_sign3 = 4'd1;
b_sign0 = 4'd9; b_sign1 = 4'd9; b_sign2 = 4'd6; b_sign3 = 4'd11;
@(posedge clk_i);
a_mant0 = 8'd7; a_mant1 = 8'd215; a_mant2 = 8'd198; a_mant3 = 8'd32;
b_mant0 = 8'd121; b_mant1 = 8'd225; b_mant2 = 8'd77; b_mant3 = 8'd120;
a_exp0 = 10'd198; a_exp1 = 10'd806; a_exp2 = 10'd836; a_exp3 = 10'd902;
b_exp0 = 10'd100; b_exp1 = 10'd468; b_exp2 = 10'd306; b_exp3 = 10'd792;
a_sign0 = 4'd8; a_sign1 = 4'd0; a_sign2 = 4'd5; a_sign3 = 4'd7;
b_sign0 = 4'd14; b_sign1 = 4'd4; b_sign2 = 4'd10; b_sign3 = 4'd4;
@(posedge clk_i);
a_mant0 = 8'd139; a_mant1 = 8'd189; a_mant2 = 8'd218; a_mant3 = 8'd235;
b_mant0 = 8'd188; b_mant1 = 8'd67; b_mant2 = 8'd9; b_mant3 = 8'd8;
a_exp0 = 10'd160; a_exp1 = 10'd283; a_exp2 = 10'd745; a_exp3 = 10'd805;
b_exp0 = 10'd900; b_exp1 = 10'd375; b_exp2 = 10'd317; b_exp3 = 10'd14;
a_sign0 = 4'd13; a_sign1 = 4'd6; a_sign2 = 4'd8; a_sign3 = 4'd5;
b_sign0 = 4'd15; b_sign1 = 4'd8; b_sign2 = 4'd16; b_sign3 = 4'd1;
@(posedge clk_i);
shared_exps0 = 8'd108;
shared_exps1 = 8'd144;
a_mant0 = 8'd245; a_mant1 = 8'd253; a_mant2 = 8'd186; a_mant3 = 8'd238;
b_mant0 = 8'd184; b_mant1 = 8'd35; b_mant2 = 8'd108; b_mant3 = 8'd117;
a_exp0 = 10'd486; a_exp1 = 10'd972; a_exp2 = 10'd64; a_exp3 = 10'd1017;
b_exp0 = 10'd70; b_exp1 = 10'd615; b_exp2 = 10'd225; b_exp3 = 10'd609;
a_sign0 = 4'd0; a_sign1 = 4'd4; a_sign2 = 4'd11; a_sign3 = 4'd7;
b_sign0 = 4'd0; b_sign1 = 4'd13; b_sign2 = 4'd12; b_sign3 = 4'd14;
@(posedge clk_i);
a_mant0 = 8'd245; a_mant1 = 8'd29; a_mant2 = 8'd191; a_mant3 = 8'd52;
b_mant0 = 8'd70; b_mant1 = 8'd83; b_mant2 = 8'd0; b_mant3 = 8'd55;
a_exp0 = 10'd740; a_exp1 = 10'd990; a_exp2 = 10'd890; a_exp3 = 10'd253;
b_exp0 = 10'd768; b_exp1 = 10'd987; b_exp2 = 10'd797; b_exp3 = 10'd369;
a_sign0 = 4'd8; a_sign1 = 4'd4; a_sign2 = 4'd10; a_sign3 = 4'd12;
b_sign0 = 4'd4; b_sign1 = 4'd11; b_sign2 = 4'd0; b_sign3 = 4'd5;
@(posedge clk_i);
a_mant0 = 8'd214; a_mant1 = 8'd54; a_mant2 = 8'd85; a_mant3 = 8'd159;
b_mant0 = 8'd19; b_mant1 = 8'd227; b_mant2 = 8'd50; b_mant3 = 8'd196;
a_exp0 = 10'd545; a_exp1 = 10'd253; a_exp2 = 10'd328; a_exp3 = 10'd422;
b_exp0 = 10'd872; b_exp1 = 10'd872; b_exp2 = 10'd740; b_exp3 = 10'd112;
a_sign0 = 4'd1; a_sign1 = 4'd9; a_sign2 = 4'd12; a_sign3 = 4'd10;
b_sign0 = 4'd16; b_sign1 = 4'd15; b_sign2 = 4'd5; b_sign3 = 4'd1;
@(posedge clk_i);
a_mant0 = 8'd185; a_mant1 = 8'd28; a_mant2 = 8'd185; a_mant3 = 8'd46;
b_mant0 = 8'd158; b_mant1 = 8'd0; b_mant2 = 8'd142; b_mant3 = 8'd180;
a_exp0 = 10'd370; a_exp1 = 10'd330; a_exp2 = 10'd380; a_exp3 = 10'd967;
b_exp0 = 10'd995; b_exp1 = 10'd19; b_exp2 = 10'd506; b_exp3 = 10'd14;
a_sign0 = 4'd10; a_sign1 = 4'd6; a_sign2 = 4'd13; a_sign3 = 4'd4;
b_sign0 = 4'd9; b_sign1 = 4'd3; b_sign2 = 4'd7; b_sign3 = 4'd11;
@(posedge clk_i);
a_mant0 = 8'd182; a_mant1 = 8'd86; a_mant2 = 8'd191; a_mant3 = 8'd195;
b_mant0 = 8'd192; b_mant1 = 8'd204; b_mant2 = 8'd110; b_mant3 = 8'd249;
a_exp0 = 10'd372; a_exp1 = 10'd225; a_exp2 = 10'd145; a_exp3 = 10'd1004;
b_exp0 = 10'd765; b_exp1 = 10'd360; b_exp2 = 10'd383; b_exp3 = 10'd201;
a_sign0 = 4'd11; a_sign1 = 4'd12; a_sign2 = 4'd10; a_sign3 = 4'd4;
b_sign0 = 4'd5; b_sign1 = 4'd3; b_sign2 = 4'd5; b_sign3 = 4'd15;
@(posedge clk_i);
a_mant0 = 8'd101; a_mant1 = 8'd67; a_mant2 = 8'd126; a_mant3 = 8'd117;
b_mant0 = 8'd238; b_mant1 = 8'd109; b_mant2 = 8'd31; b_mant3 = 8'd204;
a_exp0 = 10'd188; a_exp1 = 10'd415; a_exp2 = 10'd959; a_exp3 = 10'd529;
b_exp0 = 10'd106; b_exp1 = 10'd38; b_exp2 = 10'd697; b_exp3 = 10'd1000;
a_sign0 = 4'd3; a_sign1 = 4'd16; a_sign2 = 4'd5; a_sign3 = 4'd8;
b_sign0 = 4'd4; b_sign1 = 4'd7; b_sign2 = 4'd8; b_sign3 = 4'd13;
@(posedge clk_i);
a_mant0 = 8'd43; a_mant1 = 8'd61; a_mant2 = 8'd221; a_mant3 = 8'd71;
b_mant0 = 8'd232; b_mant1 = 8'd143; b_mant2 = 8'd75; b_mant3 = 8'd70;
a_exp0 = 10'd174; a_exp1 = 10'd442; a_exp2 = 10'd385; a_exp3 = 10'd69;
b_exp0 = 10'd521; b_exp1 = 10'd166; b_exp2 = 10'd314; b_exp3 = 10'd231;
a_sign0 = 4'd10; a_sign1 = 4'd8; a_sign2 = 4'd9; a_sign3 = 4'd4;
b_sign0 = 4'd2; b_sign1 = 4'd14; b_sign2 = 4'd0; b_sign3 = 4'd6;
@(posedge clk_i);
a_mant0 = 8'd42; a_mant1 = 8'd221; a_mant2 = 8'd49; a_mant3 = 8'd197;
b_mant0 = 8'd218; b_mant1 = 8'd255; b_mant2 = 8'd27; b_mant3 = 8'd61;
a_exp0 = 10'd113; a_exp1 = 10'd657; a_exp2 = 10'd512; a_exp3 = 10'd873;
b_exp0 = 10'd48; b_exp1 = 10'd652; b_exp2 = 10'd116; b_exp3 = 10'd509;
a_sign0 = 4'd14; a_sign1 = 4'd4; a_sign2 = 4'd8; a_sign3 = 4'd10;
b_sign0 = 4'd9; b_sign1 = 4'd9; b_sign2 = 4'd10; b_sign3 = 4'd1;
@(posedge clk_i);
shared_exps0 = 8'd147;
shared_exps1 = 8'd114;
rstn = 0;
@(posedge clk_i);
rstn = 1;
a_mant0 = 8'd108; a_mant1 = 8'd220; a_mant2 = 8'd150; a_mant3 = 8'd107;
b_mant0 = 8'd119; b_mant1 = 8'd94; b_mant2 = 8'd227; b_mant3 = 8'd253;
a_exp0 = 10'd54; a_exp1 = 10'd976; a_exp2 = 10'd543; a_exp3 = 10'd432;
b_exp0 = 10'd165; b_exp1 = 10'd1003; b_exp2 = 10'd720; b_exp3 = 10'd284;
a_sign0 = 4'd0; a_sign1 = 4'd14; a_sign2 = 4'd8; a_sign3 = 4'd7;
b_sign0 = 4'd1; b_sign1 = 4'd16; b_sign2 = 4'd7; b_sign3 = 4'd7;
@(posedge clk_i);
a_mant0 = 8'd18; a_mant1 = 8'd239; a_mant2 = 8'd122; a_mant3 = 8'd248;
b_mant0 = 8'd25; b_mant1 = 8'd75; b_mant2 = 8'd190; b_mant3 = 8'd238;
a_exp0 = 10'd423; a_exp1 = 10'd681; a_exp2 = 10'd325; a_exp3 = 10'd868;
b_exp0 = 10'd201; b_exp1 = 10'd546; b_exp2 = 10'd210; b_exp3 = 10'd847;
a_sign0 = 4'd6; a_sign1 = 4'd3; a_sign2 = 4'd5; a_sign3 = 4'd4;
b_sign0 = 4'd3; b_sign1 = 4'd3; b_sign2 = 4'd16; b_sign3 = 4'd8;
@(posedge clk_i);
a_mant0 = 8'd196; a_mant1 = 8'd167; a_mant2 = 8'd87; a_mant3 = 8'd98;
b_mant0 = 8'd217; b_mant1 = 8'd174; b_mant2 = 8'd208; b_mant3 = 8'd110;
a_exp0 = 10'd239; a_exp1 = 10'd544; a_exp2 = 10'd71; a_exp3 = 10'd144;
b_exp0 = 10'd317; b_exp1 = 10'd348; b_exp2 = 10'd179; b_exp3 = 10'd207;
a_sign0 = 4'd9; a_sign1 = 4'd2; a_sign2 = 4'd9; a_sign3 = 4'd13;
b_sign0 = 4'd10; b_sign1 = 4'd5; b_sign2 = 4'd8; b_sign3 = 4'd5;
@(posedge clk_i);
a_mant0 = 8'd38; a_mant1 = 8'd144; a_mant2 = 8'd126; a_mant3 = 8'd76;
b_mant0 = 8'd184; b_mant1 = 8'd254; b_mant2 = 8'd42; b_mant3 = 8'd159;
a_exp0 = 10'd739; a_exp1 = 10'd995; a_exp2 = 10'd136; a_exp3 = 10'd508;
b_exp0 = 10'd807; b_exp1 = 10'd554; b_exp2 = 10'd654; b_exp3 = 10'd90;
a_sign0 = 4'd0; a_sign1 = 4'd7; a_sign2 = 4'd8; a_sign3 = 4'd6;
b_sign0 = 4'd8; b_sign1 = 4'd5; b_sign2 = 4'd5; b_sign3 = 4'd0;
@(posedge clk_i);
a_mant0 = 8'd245; a_mant1 = 8'd167; a_mant2 = 8'd116; a_mant3 = 8'd141;
b_mant0 = 8'd237; b_mant1 = 8'd155; b_mant2 = 8'd57; b_mant3 = 8'd5;
a_exp0 = 10'd962; a_exp1 = 10'd990; a_exp2 = 10'd322; a_exp3 = 10'd489;
b_exp0 = 10'd110; b_exp1 = 10'd167; b_exp2 = 10'd348; b_exp3 = 10'd541;
a_sign0 = 4'd11; a_sign1 = 4'd0; a_sign2 = 4'd6; a_sign3 = 4'd16;
b_sign0 = 4'd16; b_sign1 = 4'd0; b_sign2 = 4'd13; b_sign3 = 4'd12;
@(posedge clk_i);
a_mant0 = 8'd43; a_mant1 = 8'd146; a_mant2 = 8'd15; a_mant3 = 8'd16;
b_mant0 = 8'd148; b_mant1 = 8'd76; b_mant2 = 8'd158; b_mant3 = 8'd129;
a_exp0 = 10'd24; a_exp1 = 10'd863; a_exp2 = 10'd796; a_exp3 = 10'd60;
b_exp0 = 10'd979; b_exp1 = 10'd180; b_exp2 = 10'd837; b_exp3 = 10'd376;
a_sign0 = 4'd16; a_sign1 = 4'd4; a_sign2 = 4'd10; a_sign3 = 4'd16;
b_sign0 = 4'd3; b_sign1 = 4'd11; b_sign2 = 4'd12; b_sign3 = 4'd1;
@(posedge clk_i);
a_mant0 = 8'd34; a_mant1 = 8'd40; a_mant2 = 8'd120; a_mant3 = 8'd62;
b_mant0 = 8'd182; b_mant1 = 8'd197; b_mant2 = 8'd189; b_mant3 = 8'd93;
a_exp0 = 10'd702; a_exp1 = 10'd34; a_exp2 = 10'd959; a_exp3 = 10'd706;
b_exp0 = 10'd439; b_exp1 = 10'd142; b_exp2 = 10'd689; b_exp3 = 10'd249;
a_sign0 = 4'd3; a_sign1 = 4'd11; a_sign2 = 4'd3; a_sign3 = 4'd0;
b_sign0 = 4'd7; b_sign1 = 4'd5; b_sign2 = 4'd12; b_sign3 = 4'd16;
@(posedge clk_i);
shared_exps0 = 8'd113;
shared_exps1 = 8'd150;
a_mant0 = 8'd209; a_mant1 = 8'd3; a_mant2 = 8'd106; a_mant3 = 8'd47;
b_mant0 = 8'd64; b_mant1 = 8'd162; b_mant2 = 8'd65; b_mant3 = 8'd35;
a_exp0 = 10'd672; a_exp1 = 10'd881; a_exp2 = 10'd617; a_exp3 = 10'd775;
b_exp0 = 10'd420; b_exp1 = 10'd761; b_exp2 = 10'd282; b_exp3 = 10'd938;
a_sign0 = 4'd8; a_sign1 = 4'd3; a_sign2 = 4'd0; a_sign3 = 4'd3;
b_sign0 = 4'd2; b_sign1 = 4'd0; b_sign2 = 4'd8; b_sign3 = 4'd9;
@(posedge clk_i);
a_mant0 = 8'd192; a_mant1 = 8'd128; a_mant2 = 8'd107; a_mant3 = 8'd56;
b_mant0 = 8'd34; b_mant1 = 8'd83; b_mant2 = 8'd39; b_mant3 = 8'd255;
a_exp0 = 10'd152; a_exp1 = 10'd14; a_exp2 = 10'd931; a_exp3 = 10'd586;
b_exp0 = 10'd826; b_exp1 = 10'd926; b_exp2 = 10'd10; b_exp3 = 10'd262;
a_sign0 = 4'd2; a_sign1 = 4'd16; a_sign2 = 4'd1; a_sign3 = 4'd9;
b_sign0 = 4'd8; b_sign1 = 4'd9; b_sign2 = 4'd4; b_sign3 = 4'd12;
@(posedge clk_i);
a_mant0 = 8'd8; a_mant1 = 8'd198; a_mant2 = 8'd189; a_mant3 = 8'd99;
b_mant0 = 8'd104; b_mant1 = 8'd255; b_mant2 = 8'd30; b_mant3 = 8'd13;
a_exp0 = 10'd62; a_exp1 = 10'd794; a_exp2 = 10'd700; a_exp3 = 10'd649;
b_exp0 = 10'd293; b_exp1 = 10'd122; b_exp2 = 10'd237; b_exp3 = 10'd270;
a_sign0 = 4'd16; a_sign1 = 4'd16; a_sign2 = 4'd10; a_sign3 = 4'd3;
b_sign0 = 4'd11; b_sign1 = 4'd7; b_sign2 = 4'd13; b_sign3 = 4'd2;
@(posedge clk_i);
a_mant0 = 8'd57; a_mant1 = 8'd238; a_mant2 = 8'd128; a_mant3 = 8'd143;
b_mant0 = 8'd233; b_mant1 = 8'd247; b_mant2 = 8'd252; b_mant3 = 8'd222;
a_exp0 = 10'd751; a_exp1 = 10'd975; a_exp2 = 10'd769; a_exp3 = 10'd241;
b_exp0 = 10'd170; b_exp1 = 10'd538; b_exp2 = 10'd276; b_exp3 = 10'd437;
a_sign0 = 4'd0; a_sign1 = 4'd6; a_sign2 = 4'd15; a_sign3 = 4'd7;
b_sign0 = 4'd10; b_sign1 = 4'd16; b_sign2 = 4'd1; b_sign3 = 4'd1;
@(posedge clk_i);
a_mant0 = 8'd96; a_mant1 = 8'd110; a_mant2 = 8'd47; a_mant3 = 8'd252;
b_mant0 = 8'd156; b_mant1 = 8'd0; b_mant2 = 8'd200; b_mant3 = 8'd198;
a_exp0 = 10'd685; a_exp1 = 10'd818; a_exp2 = 10'd342; a_exp3 = 10'd681;
b_exp0 = 10'd631; b_exp1 = 10'd662; b_exp2 = 10'd48; b_exp3 = 10'd616;
a_sign0 = 4'd6; a_sign1 = 4'd5; a_sign2 = 4'd2; a_sign3 = 4'd1;
b_sign0 = 4'd9; b_sign1 = 4'd10; b_sign2 = 4'd1; b_sign3 = 4'd14;
@(posedge clk_i);
a_mant0 = 8'd140; a_mant1 = 8'd225; a_mant2 = 8'd50; a_mant3 = 8'd122;
b_mant0 = 8'd148; b_mant1 = 8'd130; b_mant2 = 8'd14; b_mant3 = 8'd232;
a_exp0 = 10'd520; a_exp1 = 10'd392; a_exp2 = 10'd192; a_exp3 = 10'd639;
b_exp0 = 10'd848; b_exp1 = 10'd264; b_exp2 = 10'd247; b_exp3 = 10'd945;
a_sign0 = 4'd2; a_sign1 = 4'd15; a_sign2 = 4'd5; a_sign3 = 4'd15;
b_sign0 = 4'd5; b_sign1 = 4'd5; b_sign2 = 4'd3; b_sign3 = 4'd3;
@(posedge clk_i);
a_mant0 = 8'd25; a_mant1 = 8'd175; a_mant2 = 8'd170; a_mant3 = 8'd91;
b_mant0 = 8'd88; b_mant1 = 8'd147; b_mant2 = 8'd28; b_mant3 = 8'd242;
a_exp0 = 10'd311; a_exp1 = 10'd400; a_exp2 = 10'd324; a_exp3 = 10'd407;
b_exp0 = 10'd480; b_exp1 = 10'd926; b_exp2 = 10'd606; b_exp3 = 10'd781;
a_sign0 = 4'd1; a_sign1 = 4'd11; a_sign2 = 4'd8; a_sign3 = 4'd11;
b_sign0 = 4'd15; b_sign1 = 4'd9; b_sign2 = 4'd14; b_sign3 = 4'd15;
@(posedge clk_i);
a_mant0 = 8'd70; a_mant1 = 8'd86; a_mant2 = 8'd166; a_mant3 = 8'd145;
b_mant0 = 8'd167; b_mant1 = 8'd223; b_mant2 = 8'd254; b_mant3 = 8'd107;
a_exp0 = 10'd665; a_exp1 = 10'd448; a_exp2 = 10'd207; a_exp3 = 10'd755;
b_exp0 = 10'd421; b_exp1 = 10'd156; b_exp2 = 10'd151; b_exp3 = 10'd301;
a_sign0 = 4'd10; a_sign1 = 4'd0; a_sign2 = 4'd1; a_sign3 = 4'd6;
b_sign0 = 4'd14; b_sign1 = 4'd3; b_sign2 = 4'd0; b_sign3 = 4'd12;
@(posedge clk_i);
shared_exps0 = 8'd139;
shared_exps1 = 8'd147;
a_mant0 = 8'd99; a_mant1 = 8'd204; a_mant2 = 8'd225; a_mant3 = 8'd50;
b_mant0 = 8'd179; b_mant1 = 8'd56; b_mant2 = 8'd146; b_mant3 = 8'd10;
a_exp0 = 10'd800; a_exp1 = 10'd295; a_exp2 = 10'd21; a_exp3 = 10'd781;
b_exp0 = 10'd634; b_exp1 = 10'd682; b_exp2 = 10'd548; b_exp3 = 10'd169;
a_sign0 = 4'd8; a_sign1 = 4'd12; a_sign2 = 4'd1; a_sign3 = 4'd4;
b_sign0 = 4'd14; b_sign1 = 4'd10; b_sign2 = 4'd9; b_sign3 = 4'd11;
@(posedge clk_i);
a_mant0 = 8'd53; a_mant1 = 8'd214; a_mant2 = 8'd108; a_mant3 = 8'd105;
b_mant0 = 8'd161; b_mant1 = 8'd110; b_mant2 = 8'd6; b_mant3 = 8'd187;
a_exp0 = 10'd30; a_exp1 = 10'd574; a_exp2 = 10'd932; a_exp3 = 10'd232;
b_exp0 = 10'd655; b_exp1 = 10'd375; b_exp2 = 10'd627; b_exp3 = 10'd640;
a_sign0 = 4'd15; a_sign1 = 4'd4; a_sign2 = 4'd13; a_sign3 = 4'd5;
b_sign0 = 4'd13; b_sign1 = 4'd6; b_sign2 = 4'd14; b_sign3 = 4'd16;
@(posedge clk_i);
a_mant0 = 8'd126; a_mant1 = 8'd82; a_mant2 = 8'd53; a_mant3 = 8'd31;
b_mant0 = 8'd254; b_mant1 = 8'd207; b_mant2 = 8'd132; b_mant3 = 8'd210;
a_exp0 = 10'd971; a_exp1 = 10'd724; a_exp2 = 10'd225; a_exp3 = 10'd629;
b_exp0 = 10'd543; b_exp1 = 10'd724; b_exp2 = 10'd285; b_exp3 = 10'd851;
a_sign0 = 4'd2; a_sign1 = 4'd13; a_sign2 = 4'd14; a_sign3 = 4'd6;
b_sign0 = 4'd14; b_sign1 = 4'd11; b_sign2 = 4'd0; b_sign3 = 4'd1;
@(posedge clk_i);
a_mant0 = 8'd52; a_mant1 = 8'd118; a_mant2 = 8'd174; a_mant3 = 8'd122;
b_mant0 = 8'd253; b_mant1 = 8'd1; b_mant2 = 8'd49; b_mant3 = 8'd60;
a_exp0 = 10'd114; a_exp1 = 10'd589; a_exp2 = 10'd159; a_exp3 = 10'd919;
b_exp0 = 10'd858; b_exp1 = 10'd982; b_exp2 = 10'd661; b_exp3 = 10'd392;
a_sign0 = 4'd11; a_sign1 = 4'd1; a_sign2 = 4'd6; a_sign3 = 4'd2;
b_sign0 = 4'd10; b_sign1 = 4'd10; b_sign2 = 4'd12; b_sign3 = 4'd1;
@(posedge clk_i);
a_mant0 = 8'd239; a_mant1 = 8'd42; a_mant2 = 8'd99; a_mant3 = 8'd196;
b_mant0 = 8'd97; b_mant1 = 8'd114; b_mant2 = 8'd141; b_mant3 = 8'd208;
a_exp0 = 10'd104; a_exp1 = 10'd4; a_exp2 = 10'd158; a_exp3 = 10'd25;
b_exp0 = 10'd307; b_exp1 = 10'd346; b_exp2 = 10'd984; b_exp3 = 10'd749;
a_sign0 = 4'd16; a_sign1 = 4'd1; a_sign2 = 4'd1; a_sign3 = 4'd9;
b_sign0 = 4'd10; b_sign1 = 4'd15; b_sign2 = 4'd3; b_sign3 = 4'd15;
@(posedge clk_i);
a_mant0 = 8'd172; a_mant1 = 8'd197; a_mant2 = 8'd254; a_mant3 = 8'd214;
b_mant0 = 8'd88; b_mant1 = 8'd234; b_mant2 = 8'd220; b_mant3 = 8'd221;
a_exp0 = 10'd115; a_exp1 = 10'd331; a_exp2 = 10'd928; a_exp3 = 10'd620;
b_exp0 = 10'd841; b_exp1 = 10'd540; b_exp2 = 10'd1013; b_exp3 = 10'd690;
a_sign0 = 4'd11; a_sign1 = 4'd10; a_sign2 = 4'd11; a_sign3 = 4'd0;
b_sign0 = 4'd6; b_sign1 = 4'd14; b_sign2 = 4'd9; b_sign3 = 4'd1;
@(posedge clk_i);
a_mant0 = 8'd170; a_mant1 = 8'd94; a_mant2 = 8'd43; a_mant3 = 8'd90;
b_mant0 = 8'd63; b_mant1 = 8'd2; b_mant2 = 8'd105; b_mant3 = 8'd33;
a_exp0 = 10'd976; a_exp1 = 10'd564; a_exp2 = 10'd77; a_exp3 = 10'd880;
b_exp0 = 10'd333; b_exp1 = 10'd784; b_exp2 = 10'd774; b_exp3 = 10'd504;
a_sign0 = 4'd14; a_sign1 = 4'd6; a_sign2 = 4'd4; a_sign3 = 4'd8;
b_sign0 = 4'd2; b_sign1 = 4'd12; b_sign2 = 4'd14; b_sign3 = 4'd11;
@(posedge clk_i);
a_mant0 = 8'd27; a_mant1 = 8'd15; a_mant2 = 8'd208; a_mant3 = 8'd236;
b_mant0 = 8'd227; b_mant1 = 8'd223; b_mant2 = 8'd220; b_mant3 = 8'd173;
a_exp0 = 10'd183; a_exp1 = 10'd316; a_exp2 = 10'd657; a_exp3 = 10'd69;
b_exp0 = 10'd446; b_exp1 = 10'd881; b_exp2 = 10'd840; b_exp3 = 10'd782;
a_sign0 = 4'd6; a_sign1 = 4'd13; a_sign2 = 4'd10; a_sign3 = 4'd13;
b_sign0 = 4'd2; b_sign1 = 4'd5; b_sign2 = 4'd10; b_sign3 = 4'd14;
@(posedge clk_i);
shared_exps0 = 8'd108;
shared_exps1 = 8'd128;
a_mant0 = 8'd129; a_mant1 = 8'd43; a_mant2 = 8'd142; a_mant3 = 8'd248;
b_mant0 = 8'd157; b_mant1 = 8'd20; b_mant2 = 8'd179; b_mant3 = 8'd171;
a_exp0 = 10'd752; a_exp1 = 10'd675; a_exp2 = 10'd695; a_exp3 = 10'd716;
b_exp0 = 10'd218; b_exp1 = 10'd101; b_exp2 = 10'd75; b_exp3 = 10'd786;
a_sign0 = 4'd3; a_sign1 = 4'd15; a_sign2 = 4'd13; a_sign3 = 4'd4;
b_sign0 = 4'd14; b_sign1 = 4'd12; b_sign2 = 4'd3; b_sign3 = 4'd3;
@(posedge clk_i);
a_mant0 = 8'd34; a_mant1 = 8'd36; a_mant2 = 8'd216; a_mant3 = 8'd147;
b_mant0 = 8'd189; b_mant1 = 8'd99; b_mant2 = 8'd82; b_mant3 = 8'd241;
a_exp0 = 10'd218; a_exp1 = 10'd675; a_exp2 = 10'd228; a_exp3 = 10'd97;
b_exp0 = 10'd766; b_exp1 = 10'd898; b_exp2 = 10'd666; b_exp3 = 10'd241;
a_sign0 = 4'd7; a_sign1 = 4'd2; a_sign2 = 4'd3; a_sign3 = 4'd16;
b_sign0 = 4'd14; b_sign1 = 4'd5; b_sign2 = 4'd0; b_sign3 = 4'd9;
@(posedge clk_i);
a_mant0 = 8'd153; a_mant1 = 8'd12; a_mant2 = 8'd186; a_mant3 = 8'd150;
b_mant0 = 8'd239; b_mant1 = 8'd232; b_mant2 = 8'd53; b_mant3 = 8'd17;
a_exp0 = 10'd301; a_exp1 = 10'd703; a_exp2 = 10'd546; a_exp3 = 10'd130;
b_exp0 = 10'd249; b_exp1 = 10'd91; b_exp2 = 10'd344; b_exp3 = 10'd650;
a_sign0 = 4'd0; a_sign1 = 4'd9; a_sign2 = 4'd15; a_sign3 = 4'd4;
b_sign0 = 4'd14; b_sign1 = 4'd5; b_sign2 = 4'd15; b_sign3 = 4'd9;
@(posedge clk_i);
a_mant0 = 8'd19; a_mant1 = 8'd174; a_mant2 = 8'd35; a_mant3 = 8'd63;
b_mant0 = 8'd175; b_mant1 = 8'd73; b_mant2 = 8'd79; b_mant3 = 8'd70;
a_exp0 = 10'd853; a_exp1 = 10'd192; a_exp2 = 10'd575; a_exp3 = 10'd892;
b_exp0 = 10'd748; b_exp1 = 10'd714; b_exp2 = 10'd555; b_exp3 = 10'd607;
a_sign0 = 4'd13; a_sign1 = 4'd9; a_sign2 = 4'd7; a_sign3 = 4'd2;
b_sign0 = 4'd10; b_sign1 = 4'd10; b_sign2 = 4'd15; b_sign3 = 4'd2;
@(posedge clk_i);
a_mant0 = 8'd238; a_mant1 = 8'd74; a_mant2 = 8'd23; a_mant3 = 8'd208;
b_mant0 = 8'd255; b_mant1 = 8'd88; b_mant2 = 8'd113; b_mant3 = 8'd94;
a_exp0 = 10'd137; a_exp1 = 10'd112; a_exp2 = 10'd940; a_exp3 = 10'd191;
b_exp0 = 10'd550; b_exp1 = 10'd109; b_exp2 = 10'd473; b_exp3 = 10'd761;
a_sign0 = 4'd13; a_sign1 = 4'd12; a_sign2 = 4'd10; a_sign3 = 4'd3;
b_sign0 = 4'd3; b_sign1 = 4'd10; b_sign2 = 4'd13; b_sign3 = 4'd0;
@(posedge clk_i);
a_mant0 = 8'd92; a_mant1 = 8'd248; a_mant2 = 8'd207; a_mant3 = 8'd84;
b_mant0 = 8'd94; b_mant1 = 8'd203; b_mant2 = 8'd10; b_mant3 = 8'd129;
a_exp0 = 10'd68; a_exp1 = 10'd648; a_exp2 = 10'd941; a_exp3 = 10'd319;
b_exp0 = 10'd11; b_exp1 = 10'd529; b_exp2 = 10'd653; b_exp3 = 10'd21;
a_sign0 = 4'd0; a_sign1 = 4'd11; a_sign2 = 4'd16; a_sign3 = 4'd1;
b_sign0 = 4'd5; b_sign1 = 4'd0; b_sign2 = 4'd7; b_sign3 = 4'd12;
@(posedge clk_i);
a_mant0 = 8'd109; a_mant1 = 8'd86; a_mant2 = 8'd42; a_mant3 = 8'd94;
b_mant0 = 8'd59; b_mant1 = 8'd193; b_mant2 = 8'd14; b_mant3 = 8'd178;
a_exp0 = 10'd381; a_exp1 = 10'd516; a_exp2 = 10'd794; a_exp3 = 10'd187;
b_exp0 = 10'd858; b_exp1 = 10'd101; b_exp2 = 10'd917; b_exp3 = 10'd978;
a_sign0 = 4'd10; a_sign1 = 4'd13; a_sign2 = 4'd8; a_sign3 = 4'd14;
b_sign0 = 4'd14; b_sign1 = 4'd11; b_sign2 = 4'd15; b_sign3 = 4'd9;
@(posedge clk_i);
a_mant0 = 8'd199; a_mant1 = 8'd83; a_mant2 = 8'd83; a_mant3 = 8'd143;
b_mant0 = 8'd54; b_mant1 = 8'd203; b_mant2 = 8'd82; b_mant3 = 8'd134;
a_exp0 = 10'd965; a_exp1 = 10'd976; a_exp2 = 10'd81; a_exp3 = 10'd419;
b_exp0 = 10'd15; b_exp1 = 10'd900; b_exp2 = 10'd85; b_exp3 = 10'd242;
a_sign0 = 4'd8; a_sign1 = 4'd7; a_sign2 = 4'd11; a_sign3 = 4'd5;
b_sign0 = 4'd4; b_sign1 = 4'd2; b_sign2 = 4'd5; b_sign3 = 4'd6;
@(posedge clk_i);
shared_exps0 = 8'd127;
shared_exps1 = 8'd124;
rstn = 0;
@(posedge clk_i);
rstn = 1;
a_mant0 = 8'd136; a_mant1 = 8'd162; a_mant2 = 8'd175; a_mant3 = 8'd29;
b_mant0 = 8'd96; b_mant1 = 8'd163; b_mant2 = 8'd153; b_mant3 = 8'd236;
a_exp0 = 10'd977; a_exp1 = 10'd1005; a_exp2 = 10'd458; a_exp3 = 10'd60;
b_exp0 = 10'd877; b_exp1 = 10'd441; b_exp2 = 10'd671; b_exp3 = 10'd1016;
a_sign0 = 4'd8; a_sign1 = 4'd2; a_sign2 = 4'd10; a_sign3 = 4'd6;
b_sign0 = 4'd15; b_sign1 = 4'd11; b_sign2 = 4'd7; b_sign3 = 4'd14;
@(posedge clk_i);
a_mant0 = 8'd135; a_mant1 = 8'd154; a_mant2 = 8'd42; a_mant3 = 8'd231;
b_mant0 = 8'd194; b_mant1 = 8'd33; b_mant2 = 8'd104; b_mant3 = 8'd195;
a_exp0 = 10'd479; a_exp1 = 10'd380; a_exp2 = 10'd78; a_exp3 = 10'd271;
b_exp0 = 10'd1022; b_exp1 = 10'd819; b_exp2 = 10'd343; b_exp3 = 10'd610;
a_sign0 = 4'd2; a_sign1 = 4'd4; a_sign2 = 4'd12; a_sign3 = 4'd12;
b_sign0 = 4'd4; b_sign1 = 4'd13; b_sign2 = 4'd13; b_sign3 = 4'd15;
@(posedge clk_i);
a_mant0 = 8'd197; a_mant1 = 8'd147; a_mant2 = 8'd199; a_mant3 = 8'd154;
b_mant0 = 8'd127; b_mant1 = 8'd135; b_mant2 = 8'd151; b_mant3 = 8'd8;
a_exp0 = 10'd397; a_exp1 = 10'd1008; a_exp2 = 10'd435; a_exp3 = 10'd572;
b_exp0 = 10'd41; b_exp1 = 10'd37; b_exp2 = 10'd1009; b_exp3 = 10'd76;
a_sign0 = 4'd11; a_sign1 = 4'd10; a_sign2 = 4'd0; a_sign3 = 4'd14;
b_sign0 = 4'd16; b_sign1 = 4'd12; b_sign2 = 4'd2; b_sign3 = 4'd16;
@(posedge clk_i);
a_mant0 = 8'd199; a_mant1 = 8'd16; a_mant2 = 8'd141; a_mant3 = 8'd13;
b_mant0 = 8'd239; b_mant1 = 8'd101; b_mant2 = 8'd215; b_mant3 = 8'd165;
a_exp0 = 10'd133; a_exp1 = 10'd135; a_exp2 = 10'd945; a_exp3 = 10'd369;
b_exp0 = 10'd842; b_exp1 = 10'd963; b_exp2 = 10'd638; b_exp3 = 10'd144;
a_sign0 = 4'd9; a_sign1 = 4'd15; a_sign2 = 4'd6; a_sign3 = 4'd14;
b_sign0 = 4'd2; b_sign1 = 4'd4; b_sign2 = 4'd10; b_sign3 = 4'd0;
@(posedge clk_i);
a_mant0 = 8'd124; a_mant1 = 8'd218; a_mant2 = 8'd3; a_mant3 = 8'd167;
b_mant0 = 8'd79; b_mant1 = 8'd188; b_mant2 = 8'd185; b_mant3 = 8'd198;
a_exp0 = 10'd762; a_exp1 = 10'd759; a_exp2 = 10'd914; a_exp3 = 10'd972;
b_exp0 = 10'd564; b_exp1 = 10'd347; b_exp2 = 10'd575; b_exp3 = 10'd946;
a_sign0 = 4'd4; a_sign1 = 4'd14; a_sign2 = 4'd3; a_sign3 = 4'd8;
b_sign0 = 4'd1; b_sign1 = 4'd9; b_sign2 = 4'd1; b_sign3 = 4'd13;
@(posedge clk_i);
a_mant0 = 8'd13; a_mant1 = 8'd52; a_mant2 = 8'd71; a_mant3 = 8'd112;
b_mant0 = 8'd163; b_mant1 = 8'd93; b_mant2 = 8'd149; b_mant3 = 8'd251;
a_exp0 = 10'd284; a_exp1 = 10'd114; a_exp2 = 10'd70; a_exp3 = 10'd87;
b_exp0 = 10'd235; b_exp1 = 10'd673; b_exp2 = 10'd567; b_exp3 = 10'd168;
a_sign0 = 4'd10; a_sign1 = 4'd6; a_sign2 = 4'd3; a_sign3 = 4'd14;
b_sign0 = 4'd6; b_sign1 = 4'd10; b_sign2 = 4'd4; b_sign3 = 4'd12;
@(posedge clk_i);
a_mant0 = 8'd221; a_mant1 = 8'd205; a_mant2 = 8'd81; a_mant3 = 8'd45;
b_mant0 = 8'd25; b_mant1 = 8'd51; b_mant2 = 8'd44; b_mant3 = 8'd0;
a_exp0 = 10'd411; a_exp1 = 10'd64; a_exp2 = 10'd475; a_exp3 = 10'd959;
b_exp0 = 10'd1014; b_exp1 = 10'd479; b_exp2 = 10'd154; b_exp3 = 10'd835;
a_sign0 = 4'd12; a_sign1 = 4'd8; a_sign2 = 4'd6; a_sign3 = 4'd3;
b_sign0 = 4'd7; b_sign1 = 4'd9; b_sign2 = 4'd10; b_sign3 = 4'd10;
@(posedge clk_i);
shared_exps0 = 8'd114;
shared_exps1 = 8'd125;
a_mant0 = 8'd73; a_mant1 = 8'd198; a_mant2 = 8'd146; a_mant3 = 8'd51;
b_mant0 = 8'd23; b_mant1 = 8'd55; b_mant2 = 8'd204; b_mant3 = 8'd121;
a_exp0 = 10'd343; a_exp1 = 10'd767; a_exp2 = 10'd178; a_exp3 = 10'd534;
b_exp0 = 10'd285; b_exp1 = 10'd78; b_exp2 = 10'd73; b_exp3 = 10'd594;
a_sign0 = 4'd8; a_sign1 = 4'd1; a_sign2 = 4'd2; a_sign3 = 4'd4;
b_sign0 = 4'd7; b_sign1 = 4'd3; b_sign2 = 4'd6; b_sign3 = 4'd10;
@(posedge clk_i);
a_mant0 = 8'd36; a_mant1 = 8'd241; a_mant2 = 8'd199; a_mant3 = 8'd201;
b_mant0 = 8'd185; b_mant1 = 8'd110; b_mant2 = 8'd251; b_mant3 = 8'd125;
a_exp0 = 10'd527; a_exp1 = 10'd476; a_exp2 = 10'd8; a_exp3 = 10'd269;
b_exp0 = 10'd706; b_exp1 = 10'd632; b_exp2 = 10'd433; b_exp3 = 10'd699;
a_sign0 = 4'd1; a_sign1 = 4'd1; a_sign2 = 4'd1; a_sign3 = 4'd15;
b_sign0 = 4'd5; b_sign1 = 4'd6; b_sign2 = 4'd12; b_sign3 = 4'd6;
@(posedge clk_i);
a_mant0 = 8'd178; a_mant1 = 8'd90; a_mant2 = 8'd197; a_mant3 = 8'd17;
b_mant0 = 8'd17; b_mant1 = 8'd250; b_mant2 = 8'd148; b_mant3 = 8'd196;
a_exp0 = 10'd58; a_exp1 = 10'd690; a_exp2 = 10'd684; a_exp3 = 10'd794;
b_exp0 = 10'd303; b_exp1 = 10'd515; b_exp2 = 10'd812; b_exp3 = 10'd904;
a_sign0 = 4'd14; a_sign1 = 4'd3; a_sign2 = 4'd16; a_sign3 = 4'd8;
b_sign0 = 4'd11; b_sign1 = 4'd0; b_sign2 = 4'd2; b_sign3 = 4'd9;
@(posedge clk_i);
a_mant0 = 8'd146; a_mant1 = 8'd246; a_mant2 = 8'd118; a_mant3 = 8'd134;
b_mant0 = 8'd122; b_mant1 = 8'd240; b_mant2 = 8'd161; b_mant3 = 8'd84;
a_exp0 = 10'd223; a_exp1 = 10'd245; a_exp2 = 10'd325; a_exp3 = 10'd968;
b_exp0 = 10'd541; b_exp1 = 10'd444; b_exp2 = 10'd772; b_exp3 = 10'd764;
a_sign0 = 4'd15; a_sign1 = 4'd8; a_sign2 = 4'd8; a_sign3 = 4'd1;
b_sign0 = 4'd5; b_sign1 = 4'd4; b_sign2 = 4'd1; b_sign3 = 4'd14;
@(posedge clk_i);
a_mant0 = 8'd246; a_mant1 = 8'd224; a_mant2 = 8'd58; a_mant3 = 8'd94;
b_mant0 = 8'd211; b_mant1 = 8'd210; b_mant2 = 8'd207; b_mant3 = 8'd100;
a_exp0 = 10'd319; a_exp1 = 10'd918; a_exp2 = 10'd141; a_exp3 = 10'd550;
b_exp0 = 10'd85; b_exp1 = 10'd193; b_exp2 = 10'd729; b_exp3 = 10'd24;
a_sign0 = 4'd15; a_sign1 = 4'd9; a_sign2 = 4'd0; a_sign3 = 4'd3;
b_sign0 = 4'd8; b_sign1 = 4'd5; b_sign2 = 4'd16; b_sign3 = 4'd8;
@(posedge clk_i);
a_mant0 = 8'd196; a_mant1 = 8'd77; a_mant2 = 8'd243; a_mant3 = 8'd156;
b_mant0 = 8'd126; b_mant1 = 8'd166; b_mant2 = 8'd113; b_mant3 = 8'd59;
a_exp0 = 10'd593; a_exp1 = 10'd304; a_exp2 = 10'd259; a_exp3 = 10'd486;
b_exp0 = 10'd354; b_exp1 = 10'd21; b_exp2 = 10'd885; b_exp3 = 10'd606;
a_sign0 = 4'd0; a_sign1 = 4'd3; a_sign2 = 4'd15; a_sign3 = 4'd1;
b_sign0 = 4'd5; b_sign1 = 4'd3; b_sign2 = 4'd5; b_sign3 = 4'd5;
@(posedge clk_i);
a_mant0 = 8'd212; a_mant1 = 8'd38; a_mant2 = 8'd43; a_mant3 = 8'd154;
b_mant0 = 8'd12; b_mant1 = 8'd104; b_mant2 = 8'd95; b_mant3 = 8'd87;
a_exp0 = 10'd989; a_exp1 = 10'd507; a_exp2 = 10'd648; a_exp3 = 10'd672;
b_exp0 = 10'd965; b_exp1 = 10'd60; b_exp2 = 10'd722; b_exp3 = 10'd496;
a_sign0 = 4'd9; a_sign1 = 4'd9; a_sign2 = 4'd0; a_sign3 = 4'd3;
b_sign0 = 4'd14; b_sign1 = 4'd6; b_sign2 = 4'd1; b_sign3 = 4'd4;
@(posedge clk_i);
a_mant0 = 8'd112; a_mant1 = 8'd170; a_mant2 = 8'd217; a_mant3 = 8'd169;
b_mant0 = 8'd187; b_mant1 = 8'd30; b_mant2 = 8'd55; b_mant3 = 8'd148;
a_exp0 = 10'd792; a_exp1 = 10'd902; a_exp2 = 10'd271; a_exp3 = 10'd8;
b_exp0 = 10'd166; b_exp1 = 10'd225; b_exp2 = 10'd675; b_exp3 = 10'd1000;
a_sign0 = 4'd10; a_sign1 = 4'd10; a_sign2 = 4'd8; a_sign3 = 4'd11;
b_sign0 = 4'd2; b_sign1 = 4'd7; b_sign2 = 4'd7; b_sign3 = 4'd15;
@(posedge clk_i);
shared_exps0 = 8'd114;
shared_exps1 = 8'd131;
a_mant0 = 8'd152; a_mant1 = 8'd50; a_mant2 = 8'd98; a_mant3 = 8'd192;
b_mant0 = 8'd198; b_mant1 = 8'd167; b_mant2 = 8'd8; b_mant3 = 8'd168;
a_exp0 = 10'd157; a_exp1 = 10'd184; a_exp2 = 10'd684; a_exp3 = 10'd817;
b_exp0 = 10'd166; b_exp1 = 10'd75; b_exp2 = 10'd345; b_exp3 = 10'd692;
a_sign0 = 4'd10; a_sign1 = 4'd13; a_sign2 = 4'd10; a_sign3 = 4'd1;
b_sign0 = 4'd13; b_sign1 = 4'd10; b_sign2 = 4'd12; b_sign3 = 4'd0;
@(posedge clk_i);
a_mant0 = 8'd98; a_mant1 = 8'd150; a_mant2 = 8'd16; a_mant3 = 8'd226;
b_mant0 = 8'd254; b_mant1 = 8'd147; b_mant2 = 8'd116; b_mant3 = 8'd66;
a_exp0 = 10'd288; a_exp1 = 10'd573; a_exp2 = 10'd852; a_exp3 = 10'd372;
b_exp0 = 10'd836; b_exp1 = 10'd455; b_exp2 = 10'd1009; b_exp3 = 10'd205;
a_sign0 = 4'd13; a_sign1 = 4'd5; a_sign2 = 4'd11; a_sign3 = 4'd7;
b_sign0 = 4'd14; b_sign1 = 4'd1; b_sign2 = 4'd2; b_sign3 = 4'd10;
@(posedge clk_i);
a_mant0 = 8'd213; a_mant1 = 8'd184; a_mant2 = 8'd8; a_mant3 = 8'd121;
b_mant0 = 8'd247; b_mant1 = 8'd224; b_mant2 = 8'd207; b_mant3 = 8'd90;
a_exp0 = 10'd200; a_exp1 = 10'd159; a_exp2 = 10'd523; a_exp3 = 10'd1007;
b_exp0 = 10'd592; b_exp1 = 10'd963; b_exp2 = 10'd382; b_exp3 = 10'd351;
a_sign0 = 4'd4; a_sign1 = 4'd3; a_sign2 = 4'd7; a_sign3 = 4'd0;
b_sign0 = 4'd13; b_sign1 = 4'd11; b_sign2 = 4'd9; b_sign3 = 4'd6;
@(posedge clk_i);
a_mant0 = 8'd72; a_mant1 = 8'd138; a_mant2 = 8'd193; a_mant3 = 8'd87;
b_mant0 = 8'd133; b_mant1 = 8'd254; b_mant2 = 8'd54; b_mant3 = 8'd71;
a_exp0 = 10'd536; a_exp1 = 10'd3; a_exp2 = 10'd569; a_exp3 = 10'd514;
b_exp0 = 10'd263; b_exp1 = 10'd200; b_exp2 = 10'd214; b_exp3 = 10'd582;
a_sign0 = 4'd5; a_sign1 = 4'd12; a_sign2 = 4'd7; a_sign3 = 4'd14;
b_sign0 = 4'd3; b_sign1 = 4'd2; b_sign2 = 4'd16; b_sign3 = 4'd10;
@(posedge clk_i);
a_mant0 = 8'd7; a_mant1 = 8'd112; a_mant2 = 8'd158; a_mant3 = 8'd135;
b_mant0 = 8'd26; b_mant1 = 8'd64; b_mant2 = 8'd141; b_mant3 = 8'd110;
a_exp0 = 10'd776; a_exp1 = 10'd79; a_exp2 = 10'd148; a_exp3 = 10'd601;
b_exp0 = 10'd952; b_exp1 = 10'd381; b_exp2 = 10'd255; b_exp3 = 10'd629;
a_sign0 = 4'd5; a_sign1 = 4'd7; a_sign2 = 4'd11; a_sign3 = 4'd0;
b_sign0 = 4'd4; b_sign1 = 4'd7; b_sign2 = 4'd8; b_sign3 = 4'd4;
@(posedge clk_i);
a_mant0 = 8'd149; a_mant1 = 8'd95; a_mant2 = 8'd8; a_mant3 = 8'd244;
b_mant0 = 8'd7; b_mant1 = 8'd35; b_mant2 = 8'd40; b_mant3 = 8'd100;
a_exp0 = 10'd716; a_exp1 = 10'd728; a_exp2 = 10'd219; a_exp3 = 10'd370;
b_exp0 = 10'd634; b_exp1 = 10'd328; b_exp2 = 10'd1018; b_exp3 = 10'd956;
a_sign0 = 4'd16; a_sign1 = 4'd2; a_sign2 = 4'd5; a_sign3 = 4'd7;
b_sign0 = 4'd16; b_sign1 = 4'd1; b_sign2 = 4'd11; b_sign3 = 4'd14;
@(posedge clk_i);
a_mant0 = 8'd218; a_mant1 = 8'd25; a_mant2 = 8'd112; a_mant3 = 8'd156;
b_mant0 = 8'd203; b_mant1 = 8'd166; b_mant2 = 8'd253; b_mant3 = 8'd156;
a_exp0 = 10'd648; a_exp1 = 10'd69; a_exp2 = 10'd784; a_exp3 = 10'd847;
b_exp0 = 10'd995; b_exp1 = 10'd395; b_exp2 = 10'd508; b_exp3 = 10'd980;
a_sign0 = 4'd16; a_sign1 = 4'd2; a_sign2 = 4'd12; a_sign3 = 4'd15;
b_sign0 = 4'd1; b_sign1 = 4'd10; b_sign2 = 4'd6; b_sign3 = 4'd12;
@(posedge clk_i);
a_mant0 = 8'd239; a_mant1 = 8'd208; a_mant2 = 8'd21; a_mant3 = 8'd248;
b_mant0 = 8'd5; b_mant1 = 8'd90; b_mant2 = 8'd138; b_mant3 = 8'd172;
a_exp0 = 10'd141; a_exp1 = 10'd978; a_exp2 = 10'd115; a_exp3 = 10'd1006;
b_exp0 = 10'd657; b_exp1 = 10'd292; b_exp2 = 10'd28; b_exp3 = 10'd16;
a_sign0 = 4'd8; a_sign1 = 4'd7; a_sign2 = 4'd0; a_sign3 = 4'd8;
b_sign0 = 4'd9; b_sign1 = 4'd14; b_sign2 = 4'd7; b_sign3 = 4'd6;
@(posedge clk_i);
shared_exps0 = 8'd97;
shared_exps1 = 8'd102;
a_mant0 = 8'd166; a_mant1 = 8'd63; a_mant2 = 8'd18; a_mant3 = 8'd226;
b_mant0 = 8'd124; b_mant1 = 8'd77; b_mant2 = 8'd189; b_mant3 = 8'd82;
a_exp0 = 10'd540; a_exp1 = 10'd640; a_exp2 = 10'd302; a_exp3 = 10'd461;
b_exp0 = 10'd594; b_exp1 = 10'd882; b_exp2 = 10'd537; b_exp3 = 10'd119;
a_sign0 = 4'd5; a_sign1 = 4'd2; a_sign2 = 4'd14; a_sign3 = 4'd4;
b_sign0 = 4'd12; b_sign1 = 4'd12; b_sign2 = 4'd14; b_sign3 = 4'd11;
@(posedge clk_i);
a_mant0 = 8'd47; a_mant1 = 8'd119; a_mant2 = 8'd67; a_mant3 = 8'd50;
b_mant0 = 8'd20; b_mant1 = 8'd255; b_mant2 = 8'd34; b_mant3 = 8'd45;
a_exp0 = 10'd45; a_exp1 = 10'd749; a_exp2 = 10'd523; a_exp3 = 10'd697;
b_exp0 = 10'd1022; b_exp1 = 10'd141; b_exp2 = 10'd825; b_exp3 = 10'd809;
a_sign0 = 4'd2; a_sign1 = 4'd2; a_sign2 = 4'd2; a_sign3 = 4'd8;
b_sign0 = 4'd15; b_sign1 = 4'd3; b_sign2 = 4'd10; b_sign3 = 4'd2;
@(posedge clk_i);
a_mant0 = 8'd210; a_mant1 = 8'd135; a_mant2 = 8'd19; a_mant3 = 8'd233;
b_mant0 = 8'd4; b_mant1 = 8'd54; b_mant2 = 8'd26; b_mant3 = 8'd21;
a_exp0 = 10'd334; a_exp1 = 10'd176; a_exp2 = 10'd547; a_exp3 = 10'd87;
b_exp0 = 10'd516; b_exp1 = 10'd906; b_exp2 = 10'd546; b_exp3 = 10'd394;
a_sign0 = 4'd16; a_sign1 = 4'd15; a_sign2 = 4'd15; a_sign3 = 4'd4;
b_sign0 = 4'd1; b_sign1 = 4'd14; b_sign2 = 4'd15; b_sign3 = 4'd9;
@(posedge clk_i);
a_mant0 = 8'd63; a_mant1 = 8'd153; a_mant2 = 8'd52; a_mant3 = 8'd151;
b_mant0 = 8'd50; b_mant1 = 8'd213; b_mant2 = 8'd11; b_mant3 = 8'd30;
a_exp0 = 10'd733; a_exp1 = 10'd760; a_exp2 = 10'd919; a_exp3 = 10'd787;
b_exp0 = 10'd345; b_exp1 = 10'd765; b_exp2 = 10'd339; b_exp3 = 10'd607;
a_sign0 = 4'd1; a_sign1 = 4'd16; a_sign2 = 4'd9; a_sign3 = 4'd2;
b_sign0 = 4'd7; b_sign1 = 4'd2; b_sign2 = 4'd7; b_sign3 = 4'd0;
@(posedge clk_i);
a_mant0 = 8'd132; a_mant1 = 8'd146; a_mant2 = 8'd197; a_mant3 = 8'd230;
b_mant0 = 8'd252; b_mant1 = 8'd70; b_mant2 = 8'd214; b_mant3 = 8'd121;
a_exp0 = 10'd690; a_exp1 = 10'd881; a_exp2 = 10'd724; a_exp3 = 10'd665;
b_exp0 = 10'd945; b_exp1 = 10'd438; b_exp2 = 10'd491; b_exp3 = 10'd332;
a_sign0 = 4'd9; a_sign1 = 4'd11; a_sign2 = 4'd3; a_sign3 = 4'd0;
b_sign0 = 4'd13; b_sign1 = 4'd16; b_sign2 = 4'd1; b_sign3 = 4'd5;
@(posedge clk_i);
a_mant0 = 8'd168; a_mant1 = 8'd181; a_mant2 = 8'd231; a_mant3 = 8'd135;
b_mant0 = 8'd156; b_mant1 = 8'd74; b_mant2 = 8'd69; b_mant3 = 8'd69;
a_exp0 = 10'd513; a_exp1 = 10'd200; a_exp2 = 10'd10; a_exp3 = 10'd421;
b_exp0 = 10'd120; b_exp1 = 10'd899; b_exp2 = 10'd362; b_exp3 = 10'd330;
a_sign0 = 4'd14; a_sign1 = 4'd0; a_sign2 = 4'd16; a_sign3 = 4'd10;
b_sign0 = 4'd10; b_sign1 = 4'd6; b_sign2 = 4'd9; b_sign3 = 4'd16;
@(posedge clk_i);
a_mant0 = 8'd26; a_mant1 = 8'd178; a_mant2 = 8'd16; a_mant3 = 8'd217;
b_mant0 = 8'd154; b_mant1 = 8'd205; b_mant2 = 8'd26; b_mant3 = 8'd110;
a_exp0 = 10'd195; a_exp1 = 10'd358; a_exp2 = 10'd109; a_exp3 = 10'd339;
b_exp0 = 10'd100; b_exp1 = 10'd46; b_exp2 = 10'd821; b_exp3 = 10'd72;
a_sign0 = 4'd13; a_sign1 = 4'd11; a_sign2 = 4'd12; a_sign3 = 4'd7;
b_sign0 = 4'd9; b_sign1 = 4'd10; b_sign2 = 4'd8; b_sign3 = 4'd0;
@(posedge clk_i);
a_mant0 = 8'd94; a_mant1 = 8'd166; a_mant2 = 8'd142; a_mant3 = 8'd144;
b_mant0 = 8'd52; b_mant1 = 8'd188; b_mant2 = 8'd255; b_mant3 = 8'd173;
a_exp0 = 10'd249; a_exp1 = 10'd942; a_exp2 = 10'd736; a_exp3 = 10'd713;
b_exp0 = 10'd48; b_exp1 = 10'd150; b_exp2 = 10'd395; b_exp3 = 10'd371;
a_sign0 = 4'd2; a_sign1 = 4'd0; a_sign2 = 4'd4; a_sign3 = 4'd1;
b_sign0 = 4'd4; b_sign1 = 4'd7; b_sign2 = 4'd4; b_sign3 = 4'd8;
@(posedge clk_i);
shared_exps0 = 8'd108;
shared_exps1 = 8'd142;
rstn = 0;
@(posedge clk_i);
rstn = 1;
a_mant0 = 8'd114; a_mant1 = 8'd102; a_mant2 = 8'd249; a_mant3 = 8'd173;
b_mant0 = 8'd84; b_mant1 = 8'd21; b_mant2 = 8'd215; b_mant3 = 8'd17;
a_exp0 = 10'd195; a_exp1 = 10'd933; a_exp2 = 10'd7; a_exp3 = 10'd103;
b_exp0 = 10'd829; b_exp1 = 10'd253; b_exp2 = 10'd873; b_exp3 = 10'd25;
a_sign0 = 4'd4; a_sign1 = 4'd16; a_sign2 = 4'd16; a_sign3 = 4'd0;
b_sign0 = 4'd10; b_sign1 = 4'd7; b_sign2 = 4'd13; b_sign3 = 4'd1;
@(posedge clk_i);
a_mant0 = 8'd182; a_mant1 = 8'd133; a_mant2 = 8'd100; a_mant3 = 8'd93;
b_mant0 = 8'd36; b_mant1 = 8'd252; b_mant2 = 8'd238; b_mant3 = 8'd65;
a_exp0 = 10'd537; a_exp1 = 10'd353; a_exp2 = 10'd347; a_exp3 = 10'd502;
b_exp0 = 10'd796; b_exp1 = 10'd988; b_exp2 = 10'd649; b_exp3 = 10'd952;
a_sign0 = 4'd10; a_sign1 = 4'd5; a_sign2 = 4'd12; a_sign3 = 4'd8;
b_sign0 = 4'd4; b_sign1 = 4'd8; b_sign2 = 4'd11; b_sign3 = 4'd0;
@(posedge clk_i);
a_mant0 = 8'd19; a_mant1 = 8'd50; a_mant2 = 8'd234; a_mant3 = 8'd71;
b_mant0 = 8'd95; b_mant1 = 8'd19; b_mant2 = 8'd170; b_mant3 = 8'd128;
a_exp0 = 10'd469; a_exp1 = 10'd18; a_exp2 = 10'd231; a_exp3 = 10'd485;
b_exp0 = 10'd15; b_exp1 = 10'd934; b_exp2 = 10'd587; b_exp3 = 10'd453;
a_sign0 = 4'd2; a_sign1 = 4'd15; a_sign2 = 4'd11; a_sign3 = 4'd10;
b_sign0 = 4'd3; b_sign1 = 4'd8; b_sign2 = 4'd16; b_sign3 = 4'd11;
@(posedge clk_i);
a_mant0 = 8'd60; a_mant1 = 8'd49; a_mant2 = 8'd92; a_mant3 = 8'd61;
b_mant0 = 8'd149; b_mant1 = 8'd197; b_mant2 = 8'd162; b_mant3 = 8'd174;
a_exp0 = 10'd59; a_exp1 = 10'd50; a_exp2 = 10'd383; a_exp3 = 10'd713;
b_exp0 = 10'd459; b_exp1 = 10'd817; b_exp2 = 10'd993; b_exp3 = 10'd38;
a_sign0 = 4'd12; a_sign1 = 4'd14; a_sign2 = 4'd14; a_sign3 = 4'd14;
b_sign0 = 4'd6; b_sign1 = 4'd5; b_sign2 = 4'd15; b_sign3 = 4'd12;
@(posedge clk_i);
a_mant0 = 8'd206; a_mant1 = 8'd76; a_mant2 = 8'd43; a_mant3 = 8'd45;
b_mant0 = 8'd112; b_mant1 = 8'd141; b_mant2 = 8'd154; b_mant3 = 8'd207;
a_exp0 = 10'd893; a_exp1 = 10'd822; a_exp2 = 10'd235; a_exp3 = 10'd225;
b_exp0 = 10'd24; b_exp1 = 10'd291; b_exp2 = 10'd832; b_exp3 = 10'd932;
a_sign0 = 4'd9; a_sign1 = 4'd10; a_sign2 = 4'd9; a_sign3 = 4'd10;
b_sign0 = 4'd5; b_sign1 = 4'd11; b_sign2 = 4'd16; b_sign3 = 4'd16;
@(posedge clk_i);
a_mant0 = 8'd249; a_mant1 = 8'd117; a_mant2 = 8'd173; a_mant3 = 8'd6;
b_mant0 = 8'd143; b_mant1 = 8'd20; b_mant2 = 8'd246; b_mant3 = 8'd219;
a_exp0 = 10'd97; a_exp1 = 10'd596; a_exp2 = 10'd203; a_exp3 = 10'd146;
b_exp0 = 10'd107; b_exp1 = 10'd431; b_exp2 = 10'd625; b_exp3 = 10'd588;
a_sign0 = 4'd15; a_sign1 = 4'd10; a_sign2 = 4'd12; a_sign3 = 4'd3;
b_sign0 = 4'd7; b_sign1 = 4'd6; b_sign2 = 4'd1; b_sign3 = 4'd10;
@(posedge clk_i);
a_mant0 = 8'd142; a_mant1 = 8'd47; a_mant2 = 8'd180; a_mant3 = 8'd191;
b_mant0 = 8'd209; b_mant1 = 8'd236; b_mant2 = 8'd233; b_mant3 = 8'd138;
a_exp0 = 10'd503; a_exp1 = 10'd831; a_exp2 = 10'd1002; a_exp3 = 10'd298;
b_exp0 = 10'd455; b_exp1 = 10'd854; b_exp2 = 10'd840; b_exp3 = 10'd708;
a_sign0 = 4'd1; a_sign1 = 4'd5; a_sign2 = 4'd2; a_sign3 = 4'd5;
b_sign0 = 4'd6; b_sign1 = 4'd3; b_sign2 = 4'd2; b_sign3 = 4'd6;
@(posedge clk_i);
shared_exps0 = 8'd127;
shared_exps1 = 8'd121;
a_mant0 = 8'd62; a_mant1 = 8'd62; a_mant2 = 8'd64; a_mant3 = 8'd250;
b_mant0 = 8'd110; b_mant1 = 8'd160; b_mant2 = 8'd48; b_mant3 = 8'd128;
a_exp0 = 10'd1021; a_exp1 = 10'd117; a_exp2 = 10'd297; a_exp3 = 10'd447;
b_exp0 = 10'd420; b_exp1 = 10'd415; b_exp2 = 10'd56; b_exp3 = 10'd918;
a_sign0 = 4'd11; a_sign1 = 4'd16; a_sign2 = 4'd9; a_sign3 = 4'd8;
b_sign0 = 4'd3; b_sign1 = 4'd12; b_sign2 = 4'd8; b_sign3 = 4'd5;
@(posedge clk_i);
a_mant0 = 8'd98; a_mant1 = 8'd139; a_mant2 = 8'd140; a_mant3 = 8'd231;
b_mant0 = 8'd5; b_mant1 = 8'd131; b_mant2 = 8'd241; b_mant3 = 8'd207;
a_exp0 = 10'd141; a_exp1 = 10'd389; a_exp2 = 10'd605; a_exp3 = 10'd792;
b_exp0 = 10'd525; b_exp1 = 10'd501; b_exp2 = 10'd675; b_exp3 = 10'd238;
a_sign0 = 4'd2; a_sign1 = 4'd3; a_sign2 = 4'd11; a_sign3 = 4'd8;
b_sign0 = 4'd5; b_sign1 = 4'd13; b_sign2 = 4'd5; b_sign3 = 4'd4;
@(posedge clk_i);
a_mant0 = 8'd118; a_mant1 = 8'd10; a_mant2 = 8'd167; a_mant3 = 8'd151;
b_mant0 = 8'd162; b_mant1 = 8'd223; b_mant2 = 8'd240; b_mant3 = 8'd190;
a_exp0 = 10'd234; a_exp1 = 10'd333; a_exp2 = 10'd816; a_exp3 = 10'd380;
b_exp0 = 10'd672; b_exp1 = 10'd868; b_exp2 = 10'd302; b_exp3 = 10'd116;
a_sign0 = 4'd14; a_sign1 = 4'd1; a_sign2 = 4'd15; a_sign3 = 4'd11;
b_sign0 = 4'd5; b_sign1 = 4'd12; b_sign2 = 4'd9; b_sign3 = 4'd0;
@(posedge clk_i);
a_mant0 = 8'd252; a_mant1 = 8'd251; a_mant2 = 8'd241; a_mant3 = 8'd241;
b_mant0 = 8'd200; b_mant1 = 8'd131; b_mant2 = 8'd233; b_mant3 = 8'd210;
a_exp0 = 10'd888; a_exp1 = 10'd697; a_exp2 = 10'd999; a_exp3 = 10'd446;
b_exp0 = 10'd76; b_exp1 = 10'd1019; b_exp2 = 10'd188; b_exp3 = 10'd80;
a_sign0 = 4'd6; a_sign1 = 4'd2; a_sign2 = 4'd12; a_sign3 = 4'd2;
b_sign0 = 4'd2; b_sign1 = 4'd3; b_sign2 = 4'd13; b_sign3 = 4'd16;
@(posedge clk_i);
a_mant0 = 8'd113; a_mant1 = 8'd206; a_mant2 = 8'd136; a_mant3 = 8'd114;
b_mant0 = 8'd102; b_mant1 = 8'd20; b_mant2 = 8'd246; b_mant3 = 8'd20;
a_exp0 = 10'd949; a_exp1 = 10'd459; a_exp2 = 10'd243; a_exp3 = 10'd289;
b_exp0 = 10'd260; b_exp1 = 10'd697; b_exp2 = 10'd842; b_exp3 = 10'd750;
a_sign0 = 4'd7; a_sign1 = 4'd3; a_sign2 = 4'd13; a_sign3 = 4'd9;
b_sign0 = 4'd3; b_sign1 = 4'd15; b_sign2 = 4'd7; b_sign3 = 4'd9;
@(posedge clk_i);
a_mant0 = 8'd170; a_mant1 = 8'd111; a_mant2 = 8'd225; a_mant3 = 8'd121;
b_mant0 = 8'd204; b_mant1 = 8'd69; b_mant2 = 8'd10; b_mant3 = 8'd19;
a_exp0 = 10'd830; a_exp1 = 10'd864; a_exp2 = 10'd149; a_exp3 = 10'd564;
b_exp0 = 10'd930; b_exp1 = 10'd712; b_exp2 = 10'd457; b_exp3 = 10'd708;
a_sign0 = 4'd5; a_sign1 = 4'd1; a_sign2 = 4'd2; a_sign3 = 4'd3;
b_sign0 = 4'd0; b_sign1 = 4'd14; b_sign2 = 4'd11; b_sign3 = 4'd7;
@(posedge clk_i);
a_mant0 = 8'd4; a_mant1 = 8'd133; a_mant2 = 8'd21; a_mant3 = 8'd1;
b_mant0 = 8'd20; b_mant1 = 8'd139; b_mant2 = 8'd209; b_mant3 = 8'd119;
a_exp0 = 10'd675; a_exp1 = 10'd295; a_exp2 = 10'd558; a_exp3 = 10'd513;
b_exp0 = 10'd654; b_exp1 = 10'd32; b_exp2 = 10'd918; b_exp3 = 10'd685;
a_sign0 = 4'd12; a_sign1 = 4'd8; a_sign2 = 4'd14; a_sign3 = 4'd11;
b_sign0 = 4'd4; b_sign1 = 4'd16; b_sign2 = 4'd12; b_sign3 = 4'd9;
@(posedge clk_i);
a_mant0 = 8'd131; a_mant1 = 8'd90; a_mant2 = 8'd51; a_mant3 = 8'd147;
b_mant0 = 8'd183; b_mant1 = 8'd232; b_mant2 = 8'd122; b_mant3 = 8'd66;
a_exp0 = 10'd714; a_exp1 = 10'd994; a_exp2 = 10'd186; a_exp3 = 10'd107;
b_exp0 = 10'd886; b_exp1 = 10'd934; b_exp2 = 10'd583; b_exp3 = 10'd393;
a_sign0 = 4'd4; a_sign1 = 4'd3; a_sign2 = 4'd2; a_sign3 = 4'd1;
b_sign0 = 4'd14; b_sign1 = 4'd6; b_sign2 = 4'd5; b_sign3 = 4'd6;
@(posedge clk_i);
shared_exps0 = 8'd104;
shared_exps1 = 8'd103;
a_mant0 = 8'd230; a_mant1 = 8'd2; a_mant2 = 8'd206; a_mant3 = 8'd116;
b_mant0 = 8'd240; b_mant1 = 8'd189; b_mant2 = 8'd110; b_mant3 = 8'd172;
a_exp0 = 10'd762; a_exp1 = 10'd131; a_exp2 = 10'd990; a_exp3 = 10'd866;
b_exp0 = 10'd429; b_exp1 = 10'd439; b_exp2 = 10'd900; b_exp3 = 10'd350;
a_sign0 = 4'd3; a_sign1 = 4'd12; a_sign2 = 4'd4; a_sign3 = 4'd0;
b_sign0 = 4'd4; b_sign1 = 4'd5; b_sign2 = 4'd2; b_sign3 = 4'd8;
@(posedge clk_i);
a_mant0 = 8'd215; a_mant1 = 8'd26; a_mant2 = 8'd223; a_mant3 = 8'd249;
b_mant0 = 8'd128; b_mant1 = 8'd48; b_mant2 = 8'd113; b_mant3 = 8'd245;
a_exp0 = 10'd827; a_exp1 = 10'd967; a_exp2 = 10'd598; a_exp3 = 10'd312;
b_exp0 = 10'd865; b_exp1 = 10'd976; b_exp2 = 10'd532; b_exp3 = 10'd163;
a_sign0 = 4'd10; a_sign1 = 4'd2; a_sign2 = 4'd14; a_sign3 = 4'd14;
b_sign0 = 4'd2; b_sign1 = 4'd11; b_sign2 = 4'd16; b_sign3 = 4'd4;
@(posedge clk_i);
a_mant0 = 8'd84; a_mant1 = 8'd131; a_mant2 = 8'd12; a_mant3 = 8'd229;
b_mant0 = 8'd37; b_mant1 = 8'd64; b_mant2 = 8'd225; b_mant3 = 8'd243;
a_exp0 = 10'd788; a_exp1 = 10'd836; a_exp2 = 10'd753; a_exp3 = 10'd697;
b_exp0 = 10'd434; b_exp1 = 10'd995; b_exp2 = 10'd127; b_exp3 = 10'd928;
a_sign0 = 4'd12; a_sign1 = 4'd7; a_sign2 = 4'd5; a_sign3 = 4'd8;
b_sign0 = 4'd16; b_sign1 = 4'd12; b_sign2 = 4'd6; b_sign3 = 4'd5;
@(posedge clk_i);
a_mant0 = 8'd55; a_mant1 = 8'd41; a_mant2 = 8'd202; a_mant3 = 8'd120;
b_mant0 = 8'd243; b_mant1 = 8'd144; b_mant2 = 8'd133; b_mant3 = 8'd177;
a_exp0 = 10'd816; a_exp1 = 10'd502; a_exp2 = 10'd539; a_exp3 = 10'd552;
b_exp0 = 10'd500; b_exp1 = 10'd650; b_exp2 = 10'd176; b_exp3 = 10'd834;
a_sign0 = 4'd3; a_sign1 = 4'd13; a_sign2 = 4'd9; a_sign3 = 4'd14;
b_sign0 = 4'd1; b_sign1 = 4'd4; b_sign2 = 4'd16; b_sign3 = 4'd12;
@(posedge clk_i);
a_mant0 = 8'd185; a_mant1 = 8'd239; a_mant2 = 8'd66; a_mant3 = 8'd64;
b_mant0 = 8'd179; b_mant1 = 8'd217; b_mant2 = 8'd103; b_mant3 = 8'd134;
a_exp0 = 10'd209; a_exp1 = 10'd638; a_exp2 = 10'd696; a_exp3 = 10'd681;
b_exp0 = 10'd368; b_exp1 = 10'd263; b_exp2 = 10'd793; b_exp3 = 10'd18;
a_sign0 = 4'd9; a_sign1 = 4'd13; a_sign2 = 4'd7; a_sign3 = 4'd4;
b_sign0 = 4'd13; b_sign1 = 4'd2; b_sign2 = 4'd4; b_sign3 = 4'd0;
@(posedge clk_i);
a_mant0 = 8'd2; a_mant1 = 8'd225; a_mant2 = 8'd148; a_mant3 = 8'd48;
b_mant0 = 8'd5; b_mant1 = 8'd123; b_mant2 = 8'd140; b_mant3 = 8'd79;
a_exp0 = 10'd221; a_exp1 = 10'd878; a_exp2 = 10'd601; a_exp3 = 10'd816;
b_exp0 = 10'd577; b_exp1 = 10'd882; b_exp2 = 10'd935; b_exp3 = 10'd915;
a_sign0 = 4'd7; a_sign1 = 4'd5; a_sign2 = 4'd1; a_sign3 = 4'd14;
b_sign0 = 4'd10; b_sign1 = 4'd15; b_sign2 = 4'd10; b_sign3 = 4'd15;
@(posedge clk_i);
a_mant0 = 8'd148; a_mant1 = 8'd215; a_mant2 = 8'd221; a_mant3 = 8'd104;
b_mant0 = 8'd120; b_mant1 = 8'd117; b_mant2 = 8'd254; b_mant3 = 8'd144;
a_exp0 = 10'd750; a_exp1 = 10'd140; a_exp2 = 10'd961; a_exp3 = 10'd702;
b_exp0 = 10'd353; b_exp1 = 10'd613; b_exp2 = 10'd664; b_exp3 = 10'd679;
a_sign0 = 4'd16; a_sign1 = 4'd9; a_sign2 = 4'd12; a_sign3 = 4'd11;
b_sign0 = 4'd0; b_sign1 = 4'd1; b_sign2 = 4'd7; b_sign3 = 4'd15;
@(posedge clk_i);
a_mant0 = 8'd106; a_mant1 = 8'd136; a_mant2 = 8'd125; a_mant3 = 8'd25;
b_mant0 = 8'd69; b_mant1 = 8'd37; b_mant2 = 8'd147; b_mant3 = 8'd71;
a_exp0 = 10'd247; a_exp1 = 10'd434; a_exp2 = 10'd79; a_exp3 = 10'd789;
b_exp0 = 10'd375; b_exp1 = 10'd902; b_exp2 = 10'd44; b_exp3 = 10'd959;
a_sign0 = 4'd1; a_sign1 = 4'd5; a_sign2 = 4'd5; a_sign3 = 4'd8;
b_sign0 = 4'd11; b_sign1 = 4'd8; b_sign2 = 4'd5; b_sign3 = 4'd2;
@(posedge clk_i);
shared_exps0 = 8'd146;
shared_exps1 = 8'd138;
a_mant0 = 8'd142; a_mant1 = 8'd2; a_mant2 = 8'd70; a_mant3 = 8'd96;
b_mant0 = 8'd151; b_mant1 = 8'd83; b_mant2 = 8'd86; b_mant3 = 8'd54;
a_exp0 = 10'd371; a_exp1 = 10'd920; a_exp2 = 10'd708; a_exp3 = 10'd19;
b_exp0 = 10'd433; b_exp1 = 10'd892; b_exp2 = 10'd596; b_exp3 = 10'd549;
a_sign0 = 4'd5; a_sign1 = 4'd14; a_sign2 = 4'd0; a_sign3 = 4'd8;
b_sign0 = 4'd0; b_sign1 = 4'd15; b_sign2 = 4'd9; b_sign3 = 4'd14;
@(posedge clk_i);
a_mant0 = 8'd76; a_mant1 = 8'd73; a_mant2 = 8'd57; a_mant3 = 8'd36;
b_mant0 = 8'd29; b_mant1 = 8'd118; b_mant2 = 8'd91; b_mant3 = 8'd233;
a_exp0 = 10'd84; a_exp1 = 10'd942; a_exp2 = 10'd78; a_exp3 = 10'd364;
b_exp0 = 10'd961; b_exp1 = 10'd523; b_exp2 = 10'd958; b_exp3 = 10'd381;
a_sign0 = 4'd13; a_sign1 = 4'd13; a_sign2 = 4'd1; a_sign3 = 4'd15;
b_sign0 = 4'd11; b_sign1 = 4'd3; b_sign2 = 4'd8; b_sign3 = 4'd0;
@(posedge clk_i);
a_mant0 = 8'd203; a_mant1 = 8'd33; a_mant2 = 8'd28; a_mant3 = 8'd104;
b_mant0 = 8'd250; b_mant1 = 8'd163; b_mant2 = 8'd83; b_mant3 = 8'd194;
a_exp0 = 10'd627; a_exp1 = 10'd315; a_exp2 = 10'd698; a_exp3 = 10'd364;
b_exp0 = 10'd888; b_exp1 = 10'd1016; b_exp2 = 10'd766; b_exp3 = 10'd410;
a_sign0 = 4'd11; a_sign1 = 4'd7; a_sign2 = 4'd16; a_sign3 = 4'd9;
b_sign0 = 4'd7; b_sign1 = 4'd1; b_sign2 = 4'd10; b_sign3 = 4'd11;
@(posedge clk_i);
a_mant0 = 8'd32; a_mant1 = 8'd253; a_mant2 = 8'd2; a_mant3 = 8'd228;
b_mant0 = 8'd203; b_mant1 = 8'd70; b_mant2 = 8'd75; b_mant3 = 8'd58;
a_exp0 = 10'd586; a_exp1 = 10'd723; a_exp2 = 10'd51; a_exp3 = 10'd210;
b_exp0 = 10'd126; b_exp1 = 10'd526; b_exp2 = 10'd124; b_exp3 = 10'd147;
a_sign0 = 4'd16; a_sign1 = 4'd11; a_sign2 = 4'd10; a_sign3 = 4'd12;
b_sign0 = 4'd10; b_sign1 = 4'd13; b_sign2 = 4'd8; b_sign3 = 4'd14;
@(posedge clk_i);
a_mant0 = 8'd23; a_mant1 = 8'd30; a_mant2 = 8'd202; a_mant3 = 8'd195;
b_mant0 = 8'd111; b_mant1 = 8'd57; b_mant2 = 8'd30; b_mant3 = 8'd212;
a_exp0 = 10'd786; a_exp1 = 10'd584; a_exp2 = 10'd198; a_exp3 = 10'd574;
b_exp0 = 10'd364; b_exp1 = 10'd517; b_exp2 = 10'd957; b_exp3 = 10'd543;
a_sign0 = 4'd6; a_sign1 = 4'd3; a_sign2 = 4'd15; a_sign3 = 4'd15;
b_sign0 = 4'd9; b_sign1 = 4'd8; b_sign2 = 4'd8; b_sign3 = 4'd11;
@(posedge clk_i);
a_mant0 = 8'd219; a_mant1 = 8'd250; a_mant2 = 8'd104; a_mant3 = 8'd195;
b_mant0 = 8'd118; b_mant1 = 8'd123; b_mant2 = 8'd23; b_mant3 = 8'd95;
a_exp0 = 10'd151; a_exp1 = 10'd418; a_exp2 = 10'd476; a_exp3 = 10'd852;
b_exp0 = 10'd301; b_exp1 = 10'd717; b_exp2 = 10'd874; b_exp3 = 10'd43;
a_sign0 = 4'd13; a_sign1 = 4'd2; a_sign2 = 4'd8; a_sign3 = 4'd15;
b_sign0 = 4'd0; b_sign1 = 4'd13; b_sign2 = 4'd14; b_sign3 = 4'd16;
@(posedge clk_i);
a_mant0 = 8'd132; a_mant1 = 8'd246; a_mant2 = 8'd229; a_mant3 = 8'd195;
b_mant0 = 8'd127; b_mant1 = 8'd168; b_mant2 = 8'd210; b_mant3 = 8'd222;
a_exp0 = 10'd121; a_exp1 = 10'd84; a_exp2 = 10'd183; a_exp3 = 10'd273;
b_exp0 = 10'd311; b_exp1 = 10'd788; b_exp2 = 10'd402; b_exp3 = 10'd882;
a_sign0 = 4'd12; a_sign1 = 4'd5; a_sign2 = 4'd1; a_sign3 = 4'd9;
b_sign0 = 4'd16; b_sign1 = 4'd3; b_sign2 = 4'd1; b_sign3 = 4'd3;
@(posedge clk_i);
a_mant0 = 8'd100; a_mant1 = 8'd206; a_mant2 = 8'd141; a_mant3 = 8'd162;
b_mant0 = 8'd98; b_mant1 = 8'd138; b_mant2 = 8'd17; b_mant3 = 8'd99;
a_exp0 = 10'd597; a_exp1 = 10'd965; a_exp2 = 10'd555; a_exp3 = 10'd363;
b_exp0 = 10'd212; b_exp1 = 10'd1022; b_exp2 = 10'd342; b_exp3 = 10'd582;
a_sign0 = 4'd16; a_sign1 = 4'd10; a_sign2 = 4'd15; a_sign3 = 4'd2;
b_sign0 = 4'd4; b_sign1 = 4'd1; b_sign2 = 4'd7; b_sign3 = 4'd16;
@(posedge clk_i);
shared_exps0 = 8'd139;
shared_exps1 = 8'd139;
rstn = 0;
@(posedge clk_i);
rstn = 1;
a_mant0 = 8'd101; a_mant1 = 8'd111; a_mant2 = 8'd15; a_mant3 = 8'd122;
b_mant0 = 8'd170; b_mant1 = 8'd113; b_mant2 = 8'd110; b_mant3 = 8'd96;
a_exp0 = 10'd423; a_exp1 = 10'd426; a_exp2 = 10'd232; a_exp3 = 10'd705;
b_exp0 = 10'd480; b_exp1 = 10'd436; b_exp2 = 10'd809; b_exp3 = 10'd5;
a_sign0 = 4'd15; a_sign1 = 4'd11; a_sign2 = 4'd4; a_sign3 = 4'd15;
b_sign0 = 4'd13; b_sign1 = 4'd3; b_sign2 = 4'd9; b_sign3 = 4'd1;
@(posedge clk_i);
a_mant0 = 8'd130; a_mant1 = 8'd59; a_mant2 = 8'd35; a_mant3 = 8'd243;
b_mant0 = 8'd235; b_mant1 = 8'd92; b_mant2 = 8'd1; b_mant3 = 8'd103;
a_exp0 = 10'd238; a_exp1 = 10'd139; a_exp2 = 10'd133; a_exp3 = 10'd986;
b_exp0 = 10'd604; b_exp1 = 10'd854; b_exp2 = 10'd165; b_exp3 = 10'd278;
a_sign0 = 4'd9; a_sign1 = 4'd7; a_sign2 = 4'd4; a_sign3 = 4'd7;
b_sign0 = 4'd1; b_sign1 = 4'd16; b_sign2 = 4'd16; b_sign3 = 4'd1;
@(posedge clk_i);
a_mant0 = 8'd80; a_mant1 = 8'd193; a_mant2 = 8'd141; a_mant3 = 8'd153;
b_mant0 = 8'd205; b_mant1 = 8'd44; b_mant2 = 8'd165; b_mant3 = 8'd184;
a_exp0 = 10'd823; a_exp1 = 10'd775; a_exp2 = 10'd1001; a_exp3 = 10'd1020;
b_exp0 = 10'd195; b_exp1 = 10'd68; b_exp2 = 10'd592; b_exp3 = 10'd984;
a_sign0 = 4'd12; a_sign1 = 4'd4; a_sign2 = 4'd2; a_sign3 = 4'd16;
b_sign0 = 4'd1; b_sign1 = 4'd2; b_sign2 = 4'd14; b_sign3 = 4'd13;
@(posedge clk_i);
a_mant0 = 8'd232; a_mant1 = 8'd220; a_mant2 = 8'd211; a_mant3 = 8'd150;
b_mant0 = 8'd159; b_mant1 = 8'd182; b_mant2 = 8'd255; b_mant3 = 8'd52;
a_exp0 = 10'd976; a_exp1 = 10'd961; a_exp2 = 10'd812; a_exp3 = 10'd641;
b_exp0 = 10'd126; b_exp1 = 10'd823; b_exp2 = 10'd853; b_exp3 = 10'd870;
a_sign0 = 4'd8; a_sign1 = 4'd12; a_sign2 = 4'd12; a_sign3 = 4'd11;
b_sign0 = 4'd16; b_sign1 = 4'd0; b_sign2 = 4'd2; b_sign3 = 4'd11;
@(posedge clk_i);
a_mant0 = 8'd98; a_mant1 = 8'd152; a_mant2 = 8'd42; a_mant3 = 8'd164;
b_mant0 = 8'd243; b_mant1 = 8'd121; b_mant2 = 8'd200; b_mant3 = 8'd69;
a_exp0 = 10'd321; a_exp1 = 10'd648; a_exp2 = 10'd78; a_exp3 = 10'd728;
b_exp0 = 10'd789; b_exp1 = 10'd602; b_exp2 = 10'd517; b_exp3 = 10'd321;
a_sign0 = 4'd0; a_sign1 = 4'd9; a_sign2 = 4'd0; a_sign3 = 4'd10;
b_sign0 = 4'd2; b_sign1 = 4'd7; b_sign2 = 4'd12; b_sign3 = 4'd10;
@(posedge clk_i);
a_mant0 = 8'd14; a_mant1 = 8'd181; a_mant2 = 8'd32; a_mant3 = 8'd152;
b_mant0 = 8'd205; b_mant1 = 8'd19; b_mant2 = 8'd127; b_mant3 = 8'd23;
a_exp0 = 10'd899; a_exp1 = 10'd908; a_exp2 = 10'd365; a_exp3 = 10'd997;
b_exp0 = 10'd9; b_exp1 = 10'd614; b_exp2 = 10'd191; b_exp3 = 10'd943;
a_sign0 = 4'd3; a_sign1 = 4'd3; a_sign2 = 4'd1; a_sign3 = 4'd0;
b_sign0 = 4'd6; b_sign1 = 4'd6; b_sign2 = 4'd0; b_sign3 = 4'd0;
@(posedge clk_i);
a_mant0 = 8'd133; a_mant1 = 8'd26; a_mant2 = 8'd227; a_mant3 = 8'd203;
b_mant0 = 8'd145; b_mant1 = 8'd63; b_mant2 = 8'd56; b_mant3 = 8'd129;
a_exp0 = 10'd619; a_exp1 = 10'd903; a_exp2 = 10'd71; a_exp3 = 10'd870;
b_exp0 = 10'd909; b_exp1 = 10'd852; b_exp2 = 10'd820; b_exp3 = 10'd227;
a_sign0 = 4'd4; a_sign1 = 4'd9; a_sign2 = 4'd4; a_sign3 = 4'd11;
b_sign0 = 4'd5; b_sign1 = 4'd2; b_sign2 = 4'd2; b_sign3 = 4'd10;
@(posedge clk_i);
shared_exps0 = 8'd141;
shared_exps1 = 8'd151;
a_mant0 = 8'd92; a_mant1 = 8'd138; a_mant2 = 8'd156; a_mant3 = 8'd140;
b_mant0 = 8'd102; b_mant1 = 8'd253; b_mant2 = 8'd39; b_mant3 = 8'd119;
a_exp0 = 10'd146; a_exp1 = 10'd0; a_exp2 = 10'd747; a_exp3 = 10'd61;
b_exp0 = 10'd142; b_exp1 = 10'd154; b_exp2 = 10'd272; b_exp3 = 10'd282;
a_sign0 = 4'd11; a_sign1 = 4'd9; a_sign2 = 4'd6; a_sign3 = 4'd7;
b_sign0 = 4'd15; b_sign1 = 4'd10; b_sign2 = 4'd14; b_sign3 = 4'd1;
@(posedge clk_i);
a_mant0 = 8'd237; a_mant1 = 8'd98; a_mant2 = 8'd38; a_mant3 = 8'd66;
b_mant0 = 8'd37; b_mant1 = 8'd249; b_mant2 = 8'd200; b_mant3 = 8'd99;
a_exp0 = 10'd510; a_exp1 = 10'd974; a_exp2 = 10'd788; a_exp3 = 10'd209;
b_exp0 = 10'd56; b_exp1 = 10'd0; b_exp2 = 10'd111; b_exp3 = 10'd945;
a_sign0 = 4'd2; a_sign1 = 4'd4; a_sign2 = 4'd1; a_sign3 = 4'd10;
b_sign0 = 4'd6; b_sign1 = 4'd2; b_sign2 = 4'd16; b_sign3 = 4'd6;
@(posedge clk_i);
a_mant0 = 8'd88; a_mant1 = 8'd133; a_mant2 = 8'd241; a_mant3 = 8'd245;
b_mant0 = 8'd90; b_mant1 = 8'd244; b_mant2 = 8'd94; b_mant3 = 8'd200;
a_exp0 = 10'd856; a_exp1 = 10'd88; a_exp2 = 10'd742; a_exp3 = 10'd851;
b_exp0 = 10'd894; b_exp1 = 10'd334; b_exp2 = 10'd563; b_exp3 = 10'd362;
a_sign0 = 4'd4; a_sign1 = 4'd9; a_sign2 = 4'd9; a_sign3 = 4'd16;
b_sign0 = 4'd2; b_sign1 = 4'd2; b_sign2 = 4'd9; b_sign3 = 4'd9;
@(posedge clk_i);
a_mant0 = 8'd72; a_mant1 = 8'd162; a_mant2 = 8'd79; a_mant3 = 8'd116;
b_mant0 = 8'd88; b_mant1 = 8'd239; b_mant2 = 8'd46; b_mant3 = 8'd44;
a_exp0 = 10'd571; a_exp1 = 10'd956; a_exp2 = 10'd654; a_exp3 = 10'd782;
b_exp0 = 10'd329; b_exp1 = 10'd653; b_exp2 = 10'd253; b_exp3 = 10'd1019;
a_sign0 = 4'd5; a_sign1 = 4'd10; a_sign2 = 4'd7; a_sign3 = 4'd2;
b_sign0 = 4'd0; b_sign1 = 4'd3; b_sign2 = 4'd10; b_sign3 = 4'd7;
@(posedge clk_i);
a_mant0 = 8'd87; a_mant1 = 8'd233; a_mant2 = 8'd33; a_mant3 = 8'd58;
b_mant0 = 8'd91; b_mant1 = 8'd39; b_mant2 = 8'd36; b_mant3 = 8'd146;
a_exp0 = 10'd686; a_exp1 = 10'd95; a_exp2 = 10'd969; a_exp3 = 10'd1007;
b_exp0 = 10'd492; b_exp1 = 10'd865; b_exp2 = 10'd112; b_exp3 = 10'd312;
a_sign0 = 4'd4; a_sign1 = 4'd15; a_sign2 = 4'd10; a_sign3 = 4'd3;
b_sign0 = 4'd12; b_sign1 = 4'd5; b_sign2 = 4'd16; b_sign3 = 4'd14;
@(posedge clk_i);
a_mant0 = 8'd239; a_mant1 = 8'd36; a_mant2 = 8'd16; a_mant3 = 8'd207;
b_mant0 = 8'd39; b_mant1 = 8'd18; b_mant2 = 8'd36; b_mant3 = 8'd133;
a_exp0 = 10'd564; a_exp1 = 10'd318; a_exp2 = 10'd116; a_exp3 = 10'd164;
b_exp0 = 10'd102; b_exp1 = 10'd684; b_exp2 = 10'd251; b_exp3 = 10'd932;
a_sign0 = 4'd13; a_sign1 = 4'd15; a_sign2 = 4'd16; a_sign3 = 4'd1;
b_sign0 = 4'd4; b_sign1 = 4'd10; b_sign2 = 4'd8; b_sign3 = 4'd1;
@(posedge clk_i);
a_mant0 = 8'd130; a_mant1 = 8'd180; a_mant2 = 8'd62; a_mant3 = 8'd158;
b_mant0 = 8'd195; b_mant1 = 8'd145; b_mant2 = 8'd223; b_mant3 = 8'd72;
a_exp0 = 10'd737; a_exp1 = 10'd111; a_exp2 = 10'd419; a_exp3 = 10'd618;
b_exp0 = 10'd370; b_exp1 = 10'd940; b_exp2 = 10'd67; b_exp3 = 10'd684;
a_sign0 = 4'd9; a_sign1 = 4'd3; a_sign2 = 4'd9; a_sign3 = 4'd7;
b_sign0 = 4'd14; b_sign1 = 4'd7; b_sign2 = 4'd3; b_sign3 = 4'd0;
@(posedge clk_i);
a_mant0 = 8'd188; a_mant1 = 8'd86; a_mant2 = 8'd6; a_mant3 = 8'd81;
b_mant0 = 8'd101; b_mant1 = 8'd160; b_mant2 = 8'd222; b_mant3 = 8'd251;
a_exp0 = 10'd303; a_exp1 = 10'd885; a_exp2 = 10'd955; a_exp3 = 10'd351;
b_exp0 = 10'd22; b_exp1 = 10'd65; b_exp2 = 10'd732; b_exp3 = 10'd377;
a_sign0 = 4'd8; a_sign1 = 4'd1; a_sign2 = 4'd1; a_sign3 = 4'd1;
b_sign0 = 4'd3; b_sign1 = 4'd14; b_sign2 = 4'd3; b_sign3 = 4'd10;
@(posedge clk_i);
shared_exps0 = 8'd121;
shared_exps1 = 8'd113;
a_mant0 = 8'd100; a_mant1 = 8'd193; a_mant2 = 8'd142; a_mant3 = 8'd29;
b_mant0 = 8'd214; b_mant1 = 8'd138; b_mant2 = 8'd72; b_mant3 = 8'd143;
a_exp0 = 10'd226; a_exp1 = 10'd244; a_exp2 = 10'd799; a_exp3 = 10'd58;
b_exp0 = 10'd767; b_exp1 = 10'd569; b_exp2 = 10'd581; b_exp3 = 10'd474;
a_sign0 = 4'd12; a_sign1 = 4'd7; a_sign2 = 4'd11; a_sign3 = 4'd11;
b_sign0 = 4'd0; b_sign1 = 4'd7; b_sign2 = 4'd15; b_sign3 = 4'd10;
@(posedge clk_i);
a_mant0 = 8'd165; a_mant1 = 8'd98; a_mant2 = 8'd165; a_mant3 = 8'd54;
b_mant0 = 8'd239; b_mant1 = 8'd161; b_mant2 = 8'd99; b_mant3 = 8'd234;
a_exp0 = 10'd211; a_exp1 = 10'd537; a_exp2 = 10'd337; a_exp3 = 10'd916;
b_exp0 = 10'd795; b_exp1 = 10'd850; b_exp2 = 10'd855; b_exp3 = 10'd377;
a_sign0 = 4'd8; a_sign1 = 4'd14; a_sign2 = 4'd9; a_sign3 = 4'd6;
b_sign0 = 4'd11; b_sign1 = 4'd15; b_sign2 = 4'd7; b_sign3 = 4'd2;
@(posedge clk_i);
a_mant0 = 8'd8; a_mant1 = 8'd57; a_mant2 = 8'd118; a_mant3 = 8'd109;
b_mant0 = 8'd239; b_mant1 = 8'd189; b_mant2 = 8'd194; b_mant3 = 8'd225;
a_exp0 = 10'd201; a_exp1 = 10'd561; a_exp2 = 10'd127; a_exp3 = 10'd838;
b_exp0 = 10'd92; b_exp1 = 10'd926; b_exp2 = 10'd75; b_exp3 = 10'd500;
a_sign0 = 4'd11; a_sign1 = 4'd0; a_sign2 = 4'd4; a_sign3 = 4'd6;
b_sign0 = 4'd8; b_sign1 = 4'd1; b_sign2 = 4'd14; b_sign3 = 4'd10;
@(posedge clk_i);
a_mant0 = 8'd223; a_mant1 = 8'd4; a_mant2 = 8'd154; a_mant3 = 8'd54;
b_mant0 = 8'd99; b_mant1 = 8'd212; b_mant2 = 8'd250; b_mant3 = 8'd99;
a_exp0 = 10'd30; a_exp1 = 10'd632; a_exp2 = 10'd329; a_exp3 = 10'd871;
b_exp0 = 10'd847; b_exp1 = 10'd983; b_exp2 = 10'd202; b_exp3 = 10'd261;
a_sign0 = 4'd0; a_sign1 = 4'd5; a_sign2 = 4'd5; a_sign3 = 4'd5;
b_sign0 = 4'd4; b_sign1 = 4'd10; b_sign2 = 4'd6; b_sign3 = 4'd3;
@(posedge clk_i);
a_mant0 = 8'd131; a_mant1 = 8'd64; a_mant2 = 8'd247; a_mant3 = 8'd218;
b_mant0 = 8'd79; b_mant1 = 8'd141; b_mant2 = 8'd204; b_mant3 = 8'd222;
a_exp0 = 10'd483; a_exp1 = 10'd324; a_exp2 = 10'd83; a_exp3 = 10'd775;
b_exp0 = 10'd555; b_exp1 = 10'd169; b_exp2 = 10'd489; b_exp3 = 10'd958;
a_sign0 = 4'd12; a_sign1 = 4'd9; a_sign2 = 4'd12; a_sign3 = 4'd14;
b_sign0 = 4'd14; b_sign1 = 4'd8; b_sign2 = 4'd15; b_sign3 = 4'd13;
@(posedge clk_i);
a_mant0 = 8'd47; a_mant1 = 8'd146; a_mant2 = 8'd148; a_mant3 = 8'd155;
b_mant0 = 8'd182; b_mant1 = 8'd236; b_mant2 = 8'd37; b_mant3 = 8'd161;
a_exp0 = 10'd105; a_exp1 = 10'd643; a_exp2 = 10'd229; a_exp3 = 10'd560;
b_exp0 = 10'd661; b_exp1 = 10'd635; b_exp2 = 10'd716; b_exp3 = 10'd149;
a_sign0 = 4'd7; a_sign1 = 4'd9; a_sign2 = 4'd14; a_sign3 = 4'd5;
b_sign0 = 4'd10; b_sign1 = 4'd1; b_sign2 = 4'd13; b_sign3 = 4'd0;
@(posedge clk_i);
a_mant0 = 8'd49; a_mant1 = 8'd214; a_mant2 = 8'd205; a_mant3 = 8'd204;
b_mant0 = 8'd213; b_mant1 = 8'd158; b_mant2 = 8'd193; b_mant3 = 8'd133;
a_exp0 = 10'd471; a_exp1 = 10'd761; a_exp2 = 10'd875; a_exp3 = 10'd451;
b_exp0 = 10'd950; b_exp1 = 10'd1021; b_exp2 = 10'd66; b_exp3 = 10'd377;
a_sign0 = 4'd4; a_sign1 = 4'd4; a_sign2 = 4'd1; a_sign3 = 4'd4;
b_sign0 = 4'd7; b_sign1 = 4'd16; b_sign2 = 4'd11; b_sign3 = 4'd3;
@(posedge clk_i);
a_mant0 = 8'd153; a_mant1 = 8'd213; a_mant2 = 8'd130; a_mant3 = 8'd77;
b_mant0 = 8'd76; b_mant1 = 8'd135; b_mant2 = 8'd2; b_mant3 = 8'd210;
a_exp0 = 10'd802; a_exp1 = 10'd930; a_exp2 = 10'd224; a_exp3 = 10'd309;
b_exp0 = 10'd1015; b_exp1 = 10'd791; b_exp2 = 10'd862; b_exp3 = 10'd908;
a_sign0 = 4'd15; a_sign1 = 4'd5; a_sign2 = 4'd0; a_sign3 = 4'd2;
b_sign0 = 4'd6; b_sign1 = 4'd15; b_sign2 = 4'd15; b_sign3 = 4'd4;
@(posedge clk_i);
shared_exps0 = 8'd130;
shared_exps1 = 8'd128;
a_mant0 = 8'd71; a_mant1 = 8'd63; a_mant2 = 8'd156; a_mant3 = 8'd148;
b_mant0 = 8'd129; b_mant1 = 8'd123; b_mant2 = 8'd84; b_mant3 = 8'd201;
a_exp0 = 10'd825; a_exp1 = 10'd891; a_exp2 = 10'd569; a_exp3 = 10'd126;
b_exp0 = 10'd602; b_exp1 = 10'd552; b_exp2 = 10'd22; b_exp3 = 10'd210;
a_sign0 = 4'd14; a_sign1 = 4'd5; a_sign2 = 4'd16; a_sign3 = 4'd7;
b_sign0 = 4'd14; b_sign1 = 4'd11; b_sign2 = 4'd1; b_sign3 = 4'd12;
@(posedge clk_i);
a_mant0 = 8'd25; a_mant1 = 8'd93; a_mant2 = 8'd59; a_mant3 = 8'd233;
b_mant0 = 8'd101; b_mant1 = 8'd108; b_mant2 = 8'd13; b_mant3 = 8'd103;
a_exp0 = 10'd235; a_exp1 = 10'd775; a_exp2 = 10'd544; a_exp3 = 10'd864;
b_exp0 = 10'd850; b_exp1 = 10'd586; b_exp2 = 10'd409; b_exp3 = 10'd730;
a_sign0 = 4'd1; a_sign1 = 4'd5; a_sign2 = 4'd3; a_sign3 = 4'd5;
b_sign0 = 4'd14; b_sign1 = 4'd4; b_sign2 = 4'd1; b_sign3 = 4'd8;
@(posedge clk_i);
a_mant0 = 8'd128; a_mant1 = 8'd239; a_mant2 = 8'd228; a_mant3 = 8'd129;
b_mant0 = 8'd96; b_mant1 = 8'd1; b_mant2 = 8'd42; b_mant3 = 8'd21;
a_exp0 = 10'd630; a_exp1 = 10'd493; a_exp2 = 10'd456; a_exp3 = 10'd321;
b_exp0 = 10'd136; b_exp1 = 10'd278; b_exp2 = 10'd250; b_exp3 = 10'd928;
a_sign0 = 4'd10; a_sign1 = 4'd9; a_sign2 = 4'd1; a_sign3 = 4'd13;
b_sign0 = 4'd0; b_sign1 = 4'd0; b_sign2 = 4'd4; b_sign3 = 4'd6;
@(posedge clk_i);
a_mant0 = 8'd227; a_mant1 = 8'd75; a_mant2 = 8'd47; a_mant3 = 8'd228;
b_mant0 = 8'd112; b_mant1 = 8'd149; b_mant2 = 8'd9; b_mant3 = 8'd255;
a_exp0 = 10'd266; a_exp1 = 10'd271; a_exp2 = 10'd86; a_exp3 = 10'd366;
b_exp0 = 10'd571; b_exp1 = 10'd829; b_exp2 = 10'd498; b_exp3 = 10'd392;
a_sign0 = 4'd11; a_sign1 = 4'd10; a_sign2 = 4'd11; a_sign3 = 4'd16;
b_sign0 = 4'd8; b_sign1 = 4'd10; b_sign2 = 4'd12; b_sign3 = 4'd5;
@(posedge clk_i);
a_mant0 = 8'd102; a_mant1 = 8'd237; a_mant2 = 8'd185; a_mant3 = 8'd29;
b_mant0 = 8'd167; b_mant1 = 8'd25; b_mant2 = 8'd24; b_mant3 = 8'd223;
a_exp0 = 10'd3; a_exp1 = 10'd620; a_exp2 = 10'd807; a_exp3 = 10'd665;
b_exp0 = 10'd858; b_exp1 = 10'd616; b_exp2 = 10'd607; b_exp3 = 10'd353;
a_sign0 = 4'd6; a_sign1 = 4'd0; a_sign2 = 4'd2; a_sign3 = 4'd15;
b_sign0 = 4'd9; b_sign1 = 4'd7; b_sign2 = 4'd5; b_sign3 = 4'd5;
@(posedge clk_i);
a_mant0 = 8'd25; a_mant1 = 8'd131; a_mant2 = 8'd129; a_mant3 = 8'd198;
b_mant0 = 8'd6; b_mant1 = 8'd161; b_mant2 = 8'd54; b_mant3 = 8'd68;
a_exp0 = 10'd823; a_exp1 = 10'd789; a_exp2 = 10'd1011; a_exp3 = 10'd78;
b_exp0 = 10'd781; b_exp1 = 10'd363; b_exp2 = 10'd311; b_exp3 = 10'd477;
a_sign0 = 4'd12; a_sign1 = 4'd6; a_sign2 = 4'd13; a_sign3 = 4'd12;
b_sign0 = 4'd12; b_sign1 = 4'd1; b_sign2 = 4'd12; b_sign3 = 4'd12;
@(posedge clk_i);
a_mant0 = 8'd211; a_mant1 = 8'd138; a_mant2 = 8'd252; a_mant3 = 8'd48;
b_mant0 = 8'd55; b_mant1 = 8'd204; b_mant2 = 8'd225; b_mant3 = 8'd77;
a_exp0 = 10'd817; a_exp1 = 10'd339; a_exp2 = 10'd1021; a_exp3 = 10'd628;
b_exp0 = 10'd551; b_exp1 = 10'd640; b_exp2 = 10'd206; b_exp3 = 10'd945;
a_sign0 = 4'd9; a_sign1 = 4'd5; a_sign2 = 4'd9; a_sign3 = 4'd8;
b_sign0 = 4'd4; b_sign1 = 4'd15; b_sign2 = 4'd9; b_sign3 = 4'd3;
@(posedge clk_i);
a_mant0 = 8'd107; a_mant1 = 8'd247; a_mant2 = 8'd7; a_mant3 = 8'd30;
b_mant0 = 8'd44; b_mant1 = 8'd189; b_mant2 = 8'd222; b_mant3 = 8'd37;
a_exp0 = 10'd797; a_exp1 = 10'd437; a_exp2 = 10'd785; a_exp3 = 10'd412;
b_exp0 = 10'd554; b_exp1 = 10'd23; b_exp2 = 10'd927; b_exp3 = 10'd842;
a_sign0 = 4'd1; a_sign1 = 4'd13; a_sign2 = 4'd7; a_sign3 = 4'd15;
b_sign0 = 4'd4; b_sign1 = 4'd14; b_sign2 = 4'd10; b_sign3 = 4'd10;
@(posedge clk_i);
shared_exps0 = 8'd131;
shared_exps1 = 8'd121;
rstn = 0;
@(posedge clk_i);
rstn = 1;
a_mant0 = 8'd212; a_mant1 = 8'd20; a_mant2 = 8'd241; a_mant3 = 8'd71;
b_mant0 = 8'd38; b_mant1 = 8'd139; b_mant2 = 8'd18; b_mant3 = 8'd143;
a_exp0 = 10'd751; a_exp1 = 10'd720; a_exp2 = 10'd567; a_exp3 = 10'd75;
b_exp0 = 10'd474; b_exp1 = 10'd706; b_exp2 = 10'd354; b_exp3 = 10'd103;
a_sign0 = 4'd12; a_sign1 = 4'd13; a_sign2 = 4'd10; a_sign3 = 4'd5;
b_sign0 = 4'd6; b_sign1 = 4'd9; b_sign2 = 4'd9; b_sign3 = 4'd4;
@(posedge clk_i);
a_mant0 = 8'd203; a_mant1 = 8'd191; a_mant2 = 8'd163; a_mant3 = 8'd158;
b_mant0 = 8'd216; b_mant1 = 8'd188; b_mant2 = 8'd59; b_mant3 = 8'd170;
a_exp0 = 10'd512; a_exp1 = 10'd252; a_exp2 = 10'd310; a_exp3 = 10'd973;
b_exp0 = 10'd281; b_exp1 = 10'd507; b_exp2 = 10'd996; b_exp3 = 10'd386;
a_sign0 = 4'd1; a_sign1 = 4'd16; a_sign2 = 4'd5; a_sign3 = 4'd8;
b_sign0 = 4'd10; b_sign1 = 4'd4; b_sign2 = 4'd12; b_sign3 = 4'd9;
@(posedge clk_i);
a_mant0 = 8'd45; a_mant1 = 8'd110; a_mant2 = 8'd206; a_mant3 = 8'd71;
b_mant0 = 8'd69; b_mant1 = 8'd131; b_mant2 = 8'd160; b_mant3 = 8'd23;
a_exp0 = 10'd183; a_exp1 = 10'd142; a_exp2 = 10'd845; a_exp3 = 10'd584;
b_exp0 = 10'd796; b_exp1 = 10'd27; b_exp2 = 10'd85; b_exp3 = 10'd3;
a_sign0 = 4'd5; a_sign1 = 4'd16; a_sign2 = 4'd14; a_sign3 = 4'd3;
b_sign0 = 4'd2; b_sign1 = 4'd1; b_sign2 = 4'd9; b_sign3 = 4'd2;
@(posedge clk_i);
a_mant0 = 8'd7; a_mant1 = 8'd160; a_mant2 = 8'd126; a_mant3 = 8'd66;
b_mant0 = 8'd203; b_mant1 = 8'd63; b_mant2 = 8'd208; b_mant3 = 8'd22;
a_exp0 = 10'd940; a_exp1 = 10'd191; a_exp2 = 10'd972; a_exp3 = 10'd815;
b_exp0 = 10'd108; b_exp1 = 10'd686; b_exp2 = 10'd11; b_exp3 = 10'd80;
a_sign0 = 4'd13; a_sign1 = 4'd11; a_sign2 = 4'd1; a_sign3 = 4'd15;
b_sign0 = 4'd5; b_sign1 = 4'd16; b_sign2 = 4'd12; b_sign3 = 4'd0;
@(posedge clk_i);
a_mant0 = 8'd66; a_mant1 = 8'd133; a_mant2 = 8'd220; a_mant3 = 8'd0;
b_mant0 = 8'd244; b_mant1 = 8'd127; b_mant2 = 8'd117; b_mant3 = 8'd199;
a_exp0 = 10'd751; a_exp1 = 10'd431; a_exp2 = 10'd1001; a_exp3 = 10'd952;
b_exp0 = 10'd510; b_exp1 = 10'd377; b_exp2 = 10'd438; b_exp3 = 10'd202;
a_sign0 = 4'd8; a_sign1 = 4'd8; a_sign2 = 4'd5; a_sign3 = 4'd4;
b_sign0 = 4'd6; b_sign1 = 4'd6; b_sign2 = 4'd15; b_sign3 = 4'd13;
@(posedge clk_i);
a_mant0 = 8'd228; a_mant1 = 8'd1; a_mant2 = 8'd72; a_mant3 = 8'd19;
b_mant0 = 8'd101; b_mant1 = 8'd56; b_mant2 = 8'd108; b_mant3 = 8'd83;
a_exp0 = 10'd60; a_exp1 = 10'd733; a_exp2 = 10'd220; a_exp3 = 10'd845;
b_exp0 = 10'd703; b_exp1 = 10'd68; b_exp2 = 10'd105; b_exp3 = 10'd54;
a_sign0 = 4'd13; a_sign1 = 4'd12; a_sign2 = 4'd9; a_sign3 = 4'd4;
b_sign0 = 4'd9; b_sign1 = 4'd9; b_sign2 = 4'd9; b_sign3 = 4'd5;
@(posedge clk_i);
a_mant0 = 8'd48; a_mant1 = 8'd22; a_mant2 = 8'd125; a_mant3 = 8'd93;
b_mant0 = 8'd77; b_mant1 = 8'd7; b_mant2 = 8'd119; b_mant3 = 8'd251;
a_exp0 = 10'd683; a_exp1 = 10'd123; a_exp2 = 10'd660; a_exp3 = 10'd458;
b_exp0 = 10'd376; b_exp1 = 10'd230; b_exp2 = 10'd149; b_exp3 = 10'd839;
a_sign0 = 4'd4; a_sign1 = 4'd3; a_sign2 = 4'd12; a_sign3 = 4'd6;
b_sign0 = 4'd1; b_sign1 = 4'd3; b_sign2 = 4'd12; b_sign3 = 4'd9;
@(posedge clk_i);
shared_exps0 = 8'd135;
shared_exps1 = 8'd119;
a_mant0 = 8'd174; a_mant1 = 8'd80; a_mant2 = 8'd146; a_mant3 = 8'd83;
b_mant0 = 8'd186; b_mant1 = 8'd47; b_mant2 = 8'd179; b_mant3 = 8'd57;
a_exp0 = 10'd998; a_exp1 = 10'd885; a_exp2 = 10'd286; a_exp3 = 10'd312;
b_exp0 = 10'd677; b_exp1 = 10'd264; b_exp2 = 10'd849; b_exp3 = 10'd50;
a_sign0 = 4'd12; a_sign1 = 4'd0; a_sign2 = 4'd9; a_sign3 = 4'd4;
b_sign0 = 4'd11; b_sign1 = 4'd10; b_sign2 = 4'd4; b_sign3 = 4'd2;
@(posedge clk_i);
a_mant0 = 8'd50; a_mant1 = 8'd37; a_mant2 = 8'd191; a_mant3 = 8'd78;
b_mant0 = 8'd21; b_mant1 = 8'd121; b_mant2 = 8'd39; b_mant3 = 8'd197;
a_exp0 = 10'd495; a_exp1 = 10'd355; a_exp2 = 10'd372; a_exp3 = 10'd623;
b_exp0 = 10'd130; b_exp1 = 10'd389; b_exp2 = 10'd162; b_exp3 = 10'd66;
a_sign0 = 4'd4; a_sign1 = 4'd15; a_sign2 = 4'd10; a_sign3 = 4'd10;
b_sign0 = 4'd16; b_sign1 = 4'd14; b_sign2 = 4'd15; b_sign3 = 4'd14;
@(posedge clk_i);
a_mant0 = 8'd109; a_mant1 = 8'd112; a_mant2 = 8'd98; a_mant3 = 8'd105;
b_mant0 = 8'd117; b_mant1 = 8'd87; b_mant2 = 8'd205; b_mant3 = 8'd18;
a_exp0 = 10'd15; a_exp1 = 10'd184; a_exp2 = 10'd403; a_exp3 = 10'd95;
b_exp0 = 10'd195; b_exp1 = 10'd545; b_exp2 = 10'd318; b_exp3 = 10'd148;
a_sign0 = 4'd5; a_sign1 = 4'd10; a_sign2 = 4'd9; a_sign3 = 4'd8;
b_sign0 = 4'd6; b_sign1 = 4'd13; b_sign2 = 4'd16; b_sign3 = 4'd4;
@(posedge clk_i);
a_mant0 = 8'd248; a_mant1 = 8'd210; a_mant2 = 8'd66; a_mant3 = 8'd4;
b_mant0 = 8'd214; b_mant1 = 8'd58; b_mant2 = 8'd26; b_mant3 = 8'd143;
a_exp0 = 10'd233; a_exp1 = 10'd983; a_exp2 = 10'd614; a_exp3 = 10'd913;
b_exp0 = 10'd666; b_exp1 = 10'd661; b_exp2 = 10'd747; b_exp3 = 10'd322;
a_sign0 = 4'd9; a_sign1 = 4'd3; a_sign2 = 4'd5; a_sign3 = 4'd10;
b_sign0 = 4'd1; b_sign1 = 4'd13; b_sign2 = 4'd13; b_sign3 = 4'd11;
@(posedge clk_i);
a_mant0 = 8'd191; a_mant1 = 8'd129; a_mant2 = 8'd200; a_mant3 = 8'd29;
b_mant0 = 8'd111; b_mant1 = 8'd141; b_mant2 = 8'd244; b_mant3 = 8'd240;
a_exp0 = 10'd87; a_exp1 = 10'd665; a_exp2 = 10'd64; a_exp3 = 10'd1008;
b_exp0 = 10'd264; b_exp1 = 10'd407; b_exp2 = 10'd100; b_exp3 = 10'd1009;
a_sign0 = 4'd4; a_sign1 = 4'd13; a_sign2 = 4'd1; a_sign3 = 4'd14;
b_sign0 = 4'd14; b_sign1 = 4'd7; b_sign2 = 4'd6; b_sign3 = 4'd12;
@(posedge clk_i);
a_mant0 = 8'd9; a_mant1 = 8'd43; a_mant2 = 8'd14; a_mant3 = 8'd56;
b_mant0 = 8'd170; b_mant1 = 8'd204; b_mant2 = 8'd43; b_mant3 = 8'd190;
a_exp0 = 10'd395; a_exp1 = 10'd1013; a_exp2 = 10'd830; a_exp3 = 10'd96;
b_exp0 = 10'd144; b_exp1 = 10'd609; b_exp2 = 10'd514; b_exp3 = 10'd374;
a_sign0 = 4'd6; a_sign1 = 4'd1; a_sign2 = 4'd2; a_sign3 = 4'd7;
b_sign0 = 4'd14; b_sign1 = 4'd11; b_sign2 = 4'd0; b_sign3 = 4'd13;
@(posedge clk_i);
a_mant0 = 8'd148; a_mant1 = 8'd40; a_mant2 = 8'd95; a_mant3 = 8'd35;
b_mant0 = 8'd16; b_mant1 = 8'd60; b_mant2 = 8'd31; b_mant3 = 8'd89;
a_exp0 = 10'd964; a_exp1 = 10'd19; a_exp2 = 10'd626; a_exp3 = 10'd5;
b_exp0 = 10'd475; b_exp1 = 10'd732; b_exp2 = 10'd647; b_exp3 = 10'd280;
a_sign0 = 4'd9; a_sign1 = 4'd12; a_sign2 = 4'd8; a_sign3 = 4'd0;
b_sign0 = 4'd6; b_sign1 = 4'd6; b_sign2 = 4'd2; b_sign3 = 4'd9;
@(posedge clk_i);
a_mant0 = 8'd235; a_mant1 = 8'd111; a_mant2 = 8'd48; a_mant3 = 8'd13;
b_mant0 = 8'd127; b_mant1 = 8'd123; b_mant2 = 8'd173; b_mant3 = 8'd74;
a_exp0 = 10'd532; a_exp1 = 10'd368; a_exp2 = 10'd170; a_exp3 = 10'd387;
b_exp0 = 10'd594; b_exp1 = 10'd366; b_exp2 = 10'd578; b_exp3 = 10'd99;
a_sign0 = 4'd15; a_sign1 = 4'd16; a_sign2 = 4'd11; a_sign3 = 4'd4;
b_sign0 = 4'd4; b_sign1 = 4'd12; b_sign2 = 4'd16; b_sign3 = 4'd8;
@(posedge clk_i);
shared_exps0 = 8'd143;
shared_exps1 = 8'd115;
a_mant0 = 8'd163; a_mant1 = 8'd203; a_mant2 = 8'd138; a_mant3 = 8'd204;
b_mant0 = 8'd119; b_mant1 = 8'd229; b_mant2 = 8'd162; b_mant3 = 8'd87;
a_exp0 = 10'd644; a_exp1 = 10'd533; a_exp2 = 10'd853; a_exp3 = 10'd484;
b_exp0 = 10'd303; b_exp1 = 10'd91; b_exp2 = 10'd879; b_exp3 = 10'd853;
a_sign0 = 4'd9; a_sign1 = 4'd4; a_sign2 = 4'd13; a_sign3 = 4'd8;
b_sign0 = 4'd12; b_sign1 = 4'd14; b_sign2 = 4'd16; b_sign3 = 4'd8;
@(posedge clk_i);
a_mant0 = 8'd141; a_mant1 = 8'd39; a_mant2 = 8'd132; a_mant3 = 8'd146;
b_mant0 = 8'd148; b_mant1 = 8'd138; b_mant2 = 8'd72; b_mant3 = 8'd48;
a_exp0 = 10'd633; a_exp1 = 10'd106; a_exp2 = 10'd997; a_exp3 = 10'd380;
b_exp0 = 10'd929; b_exp1 = 10'd253; b_exp2 = 10'd349; b_exp3 = 10'd864;
a_sign0 = 4'd11; a_sign1 = 4'd12; a_sign2 = 4'd15; a_sign3 = 4'd5;
b_sign0 = 4'd1; b_sign1 = 4'd4; b_sign2 = 4'd9; b_sign3 = 4'd0;
@(posedge clk_i);
a_mant0 = 8'd224; a_mant1 = 8'd171; a_mant2 = 8'd193; a_mant3 = 8'd207;
b_mant0 = 8'd212; b_mant1 = 8'd50; b_mant2 = 8'd98; b_mant3 = 8'd96;
a_exp0 = 10'd365; a_exp1 = 10'd152; a_exp2 = 10'd878; a_exp3 = 10'd200;
b_exp0 = 10'd893; b_exp1 = 10'd515; b_exp2 = 10'd50; b_exp3 = 10'd952;
a_sign0 = 4'd9; a_sign1 = 4'd4; a_sign2 = 4'd5; a_sign3 = 4'd2;
b_sign0 = 4'd16; b_sign1 = 4'd9; b_sign2 = 4'd5; b_sign3 = 4'd8;
@(posedge clk_i);
a_mant0 = 8'd56; a_mant1 = 8'd152; a_mant2 = 8'd140; a_mant3 = 8'd74;
b_mant0 = 8'd149; b_mant1 = 8'd215; b_mant2 = 8'd197; b_mant3 = 8'd149;
a_exp0 = 10'd683; a_exp1 = 10'd834; a_exp2 = 10'd987; a_exp3 = 10'd159;
b_exp0 = 10'd948; b_exp1 = 10'd290; b_exp2 = 10'd788; b_exp3 = 10'd988;
a_sign0 = 4'd15; a_sign1 = 4'd10; a_sign2 = 4'd14; a_sign3 = 4'd0;
b_sign0 = 4'd12; b_sign1 = 4'd12; b_sign2 = 4'd5; b_sign3 = 4'd1;
@(posedge clk_i);
a_mant0 = 8'd76; a_mant1 = 8'd206; a_mant2 = 8'd117; a_mant3 = 8'd177;
b_mant0 = 8'd202; b_mant1 = 8'd173; b_mant2 = 8'd206; b_mant3 = 8'd31;
a_exp0 = 10'd662; a_exp1 = 10'd6; a_exp2 = 10'd246; a_exp3 = 10'd928;
b_exp0 = 10'd66; b_exp1 = 10'd1018; b_exp2 = 10'd374; b_exp3 = 10'd868;
a_sign0 = 4'd3; a_sign1 = 4'd12; a_sign2 = 4'd3; a_sign3 = 4'd16;
b_sign0 = 4'd1; b_sign1 = 4'd7; b_sign2 = 4'd12; b_sign3 = 4'd2;
@(posedge clk_i);
a_mant0 = 8'd50; a_mant1 = 8'd165; a_mant2 = 8'd42; a_mant3 = 8'd27;
b_mant0 = 8'd182; b_mant1 = 8'd197; b_mant2 = 8'd122; b_mant3 = 8'd55;
a_exp0 = 10'd168; a_exp1 = 10'd647; a_exp2 = 10'd637; a_exp3 = 10'd268;
b_exp0 = 10'd905; b_exp1 = 10'd94; b_exp2 = 10'd51; b_exp3 = 10'd556;
a_sign0 = 4'd6; a_sign1 = 4'd6; a_sign2 = 4'd13; a_sign3 = 4'd11;
b_sign0 = 4'd8; b_sign1 = 4'd8; b_sign2 = 4'd11; b_sign3 = 4'd12;
@(posedge clk_i);
a_mant0 = 8'd12; a_mant1 = 8'd236; a_mant2 = 8'd35; a_mant3 = 8'd84;
b_mant0 = 8'd253; b_mant1 = 8'd251; b_mant2 = 8'd11; b_mant3 = 8'd103;
a_exp0 = 10'd362; a_exp1 = 10'd425; a_exp2 = 10'd379; a_exp3 = 10'd143;
b_exp0 = 10'd587; b_exp1 = 10'd611; b_exp2 = 10'd844; b_exp3 = 10'd824;
a_sign0 = 4'd8; a_sign1 = 4'd5; a_sign2 = 4'd1; a_sign3 = 4'd8;
b_sign0 = 4'd11; b_sign1 = 4'd0; b_sign2 = 4'd13; b_sign3 = 4'd4;
@(posedge clk_i);
a_mant0 = 8'd69; a_mant1 = 8'd211; a_mant2 = 8'd105; a_mant3 = 8'd90;
b_mant0 = 8'd43; b_mant1 = 8'd242; b_mant2 = 8'd29; b_mant3 = 8'd133;
a_exp0 = 10'd563; a_exp1 = 10'd317; a_exp2 = 10'd786; a_exp3 = 10'd294;
b_exp0 = 10'd687; b_exp1 = 10'd642; b_exp2 = 10'd686; b_exp3 = 10'd160;
a_sign0 = 4'd16; a_sign1 = 4'd6; a_sign2 = 4'd4; a_sign3 = 4'd3;
b_sign0 = 4'd0; b_sign1 = 4'd9; b_sign2 = 4'd0; b_sign3 = 4'd3;
@(posedge clk_i);
shared_exps0 = 8'd129;
shared_exps1 = 8'd130;
a_mant0 = 8'd203; a_mant1 = 8'd174; a_mant2 = 8'd189; a_mant3 = 8'd92;
b_mant0 = 8'd213; b_mant1 = 8'd52; b_mant2 = 8'd69; b_mant3 = 8'd22;
a_exp0 = 10'd137; a_exp1 = 10'd755; a_exp2 = 10'd238; a_exp3 = 10'd1000;
b_exp0 = 10'd292; b_exp1 = 10'd525; b_exp2 = 10'd618; b_exp3 = 10'd324;
a_sign0 = 4'd5; a_sign1 = 4'd12; a_sign2 = 4'd11; a_sign3 = 4'd2;
b_sign0 = 4'd9; b_sign1 = 4'd8; b_sign2 = 4'd16; b_sign3 = 4'd10;
@(posedge clk_i);
a_mant0 = 8'd160; a_mant1 = 8'd131; a_mant2 = 8'd167; a_mant3 = 8'd193;
b_mant0 = 8'd33; b_mant1 = 8'd5; b_mant2 = 8'd38; b_mant3 = 8'd220;
a_exp0 = 10'd862; a_exp1 = 10'd26; a_exp2 = 10'd201; a_exp3 = 10'd109;
b_exp0 = 10'd84; b_exp1 = 10'd169; b_exp2 = 10'd704; b_exp3 = 10'd629;
a_sign0 = 4'd0; a_sign1 = 4'd12; a_sign2 = 4'd11; a_sign3 = 4'd16;
b_sign0 = 4'd11; b_sign1 = 4'd3; b_sign2 = 4'd2; b_sign3 = 4'd12;
@(posedge clk_i);
a_mant0 = 8'd65; a_mant1 = 8'd53; a_mant2 = 8'd191; a_mant3 = 8'd124;
b_mant0 = 8'd58; b_mant1 = 8'd192; b_mant2 = 8'd23; b_mant3 = 8'd29;
a_exp0 = 10'd982; a_exp1 = 10'd963; a_exp2 = 10'd29; a_exp3 = 10'd729;
b_exp0 = 10'd821; b_exp1 = 10'd499; b_exp2 = 10'd378; b_exp3 = 10'd580;
a_sign0 = 4'd15; a_sign1 = 4'd15; a_sign2 = 4'd15; a_sign3 = 4'd16;
b_sign0 = 4'd10; b_sign1 = 4'd0; b_sign2 = 4'd5; b_sign3 = 4'd9;
@(posedge clk_i);
a_mant0 = 8'd220; a_mant1 = 8'd113; a_mant2 = 8'd136; a_mant3 = 8'd253;
b_mant0 = 8'd46; b_mant1 = 8'd119; b_mant2 = 8'd91; b_mant3 = 8'd44;
a_exp0 = 10'd33; a_exp1 = 10'd960; a_exp2 = 10'd507; a_exp3 = 10'd699;
b_exp0 = 10'd483; b_exp1 = 10'd267; b_exp2 = 10'd212; b_exp3 = 10'd307;
a_sign0 = 4'd7; a_sign1 = 4'd0; a_sign2 = 4'd2; a_sign3 = 4'd3;
b_sign0 = 4'd3; b_sign1 = 4'd0; b_sign2 = 4'd6; b_sign3 = 4'd10;
@(posedge clk_i);
a_mant0 = 8'd66; a_mant1 = 8'd136; a_mant2 = 8'd197; a_mant3 = 8'd139;
b_mant0 = 8'd185; b_mant1 = 8'd211; b_mant2 = 8'd143; b_mant3 = 8'd246;
a_exp0 = 10'd210; a_exp1 = 10'd872; a_exp2 = 10'd321; a_exp3 = 10'd354;
b_exp0 = 10'd799; b_exp1 = 10'd700; b_exp2 = 10'd947; b_exp3 = 10'd885;
a_sign0 = 4'd7; a_sign1 = 4'd16; a_sign2 = 4'd2; a_sign3 = 4'd11;
b_sign0 = 4'd5; b_sign1 = 4'd14; b_sign2 = 4'd12; b_sign3 = 4'd14;
@(posedge clk_i);
a_mant0 = 8'd28; a_mant1 = 8'd140; a_mant2 = 8'd188; a_mant3 = 8'd77;
b_mant0 = 8'd18; b_mant1 = 8'd7; b_mant2 = 8'd91; b_mant3 = 8'd241;
a_exp0 = 10'd219; a_exp1 = 10'd694; a_exp2 = 10'd869; a_exp3 = 10'd314;
b_exp0 = 10'd13; b_exp1 = 10'd42; b_exp2 = 10'd122; b_exp3 = 10'd831;
a_sign0 = 4'd9; a_sign1 = 4'd0; a_sign2 = 4'd7; a_sign3 = 4'd8;
b_sign0 = 4'd13; b_sign1 = 4'd1; b_sign2 = 4'd1; b_sign3 = 4'd10;
@(posedge clk_i);
a_mant0 = 8'd157; a_mant1 = 8'd248; a_mant2 = 8'd24; a_mant3 = 8'd173;
b_mant0 = 8'd103; b_mant1 = 8'd98; b_mant2 = 8'd203; b_mant3 = 8'd7;
a_exp0 = 10'd235; a_exp1 = 10'd578; a_exp2 = 10'd629; a_exp3 = 10'd888;
b_exp0 = 10'd203; b_exp1 = 10'd509; b_exp2 = 10'd59; b_exp3 = 10'd261;
a_sign0 = 4'd12; a_sign1 = 4'd8; a_sign2 = 4'd5; a_sign3 = 4'd2;
b_sign0 = 4'd13; b_sign1 = 4'd16; b_sign2 = 4'd6; b_sign3 = 4'd2;
@(posedge clk_i);
a_mant0 = 8'd44; a_mant1 = 8'd219; a_mant2 = 8'd171; a_mant3 = 8'd197;
b_mant0 = 8'd60; b_mant1 = 8'd253; b_mant2 = 8'd6; b_mant3 = 8'd23;
a_exp0 = 10'd615; a_exp1 = 10'd834; a_exp2 = 10'd657; a_exp3 = 10'd493;
b_exp0 = 10'd229; b_exp1 = 10'd734; b_exp2 = 10'd241; b_exp3 = 10'd608;
a_sign0 = 4'd9; a_sign1 = 4'd15; a_sign2 = 4'd14; a_sign3 = 4'd7;
b_sign0 = 4'd3; b_sign1 = 4'd1; b_sign2 = 4'd6; b_sign3 = 4'd1;
@(posedge clk_i);
shared_exps0 = 8'd132;
shared_exps1 = 8'd111;
rstn = 0;
@(posedge clk_i);
rstn = 1;
a_mant0 = 8'd125; a_mant1 = 8'd102; a_mant2 = 8'd125; a_mant3 = 8'd145;
b_mant0 = 8'd134; b_mant1 = 8'd239; b_mant2 = 8'd118; b_mant3 = 8'd169;
a_exp0 = 10'd250; a_exp1 = 10'd170; a_exp2 = 10'd838; a_exp3 = 10'd54;
b_exp0 = 10'd880; b_exp1 = 10'd294; b_exp2 = 10'd909; b_exp3 = 10'd845;
a_sign0 = 4'd16; a_sign1 = 4'd12; a_sign2 = 4'd13; a_sign3 = 4'd14;
b_sign0 = 4'd16; b_sign1 = 4'd2; b_sign2 = 4'd13; b_sign3 = 4'd9;
@(posedge clk_i);
a_mant0 = 8'd89; a_mant1 = 8'd115; a_mant2 = 8'd33; a_mant3 = 8'd69;
b_mant0 = 8'd64; b_mant1 = 8'd53; b_mant2 = 8'd178; b_mant3 = 8'd152;
a_exp0 = 10'd459; a_exp1 = 10'd727; a_exp2 = 10'd574; a_exp3 = 10'd309;
b_exp0 = 10'd441; b_exp1 = 10'd966; b_exp2 = 10'd940; b_exp3 = 10'd985;
a_sign0 = 4'd15; a_sign1 = 4'd4; a_sign2 = 4'd12; a_sign3 = 4'd10;
b_sign0 = 4'd1; b_sign1 = 4'd12; b_sign2 = 4'd4; b_sign3 = 4'd0;
@(posedge clk_i);
a_mant0 = 8'd153; a_mant1 = 8'd150; a_mant2 = 8'd104; a_mant3 = 8'd89;
b_mant0 = 8'd167; b_mant1 = 8'd163; b_mant2 = 8'd235; b_mant3 = 8'd181;
a_exp0 = 10'd986; a_exp1 = 10'd72; a_exp2 = 10'd0; a_exp3 = 10'd1007;
b_exp0 = 10'd705; b_exp1 = 10'd856; b_exp2 = 10'd363; b_exp3 = 10'd757;
a_sign0 = 4'd6; a_sign1 = 4'd11; a_sign2 = 4'd12; a_sign3 = 4'd12;
b_sign0 = 4'd10; b_sign1 = 4'd2; b_sign2 = 4'd0; b_sign3 = 4'd8;
@(posedge clk_i);
a_mant0 = 8'd55; a_mant1 = 8'd45; a_mant2 = 8'd245; a_mant3 = 8'd61;
b_mant0 = 8'd73; b_mant1 = 8'd34; b_mant2 = 8'd8; b_mant3 = 8'd146;
a_exp0 = 10'd507; a_exp1 = 10'd248; a_exp2 = 10'd532; a_exp3 = 10'd88;
b_exp0 = 10'd553; b_exp1 = 10'd597; b_exp2 = 10'd249; b_exp3 = 10'd840;
a_sign0 = 4'd11; a_sign1 = 4'd1; a_sign2 = 4'd5; a_sign3 = 4'd15;
b_sign0 = 4'd7; b_sign1 = 4'd3; b_sign2 = 4'd6; b_sign3 = 4'd9;
@(posedge clk_i);
a_mant0 = 8'd234; a_mant1 = 8'd200; a_mant2 = 8'd148; a_mant3 = 8'd206;
b_mant0 = 8'd92; b_mant1 = 8'd195; b_mant2 = 8'd103; b_mant3 = 8'd226;
a_exp0 = 10'd33; a_exp1 = 10'd718; a_exp2 = 10'd1020; a_exp3 = 10'd79;
b_exp0 = 10'd104; b_exp1 = 10'd235; b_exp2 = 10'd123; b_exp3 = 10'd562;
a_sign0 = 4'd12; a_sign1 = 4'd15; a_sign2 = 4'd10; a_sign3 = 4'd16;
b_sign0 = 4'd15; b_sign1 = 4'd7; b_sign2 = 4'd5; b_sign3 = 4'd5;
@(posedge clk_i);
a_mant0 = 8'd212; a_mant1 = 8'd8; a_mant2 = 8'd189; a_mant3 = 8'd87;
b_mant0 = 8'd43; b_mant1 = 8'd140; b_mant2 = 8'd155; b_mant3 = 8'd158;
a_exp0 = 10'd969; a_exp1 = 10'd715; a_exp2 = 10'd850; a_exp3 = 10'd478;
b_exp0 = 10'd768; b_exp1 = 10'd925; b_exp2 = 10'd22; b_exp3 = 10'd105;
a_sign0 = 4'd9; a_sign1 = 4'd8; a_sign2 = 4'd3; a_sign3 = 4'd8;
b_sign0 = 4'd12; b_sign1 = 4'd12; b_sign2 = 4'd12; b_sign3 = 4'd0;
@(posedge clk_i);
a_mant0 = 8'd237; a_mant1 = 8'd144; a_mant2 = 8'd145; a_mant3 = 8'd223;
b_mant0 = 8'd153; b_mant1 = 8'd65; b_mant2 = 8'd136; b_mant3 = 8'd193;
a_exp0 = 10'd679; a_exp1 = 10'd139; a_exp2 = 10'd321; a_exp3 = 10'd565;
b_exp0 = 10'd674; b_exp1 = 10'd137; b_exp2 = 10'd650; b_exp3 = 10'd839;
a_sign0 = 4'd16; a_sign1 = 4'd9; a_sign2 = 4'd8; a_sign3 = 4'd14;
b_sign0 = 4'd9; b_sign1 = 4'd9; b_sign2 = 4'd6; b_sign3 = 4'd2;
@(posedge clk_i);
shared_exps0 = 8'd95;
shared_exps1 = 8'd121;
a_mant0 = 8'd29; a_mant1 = 8'd124; a_mant2 = 8'd205; a_mant3 = 8'd194;
b_mant0 = 8'd87; b_mant1 = 8'd102; b_mant2 = 8'd180; b_mant3 = 8'd162;
a_exp0 = 10'd201; a_exp1 = 10'd399; a_exp2 = 10'd54; a_exp3 = 10'd194;
b_exp0 = 10'd185; b_exp1 = 10'd807; b_exp2 = 10'd448; b_exp3 = 10'd747;
a_sign0 = 4'd1; a_sign1 = 4'd16; a_sign2 = 4'd6; a_sign3 = 4'd12;
b_sign0 = 4'd2; b_sign1 = 4'd8; b_sign2 = 4'd0; b_sign3 = 4'd15;
@(posedge clk_i);
a_mant0 = 8'd112; a_mant1 = 8'd112; a_mant2 = 8'd109; a_mant3 = 8'd147;
b_mant0 = 8'd223; b_mant1 = 8'd236; b_mant2 = 8'd230; b_mant3 = 8'd183;
a_exp0 = 10'd175; a_exp1 = 10'd508; a_exp2 = 10'd813; a_exp3 = 10'd552;
b_exp0 = 10'd651; b_exp1 = 10'd666; b_exp2 = 10'd858; b_exp3 = 10'd789;
a_sign0 = 4'd9; a_sign1 = 4'd3; a_sign2 = 4'd16; a_sign3 = 4'd7;
b_sign0 = 4'd1; b_sign1 = 4'd14; b_sign2 = 4'd12; b_sign3 = 4'd8;
@(posedge clk_i);
a_mant0 = 8'd92; a_mant1 = 8'd109; a_mant2 = 8'd131; a_mant3 = 8'd234;
b_mant0 = 8'd167; b_mant1 = 8'd214; b_mant2 = 8'd59; b_mant3 = 8'd65;
a_exp0 = 10'd400; a_exp1 = 10'd353; a_exp2 = 10'd296; a_exp3 = 10'd371;
b_exp0 = 10'd624; b_exp1 = 10'd635; b_exp2 = 10'd582; b_exp3 = 10'd567;
a_sign0 = 4'd1; a_sign1 = 4'd11; a_sign2 = 4'd11; a_sign3 = 4'd2;
b_sign0 = 4'd12; b_sign1 = 4'd10; b_sign2 = 4'd15; b_sign3 = 4'd4;
@(posedge clk_i);
a_mant0 = 8'd53; a_mant1 = 8'd101; a_mant2 = 8'd191; a_mant3 = 8'd132;
b_mant0 = 8'd3; b_mant1 = 8'd26; b_mant2 = 8'd134; b_mant3 = 8'd131;
a_exp0 = 10'd510; a_exp1 = 10'd941; a_exp2 = 10'd462; a_exp3 = 10'd78;
b_exp0 = 10'd622; b_exp1 = 10'd217; b_exp2 = 10'd963; b_exp3 = 10'd47;
a_sign0 = 4'd15; a_sign1 = 4'd11; a_sign2 = 4'd8; a_sign3 = 4'd12;
b_sign0 = 4'd9; b_sign1 = 4'd2; b_sign2 = 4'd5; b_sign3 = 4'd10;
@(posedge clk_i);
a_mant0 = 8'd200; a_mant1 = 8'd171; a_mant2 = 8'd127; a_mant3 = 8'd177;
b_mant0 = 8'd143; b_mant1 = 8'd6; b_mant2 = 8'd246; b_mant3 = 8'd236;
a_exp0 = 10'd543; a_exp1 = 10'd132; a_exp2 = 10'd205; a_exp3 = 10'd603;
b_exp0 = 10'd371; b_exp1 = 10'd287; b_exp2 = 10'd333; b_exp3 = 10'd978;
a_sign0 = 4'd1; a_sign1 = 4'd5; a_sign2 = 4'd7; a_sign3 = 4'd8;
b_sign0 = 4'd1; b_sign1 = 4'd10; b_sign2 = 4'd9; b_sign3 = 4'd0;
@(posedge clk_i);
a_mant0 = 8'd209; a_mant1 = 8'd53; a_mant2 = 8'd250; a_mant3 = 8'd139;
b_mant0 = 8'd238; b_mant1 = 8'd14; b_mant2 = 8'd115; b_mant3 = 8'd111;
a_exp0 = 10'd219; a_exp1 = 10'd667; a_exp2 = 10'd998; a_exp3 = 10'd299;
b_exp0 = 10'd776; b_exp1 = 10'd598; b_exp2 = 10'd231; b_exp3 = 10'd881;
a_sign0 = 4'd13; a_sign1 = 4'd5; a_sign2 = 4'd1; a_sign3 = 4'd8;
b_sign0 = 4'd0; b_sign1 = 4'd7; b_sign2 = 4'd2; b_sign3 = 4'd12;
@(posedge clk_i);
a_mant0 = 8'd242; a_mant1 = 8'd185; a_mant2 = 8'd110; a_mant3 = 8'd58;
b_mant0 = 8'd127; b_mant1 = 8'd207; b_mant2 = 8'd86; b_mant3 = 8'd31;
a_exp0 = 10'd327; a_exp1 = 10'd412; a_exp2 = 10'd835; a_exp3 = 10'd558;
b_exp0 = 10'd212; b_exp1 = 10'd390; b_exp2 = 10'd860; b_exp3 = 10'd138;
a_sign0 = 4'd3; a_sign1 = 4'd2; a_sign2 = 4'd4; a_sign3 = 4'd15;
b_sign0 = 4'd15; b_sign1 = 4'd0; b_sign2 = 4'd10; b_sign3 = 4'd4;
@(posedge clk_i);
a_mant0 = 8'd170; a_mant1 = 8'd140; a_mant2 = 8'd126; a_mant3 = 8'd45;
b_mant0 = 8'd57; b_mant1 = 8'd176; b_mant2 = 8'd192; b_mant3 = 8'd232;
a_exp0 = 10'd857; a_exp1 = 10'd151; a_exp2 = 10'd756; a_exp3 = 10'd165;
b_exp0 = 10'd910; b_exp1 = 10'd221; b_exp2 = 10'd126; b_exp3 = 10'd244;
a_sign0 = 4'd10; a_sign1 = 4'd4; a_sign2 = 4'd13; a_sign3 = 4'd15;
b_sign0 = 4'd0; b_sign1 = 4'd1; b_sign2 = 4'd0; b_sign3 = 4'd1;
@(posedge clk_i);
shared_exps0 = 8'd125;
shared_exps1 = 8'd112;
a_mant0 = 8'd196; a_mant1 = 8'd130; a_mant2 = 8'd5; a_mant3 = 8'd183;
b_mant0 = 8'd58; b_mant1 = 8'd224; b_mant2 = 8'd74; b_mant3 = 8'd34;
a_exp0 = 10'd299; a_exp1 = 10'd710; a_exp2 = 10'd647; a_exp3 = 10'd924;
b_exp0 = 10'd118; b_exp1 = 10'd421; b_exp2 = 10'd962; b_exp3 = 10'd254;
a_sign0 = 4'd2; a_sign1 = 4'd5; a_sign2 = 4'd13; a_sign3 = 4'd4;
b_sign0 = 4'd4; b_sign1 = 4'd14; b_sign2 = 4'd12; b_sign3 = 4'd3;
@(posedge clk_i);
a_mant0 = 8'd198; a_mant1 = 8'd83; a_mant2 = 8'd55; a_mant3 = 8'd47;
b_mant0 = 8'd8; b_mant1 = 8'd245; b_mant2 = 8'd188; b_mant3 = 8'd187;
a_exp0 = 10'd640; a_exp1 = 10'd740; a_exp2 = 10'd251; a_exp3 = 10'd913;
b_exp0 = 10'd119; b_exp1 = 10'd432; b_exp2 = 10'd833; b_exp3 = 10'd829;
a_sign0 = 4'd8; a_sign1 = 4'd8; a_sign2 = 4'd9; a_sign3 = 4'd9;
b_sign0 = 4'd10; b_sign1 = 4'd1; b_sign2 = 4'd4; b_sign3 = 4'd10;
@(posedge clk_i);
a_mant0 = 8'd141; a_mant1 = 8'd253; a_mant2 = 8'd89; a_mant3 = 8'd138;
b_mant0 = 8'd245; b_mant1 = 8'd69; b_mant2 = 8'd225; b_mant3 = 8'd214;
a_exp0 = 10'd148; a_exp1 = 10'd929; a_exp2 = 10'd978; a_exp3 = 10'd911;
b_exp0 = 10'd844; b_exp1 = 10'd616; b_exp2 = 10'd26; b_exp3 = 10'd705;
a_sign0 = 4'd6; a_sign1 = 4'd13; a_sign2 = 4'd7; a_sign3 = 4'd9;
b_sign0 = 4'd16; b_sign1 = 4'd8; b_sign2 = 4'd3; b_sign3 = 4'd16;
@(posedge clk_i);
a_mant0 = 8'd198; a_mant1 = 8'd129; a_mant2 = 8'd255; a_mant3 = 8'd54;
b_mant0 = 8'd32; b_mant1 = 8'd3; b_mant2 = 8'd220; b_mant3 = 8'd158;
a_exp0 = 10'd40; a_exp1 = 10'd105; a_exp2 = 10'd770; a_exp3 = 10'd819;
b_exp0 = 10'd60; b_exp1 = 10'd246; b_exp2 = 10'd390; b_exp3 = 10'd389;
a_sign0 = 4'd0; a_sign1 = 4'd6; a_sign2 = 4'd16; a_sign3 = 4'd4;
b_sign0 = 4'd6; b_sign1 = 4'd0; b_sign2 = 4'd14; b_sign3 = 4'd4;
@(posedge clk_i);
a_mant0 = 8'd149; a_mant1 = 8'd143; a_mant2 = 8'd231; a_mant3 = 8'd117;
b_mant0 = 8'd8; b_mant1 = 8'd45; b_mant2 = 8'd3; b_mant3 = 8'd147;
a_exp0 = 10'd92; a_exp1 = 10'd434; a_exp2 = 10'd969; a_exp3 = 10'd322;
b_exp0 = 10'd675; b_exp1 = 10'd503; b_exp2 = 10'd748; b_exp3 = 10'd799;
a_sign0 = 4'd3; a_sign1 = 4'd15; a_sign2 = 4'd12; a_sign3 = 4'd16;
b_sign0 = 4'd2; b_sign1 = 4'd3; b_sign2 = 4'd13; b_sign3 = 4'd8;
@(posedge clk_i);
a_mant0 = 8'd105; a_mant1 = 8'd70; a_mant2 = 8'd165; a_mant3 = 8'd227;
b_mant0 = 8'd168; b_mant1 = 8'd194; b_mant2 = 8'd36; b_mant3 = 8'd20;
a_exp0 = 10'd807; a_exp1 = 10'd487; a_exp2 = 10'd698; a_exp3 = 10'd347;
b_exp0 = 10'd582; b_exp1 = 10'd605; b_exp2 = 10'd243; b_exp3 = 10'd260;
a_sign0 = 4'd3; a_sign1 = 4'd6; a_sign2 = 4'd10; a_sign3 = 4'd13;
b_sign0 = 4'd15; b_sign1 = 4'd8; b_sign2 = 4'd8; b_sign3 = 4'd8;
@(posedge clk_i);
a_mant0 = 8'd57; a_mant1 = 8'd182; a_mant2 = 8'd13; a_mant3 = 8'd79;
b_mant0 = 8'd51; b_mant1 = 8'd140; b_mant2 = 8'd214; b_mant3 = 8'd220;
a_exp0 = 10'd141; a_exp1 = 10'd494; a_exp2 = 10'd8; a_exp3 = 10'd175;
b_exp0 = 10'd310; b_exp1 = 10'd785; b_exp2 = 10'd657; b_exp3 = 10'd954;
a_sign0 = 4'd0; a_sign1 = 4'd15; a_sign2 = 4'd12; a_sign3 = 4'd0;
b_sign0 = 4'd9; b_sign1 = 4'd14; b_sign2 = 4'd7; b_sign3 = 4'd1;
@(posedge clk_i);
a_mant0 = 8'd249; a_mant1 = 8'd47; a_mant2 = 8'd211; a_mant3 = 8'd136;
b_mant0 = 8'd51; b_mant1 = 8'd30; b_mant2 = 8'd249; b_mant3 = 8'd197;
a_exp0 = 10'd590; a_exp1 = 10'd258; a_exp2 = 10'd313; a_exp3 = 10'd512;
b_exp0 = 10'd93; b_exp1 = 10'd20; b_exp2 = 10'd440; b_exp3 = 10'd414;
a_sign0 = 4'd0; a_sign1 = 4'd2; a_sign2 = 4'd11; a_sign3 = 4'd13;
b_sign0 = 4'd9; b_sign1 = 4'd9; b_sign2 = 4'd14; b_sign3 = 4'd3;
@(posedge clk_i);
shared_exps0 = 8'd137;
shared_exps1 = 8'd140;
a_mant0 = 8'd84; a_mant1 = 8'd232; a_mant2 = 8'd20; a_mant3 = 8'd204;
b_mant0 = 8'd217; b_mant1 = 8'd123; b_mant2 = 8'd207; b_mant3 = 8'd246;
a_exp0 = 10'd988; a_exp1 = 10'd391; a_exp2 = 10'd414; a_exp3 = 10'd508;
b_exp0 = 10'd743; b_exp1 = 10'd100; b_exp2 = 10'd663; b_exp3 = 10'd615;
a_sign0 = 4'd15; a_sign1 = 4'd2; a_sign2 = 4'd0; a_sign3 = 4'd9;
b_sign0 = 4'd5; b_sign1 = 4'd2; b_sign2 = 4'd15; b_sign3 = 4'd16;
@(posedge clk_i);
a_mant0 = 8'd50; a_mant1 = 8'd165; a_mant2 = 8'd165; a_mant3 = 8'd183;
b_mant0 = 8'd213; b_mant1 = 8'd117; b_mant2 = 8'd237; b_mant3 = 8'd175;
a_exp0 = 10'd676; a_exp1 = 10'd578; a_exp2 = 10'd99; a_exp3 = 10'd354;
b_exp0 = 10'd38; b_exp1 = 10'd326; b_exp2 = 10'd7; b_exp3 = 10'd998;
a_sign0 = 4'd8; a_sign1 = 4'd15; a_sign2 = 4'd10; a_sign3 = 4'd1;
b_sign0 = 4'd9; b_sign1 = 4'd16; b_sign2 = 4'd12; b_sign3 = 4'd5;
@(posedge clk_i);
a_mant0 = 8'd243; a_mant1 = 8'd178; a_mant2 = 8'd200; a_mant3 = 8'd192;
b_mant0 = 8'd149; b_mant1 = 8'd216; b_mant2 = 8'd201; b_mant3 = 8'd240;
a_exp0 = 10'd279; a_exp1 = 10'd206; a_exp2 = 10'd887; a_exp3 = 10'd133;
b_exp0 = 10'd283; b_exp1 = 10'd419; b_exp2 = 10'd200; b_exp3 = 10'd442;
a_sign0 = 4'd8; a_sign1 = 4'd0; a_sign2 = 4'd4; a_sign3 = 4'd10;
b_sign0 = 4'd13; b_sign1 = 4'd13; b_sign2 = 4'd16; b_sign3 = 4'd0;
@(posedge clk_i);
a_mant0 = 8'd143; a_mant1 = 8'd36; a_mant2 = 8'd252; a_mant3 = 8'd146;
b_mant0 = 8'd223; b_mant1 = 8'd255; b_mant2 = 8'd225; b_mant3 = 8'd30;
a_exp0 = 10'd129; a_exp1 = 10'd929; a_exp2 = 10'd433; a_exp3 = 10'd91;
b_exp0 = 10'd676; b_exp1 = 10'd475; b_exp2 = 10'd569; b_exp3 = 10'd315;
a_sign0 = 4'd4; a_sign1 = 4'd1; a_sign2 = 4'd0; a_sign3 = 4'd14;
b_sign0 = 4'd16; b_sign1 = 4'd13; b_sign2 = 4'd6; b_sign3 = 4'd7;
@(posedge clk_i);
a_mant0 = 8'd151; a_mant1 = 8'd211; a_mant2 = 8'd243; a_mant3 = 8'd204;
b_mant0 = 8'd39; b_mant1 = 8'd136; b_mant2 = 8'd44; b_mant3 = 8'd250;
a_exp0 = 10'd440; a_exp1 = 10'd807; a_exp2 = 10'd870; a_exp3 = 10'd124;
b_exp0 = 10'd373; b_exp1 = 10'd659; b_exp2 = 10'd840; b_exp3 = 10'd623;
a_sign0 = 4'd10; a_sign1 = 4'd4; a_sign2 = 4'd14; a_sign3 = 4'd14;
b_sign0 = 4'd9; b_sign1 = 4'd9; b_sign2 = 4'd3; b_sign3 = 4'd12;
@(posedge clk_i);
a_mant0 = 8'd102; a_mant1 = 8'd203; a_mant2 = 8'd251; a_mant3 = 8'd36;
b_mant0 = 8'd55; b_mant1 = 8'd211; b_mant2 = 8'd100; b_mant3 = 8'd76;
a_exp0 = 10'd85; a_exp1 = 10'd354; a_exp2 = 10'd94; a_exp3 = 10'd986;
b_exp0 = 10'd551; b_exp1 = 10'd212; b_exp2 = 10'd447; b_exp3 = 10'd44;
a_sign0 = 4'd10; a_sign1 = 4'd13; a_sign2 = 4'd2; a_sign3 = 4'd11;
b_sign0 = 4'd4; b_sign1 = 4'd6; b_sign2 = 4'd12; b_sign3 = 4'd3;
@(posedge clk_i);
a_mant0 = 8'd76; a_mant1 = 8'd200; a_mant2 = 8'd59; a_mant3 = 8'd96;
b_mant0 = 8'd46; b_mant1 = 8'd134; b_mant2 = 8'd249; b_mant3 = 8'd197;
a_exp0 = 10'd748; a_exp1 = 10'd435; a_exp2 = 10'd66; a_exp3 = 10'd420;
b_exp0 = 10'd657; b_exp1 = 10'd348; b_exp2 = 10'd602; b_exp3 = 10'd225;
a_sign0 = 4'd9; a_sign1 = 4'd7; a_sign2 = 4'd13; a_sign3 = 4'd3;
b_sign0 = 4'd9; b_sign1 = 4'd13; b_sign2 = 4'd16; b_sign3 = 4'd9;
@(posedge clk_i);
a_mant0 = 8'd232; a_mant1 = 8'd20; a_mant2 = 8'd216; a_mant3 = 8'd57;
b_mant0 = 8'd51; b_mant1 = 8'd111; b_mant2 = 8'd158; b_mant3 = 8'd112;
a_exp0 = 10'd602; a_exp1 = 10'd376; a_exp2 = 10'd690; a_exp3 = 10'd229;
b_exp0 = 10'd434; b_exp1 = 10'd811; b_exp2 = 10'd223; b_exp3 = 10'd523;
a_sign0 = 4'd15; a_sign1 = 4'd14; a_sign2 = 4'd7; a_sign3 = 4'd15;
b_sign0 = 4'd1; b_sign1 = 4'd8; b_sign2 = 4'd10; b_sign3 = 4'd12;
@(posedge clk_i);
shared_exps0 = 8'd137;
shared_exps1 = 8'd114;
rstn = 0;
@(posedge clk_i);
rstn = 1;
a_mant0 = 8'd20; a_mant1 = 8'd13; a_mant2 = 8'd119; a_mant3 = 8'd233;
b_mant0 = 8'd116; b_mant1 = 8'd195; b_mant2 = 8'd177; b_mant3 = 8'd185;
a_exp0 = 10'd774; a_exp1 = 10'd385; a_exp2 = 10'd974; a_exp3 = 10'd11;
b_exp0 = 10'd951; b_exp1 = 10'd470; b_exp2 = 10'd73; b_exp3 = 10'd482;
a_sign0 = 4'd16; a_sign1 = 4'd3; a_sign2 = 4'd15; a_sign3 = 4'd11;
b_sign0 = 4'd12; b_sign1 = 4'd11; b_sign2 = 4'd15; b_sign3 = 4'd6;
@(posedge clk_i);
a_mant0 = 8'd35; a_mant1 = 8'd115; a_mant2 = 8'd240; a_mant3 = 8'd93;
b_mant0 = 8'd57; b_mant1 = 8'd237; b_mant2 = 8'd161; b_mant3 = 8'd78;
a_exp0 = 10'd10; a_exp1 = 10'd374; a_exp2 = 10'd557; a_exp3 = 10'd788;
b_exp0 = 10'd389; b_exp1 = 10'd229; b_exp2 = 10'd536; b_exp3 = 10'd196;
a_sign0 = 4'd14; a_sign1 = 4'd8; a_sign2 = 4'd10; a_sign3 = 4'd0;
b_sign0 = 4'd11; b_sign1 = 4'd13; b_sign2 = 4'd8; b_sign3 = 4'd12;
@(posedge clk_i);
a_mant0 = 8'd78; a_mant1 = 8'd216; a_mant2 = 8'd230; a_mant3 = 8'd141;
b_mant0 = 8'd183; b_mant1 = 8'd228; b_mant2 = 8'd202; b_mant3 = 8'd176;
a_exp0 = 10'd931; a_exp1 = 10'd544; a_exp2 = 10'd83; a_exp3 = 10'd689;
b_exp0 = 10'd829; b_exp1 = 10'd402; b_exp2 = 10'd85; b_exp3 = 10'd743;
a_sign0 = 4'd12; a_sign1 = 4'd7; a_sign2 = 4'd5; a_sign3 = 4'd10;
b_sign0 = 4'd7; b_sign1 = 4'd0; b_sign2 = 4'd1; b_sign3 = 4'd8;
@(posedge clk_i);
a_mant0 = 8'd180; a_mant1 = 8'd155; a_mant2 = 8'd98; a_mant3 = 8'd15;
b_mant0 = 8'd225; b_mant1 = 8'd178; b_mant2 = 8'd182; b_mant3 = 8'd168;
a_exp0 = 10'd206; a_exp1 = 10'd299; a_exp2 = 10'd311; a_exp3 = 10'd700;
b_exp0 = 10'd184; b_exp1 = 10'd167; b_exp2 = 10'd721; b_exp3 = 10'd437;
a_sign0 = 4'd12; a_sign1 = 4'd13; a_sign2 = 4'd14; a_sign3 = 4'd1;
b_sign0 = 4'd2; b_sign1 = 4'd13; b_sign2 = 4'd15; b_sign3 = 4'd14;
@(posedge clk_i);
a_mant0 = 8'd234; a_mant1 = 8'd145; a_mant2 = 8'd88; a_mant3 = 8'd203;
b_mant0 = 8'd218; b_mant1 = 8'd239; b_mant2 = 8'd90; b_mant3 = 8'd250;
a_exp0 = 10'd501; a_exp1 = 10'd615; a_exp2 = 10'd605; a_exp3 = 10'd902;
b_exp0 = 10'd293; b_exp1 = 10'd343; b_exp2 = 10'd225; b_exp3 = 10'd389;
a_sign0 = 4'd0; a_sign1 = 4'd12; a_sign2 = 4'd12; a_sign3 = 4'd4;
b_sign0 = 4'd4; b_sign1 = 4'd5; b_sign2 = 4'd3; b_sign3 = 4'd16;
@(posedge clk_i);
a_mant0 = 8'd182; a_mant1 = 8'd162; a_mant2 = 8'd75; a_mant3 = 8'd99;
b_mant0 = 8'd145; b_mant1 = 8'd109; b_mant2 = 8'd31; b_mant3 = 8'd32;
a_exp0 = 10'd981; a_exp1 = 10'd139; a_exp2 = 10'd639; a_exp3 = 10'd791;
b_exp0 = 10'd362; b_exp1 = 10'd735; b_exp2 = 10'd302; b_exp3 = 10'd504;
a_sign0 = 4'd4; a_sign1 = 4'd1; a_sign2 = 4'd14; a_sign3 = 4'd14;
b_sign0 = 4'd2; b_sign1 = 4'd2; b_sign2 = 4'd14; b_sign3 = 4'd7;
@(posedge clk_i);
a_mant0 = 8'd145; a_mant1 = 8'd14; a_mant2 = 8'd99; a_mant3 = 8'd21;
b_mant0 = 8'd147; b_mant1 = 8'd163; b_mant2 = 8'd81; b_mant3 = 8'd193;
a_exp0 = 10'd694; a_exp1 = 10'd123; a_exp2 = 10'd851; a_exp3 = 10'd744;
b_exp0 = 10'd732; b_exp1 = 10'd729; b_exp2 = 10'd64; b_exp3 = 10'd623;
a_sign0 = 4'd13; a_sign1 = 4'd7; a_sign2 = 4'd4; a_sign3 = 4'd8;
b_sign0 = 4'd9; b_sign1 = 4'd6; b_sign2 = 4'd8; b_sign3 = 4'd8;
@(posedge clk_i);
shared_exps0 = 8'd96;
shared_exps1 = 8'd119;
a_mant0 = 8'd139; a_mant1 = 8'd103; a_mant2 = 8'd164; a_mant3 = 8'd169;
b_mant0 = 8'd145; b_mant1 = 8'd38; b_mant2 = 8'd91; b_mant3 = 8'd56;
a_exp0 = 10'd230; a_exp1 = 10'd451; a_exp2 = 10'd472; a_exp3 = 10'd464;
b_exp0 = 10'd492; b_exp1 = 10'd430; b_exp2 = 10'd736; b_exp3 = 10'd260;
a_sign0 = 4'd12; a_sign1 = 4'd16; a_sign2 = 4'd5; a_sign3 = 4'd0;
b_sign0 = 4'd0; b_sign1 = 4'd1; b_sign2 = 4'd16; b_sign3 = 4'd14;
@(posedge clk_i);
a_mant0 = 8'd134; a_mant1 = 8'd188; a_mant2 = 8'd236; a_mant3 = 8'd84;
b_mant0 = 8'd156; b_mant1 = 8'd219; b_mant2 = 8'd20; b_mant3 = 8'd245;
a_exp0 = 10'd759; a_exp1 = 10'd912; a_exp2 = 10'd642; a_exp3 = 10'd210;
b_exp0 = 10'd45; b_exp1 = 10'd122; b_exp2 = 10'd702; b_exp3 = 10'd300;
a_sign0 = 4'd7; a_sign1 = 4'd10; a_sign2 = 4'd13; a_sign3 = 4'd9;
b_sign0 = 4'd13; b_sign1 = 4'd1; b_sign2 = 4'd5; b_sign3 = 4'd6;
@(posedge clk_i);
a_mant0 = 8'd161; a_mant1 = 8'd131; a_mant2 = 8'd232; a_mant3 = 8'd129;
b_mant0 = 8'd236; b_mant1 = 8'd26; b_mant2 = 8'd234; b_mant3 = 8'd219;
a_exp0 = 10'd102; a_exp1 = 10'd120; a_exp2 = 10'd896; a_exp3 = 10'd61;
b_exp0 = 10'd397; b_exp1 = 10'd621; b_exp2 = 10'd54; b_exp3 = 10'd859;
a_sign0 = 4'd13; a_sign1 = 4'd7; a_sign2 = 4'd3; a_sign3 = 4'd7;
b_sign0 = 4'd1; b_sign1 = 4'd5; b_sign2 = 4'd16; b_sign3 = 4'd4;
@(posedge clk_i);
a_mant0 = 8'd0; a_mant1 = 8'd246; a_mant2 = 8'd199; a_mant3 = 8'd21;
b_mant0 = 8'd182; b_mant1 = 8'd35; b_mant2 = 8'd59; b_mant3 = 8'd238;
a_exp0 = 10'd352; a_exp1 = 10'd799; a_exp2 = 10'd459; a_exp3 = 10'd303;
b_exp0 = 10'd607; b_exp1 = 10'd600; b_exp2 = 10'd509; b_exp3 = 10'd16;
a_sign0 = 4'd10; a_sign1 = 4'd10; a_sign2 = 4'd9; a_sign3 = 4'd8;
b_sign0 = 4'd2; b_sign1 = 4'd8; b_sign2 = 4'd3; b_sign3 = 4'd1;
@(posedge clk_i);
a_mant0 = 8'd237; a_mant1 = 8'd252; a_mant2 = 8'd172; a_mant3 = 8'd221;
b_mant0 = 8'd146; b_mant1 = 8'd135; b_mant2 = 8'd20; b_mant3 = 8'd29;
a_exp0 = 10'd1015; a_exp1 = 10'd351; a_exp2 = 10'd683; a_exp3 = 10'd174;
b_exp0 = 10'd917; b_exp1 = 10'd604; b_exp2 = 10'd394; b_exp3 = 10'd182;
a_sign0 = 4'd15; a_sign1 = 4'd11; a_sign2 = 4'd1; a_sign3 = 4'd14;
b_sign0 = 4'd12; b_sign1 = 4'd13; b_sign2 = 4'd15; b_sign3 = 4'd10;
@(posedge clk_i);
a_mant0 = 8'd175; a_mant1 = 8'd109; a_mant2 = 8'd247; a_mant3 = 8'd119;
b_mant0 = 8'd202; b_mant1 = 8'd68; b_mant2 = 8'd142; b_mant3 = 8'd210;
a_exp0 = 10'd465; a_exp1 = 10'd347; a_exp2 = 10'd74; a_exp3 = 10'd463;
b_exp0 = 10'd696; b_exp1 = 10'd328; b_exp2 = 10'd965; b_exp3 = 10'd807;
a_sign0 = 4'd0; a_sign1 = 4'd9; a_sign2 = 4'd4; a_sign3 = 4'd3;
b_sign0 = 4'd5; b_sign1 = 4'd2; b_sign2 = 4'd8; b_sign3 = 4'd3;
@(posedge clk_i);
a_mant0 = 8'd158; a_mant1 = 8'd221; a_mant2 = 8'd44; a_mant3 = 8'd57;
b_mant0 = 8'd101; b_mant1 = 8'd33; b_mant2 = 8'd147; b_mant3 = 8'd197;
a_exp0 = 10'd719; a_exp1 = 10'd794; a_exp2 = 10'd368; a_exp3 = 10'd884;
b_exp0 = 10'd225; b_exp1 = 10'd372; b_exp2 = 10'd913; b_exp3 = 10'd360;
a_sign0 = 4'd11; a_sign1 = 4'd0; a_sign2 = 4'd7; a_sign3 = 4'd10;
b_sign0 = 4'd8; b_sign1 = 4'd10; b_sign2 = 4'd1; b_sign3 = 4'd1;
@(posedge clk_i);
a_mant0 = 8'd39; a_mant1 = 8'd123; a_mant2 = 8'd191; a_mant3 = 8'd123;
b_mant0 = 8'd45; b_mant1 = 8'd74; b_mant2 = 8'd181; b_mant3 = 8'd127;
a_exp0 = 10'd24; a_exp1 = 10'd959; a_exp2 = 10'd211; a_exp3 = 10'd148;
b_exp0 = 10'd915; b_exp1 = 10'd867; b_exp2 = 10'd622; b_exp3 = 10'd492;
a_sign0 = 4'd8; a_sign1 = 4'd4; a_sign2 = 4'd3; a_sign3 = 4'd6;
b_sign0 = 4'd5; b_sign1 = 4'd16; b_sign2 = 4'd16; b_sign3 = 4'd2;
@(posedge clk_i);
shared_exps0 = 8'd137;
shared_exps1 = 8'd128;
a_mant0 = 8'd199; a_mant1 = 8'd160; a_mant2 = 8'd205; a_mant3 = 8'd84;
b_mant0 = 8'd115; b_mant1 = 8'd241; b_mant2 = 8'd67; b_mant3 = 8'd33;
a_exp0 = 10'd216; a_exp1 = 10'd983; a_exp2 = 10'd473; a_exp3 = 10'd207;
b_exp0 = 10'd877; b_exp1 = 10'd624; b_exp2 = 10'd948; b_exp3 = 10'd850;
a_sign0 = 4'd4; a_sign1 = 4'd10; a_sign2 = 4'd0; a_sign3 = 4'd10;
b_sign0 = 4'd8; b_sign1 = 4'd9; b_sign2 = 4'd2; b_sign3 = 4'd6;
@(posedge clk_i);
a_mant0 = 8'd164; a_mant1 = 8'd58; a_mant2 = 8'd34; a_mant3 = 8'd63;
b_mant0 = 8'd216; b_mant1 = 8'd83; b_mant2 = 8'd2; b_mant3 = 8'd2;
a_exp0 = 10'd932; a_exp1 = 10'd922; a_exp2 = 10'd194; a_exp3 = 10'd409;
b_exp0 = 10'd818; b_exp1 = 10'd70; b_exp2 = 10'd498; b_exp3 = 10'd1015;
a_sign0 = 4'd10; a_sign1 = 4'd5; a_sign2 = 4'd7; a_sign3 = 4'd6;
b_sign0 = 4'd10; b_sign1 = 4'd11; b_sign2 = 4'd14; b_sign3 = 4'd1;
@(posedge clk_i);
a_mant0 = 8'd192; a_mant1 = 8'd121; a_mant2 = 8'd197; a_mant3 = 8'd198;
b_mant0 = 8'd211; b_mant1 = 8'd115; b_mant2 = 8'd33; b_mant3 = 8'd28;
a_exp0 = 10'd496; a_exp1 = 10'd677; a_exp2 = 10'd130; a_exp3 = 10'd856;
b_exp0 = 10'd370; b_exp1 = 10'd672; b_exp2 = 10'd357; b_exp3 = 10'd186;
a_sign0 = 4'd8; a_sign1 = 4'd2; a_sign2 = 4'd15; a_sign3 = 4'd0;
b_sign0 = 4'd1; b_sign1 = 4'd10; b_sign2 = 4'd1; b_sign3 = 4'd4;
@(posedge clk_i);
a_mant0 = 8'd63; a_mant1 = 8'd94; a_mant2 = 8'd147; a_mant3 = 8'd79;
b_mant0 = 8'd19; b_mant1 = 8'd10; b_mant2 = 8'd153; b_mant3 = 8'd207;
a_exp0 = 10'd442; a_exp1 = 10'd114; a_exp2 = 10'd451; a_exp3 = 10'd755;
b_exp0 = 10'd737; b_exp1 = 10'd944; b_exp2 = 10'd277; b_exp3 = 10'd869;
a_sign0 = 4'd1; a_sign1 = 4'd3; a_sign2 = 4'd2; a_sign3 = 4'd6;
b_sign0 = 4'd14; b_sign1 = 4'd5; b_sign2 = 4'd1; b_sign3 = 4'd10;
@(posedge clk_i);
a_mant0 = 8'd97; a_mant1 = 8'd82; a_mant2 = 8'd13; a_mant3 = 8'd87;
b_mant0 = 8'd0; b_mant1 = 8'd240; b_mant2 = 8'd109; b_mant3 = 8'd43;
a_exp0 = 10'd911; a_exp1 = 10'd478; a_exp2 = 10'd516; a_exp3 = 10'd224;
b_exp0 = 10'd461; b_exp1 = 10'd940; b_exp2 = 10'd107; b_exp3 = 10'd326;
a_sign0 = 4'd16; a_sign1 = 4'd5; a_sign2 = 4'd4; a_sign3 = 4'd4;
b_sign0 = 4'd8; b_sign1 = 4'd13; b_sign2 = 4'd8; b_sign3 = 4'd2;
@(posedge clk_i);
a_mant0 = 8'd116; a_mant1 = 8'd157; a_mant2 = 8'd209; a_mant3 = 8'd211;
b_mant0 = 8'd63; b_mant1 = 8'd122; b_mant2 = 8'd47; b_mant3 = 8'd28;
a_exp0 = 10'd324; a_exp1 = 10'd988; a_exp2 = 10'd5; a_exp3 = 10'd472;
b_exp0 = 10'd324; b_exp1 = 10'd447; b_exp2 = 10'd578; b_exp3 = 10'd966;
a_sign0 = 4'd16; a_sign1 = 4'd16; a_sign2 = 4'd15; a_sign3 = 4'd7;
b_sign0 = 4'd2; b_sign1 = 4'd15; b_sign2 = 4'd0; b_sign3 = 4'd15;
@(posedge clk_i);
a_mant0 = 8'd179; a_mant1 = 8'd225; a_mant2 = 8'd64; a_mant3 = 8'd137;
b_mant0 = 8'd13; b_mant1 = 8'd116; b_mant2 = 8'd175; b_mant3 = 8'd243;
a_exp0 = 10'd405; a_exp1 = 10'd526; a_exp2 = 10'd93; a_exp3 = 10'd679;
b_exp0 = 10'd341; b_exp1 = 10'd936; b_exp2 = 10'd201; b_exp3 = 10'd422;
a_sign0 = 4'd8; a_sign1 = 4'd0; a_sign2 = 4'd4; a_sign3 = 4'd9;
b_sign0 = 4'd6; b_sign1 = 4'd1; b_sign2 = 4'd10; b_sign3 = 4'd16;
@(posedge clk_i);
a_mant0 = 8'd108; a_mant1 = 8'd122; a_mant2 = 8'd188; a_mant3 = 8'd179;
b_mant0 = 8'd99; b_mant1 = 8'd235; b_mant2 = 8'd210; b_mant3 = 8'd172;
a_exp0 = 10'd768; a_exp1 = 10'd845; a_exp2 = 10'd53; a_exp3 = 10'd349;
b_exp0 = 10'd802; b_exp1 = 10'd483; b_exp2 = 10'd960; b_exp3 = 10'd368;
a_sign0 = 4'd2; a_sign1 = 4'd8; a_sign2 = 4'd13; a_sign3 = 4'd6;
b_sign0 = 4'd15; b_sign1 = 4'd3; b_sign2 = 4'd1; b_sign3 = 4'd6;
@(posedge clk_i);
shared_exps0 = 8'd124;
shared_exps1 = 8'd124;
a_mant0 = 8'd66; a_mant1 = 8'd88; a_mant2 = 8'd55; a_mant3 = 8'd7;
b_mant0 = 8'd48; b_mant1 = 8'd93; b_mant2 = 8'd161; b_mant3 = 8'd84;
a_exp0 = 10'd536; a_exp1 = 10'd678; a_exp2 = 10'd242; a_exp3 = 10'd861;
b_exp0 = 10'd6; b_exp1 = 10'd447; b_exp2 = 10'd498; b_exp3 = 10'd740;
a_sign0 = 4'd12; a_sign1 = 4'd6; a_sign2 = 4'd7; a_sign3 = 4'd10;
b_sign0 = 4'd3; b_sign1 = 4'd2; b_sign2 = 4'd4; b_sign3 = 4'd0;
@(posedge clk_i);
a_mant0 = 8'd131; a_mant1 = 8'd205; a_mant2 = 8'd167; a_mant3 = 8'd147;
b_mant0 = 8'd160; b_mant1 = 8'd194; b_mant2 = 8'd13; b_mant3 = 8'd40;
a_exp0 = 10'd83; a_exp1 = 10'd315; a_exp2 = 10'd807; a_exp3 = 10'd414;
b_exp0 = 10'd573; b_exp1 = 10'd625; b_exp2 = 10'd13; b_exp3 = 10'd738;
a_sign0 = 4'd5; a_sign1 = 4'd16; a_sign2 = 4'd6; a_sign3 = 4'd8;
b_sign0 = 4'd1; b_sign1 = 4'd12; b_sign2 = 4'd10; b_sign3 = 4'd6;
@(posedge clk_i);
a_mant0 = 8'd214; a_mant1 = 8'd194; a_mant2 = 8'd63; a_mant3 = 8'd111;
b_mant0 = 8'd224; b_mant1 = 8'd117; b_mant2 = 8'd201; b_mant3 = 8'd243;
a_exp0 = 10'd340; a_exp1 = 10'd934; a_exp2 = 10'd155; a_exp3 = 10'd395;
b_exp0 = 10'd404; b_exp1 = 10'd193; b_exp2 = 10'd210; b_exp3 = 10'd368;
a_sign0 = 4'd11; a_sign1 = 4'd0; a_sign2 = 4'd6; a_sign3 = 4'd9;
b_sign0 = 4'd6; b_sign1 = 4'd14; b_sign2 = 4'd12; b_sign3 = 4'd0;
@(posedge clk_i);
a_mant0 = 8'd6; a_mant1 = 8'd60; a_mant2 = 8'd202; a_mant3 = 8'd20;
b_mant0 = 8'd125; b_mant1 = 8'd177; b_mant2 = 8'd238; b_mant3 = 8'd229;
a_exp0 = 10'd83; a_exp1 = 10'd1007; a_exp2 = 10'd885; a_exp3 = 10'd387;
b_exp0 = 10'd350; b_exp1 = 10'd843; b_exp2 = 10'd43; b_exp3 = 10'd884;
a_sign0 = 4'd11; a_sign1 = 4'd0; a_sign2 = 4'd7; a_sign3 = 4'd0;
b_sign0 = 4'd10; b_sign1 = 4'd11; b_sign2 = 4'd5; b_sign3 = 4'd14;
@(posedge clk_i);
a_mant0 = 8'd203; a_mant1 = 8'd119; a_mant2 = 8'd252; a_mant3 = 8'd111;
b_mant0 = 8'd240; b_mant1 = 8'd153; b_mant2 = 8'd141; b_mant3 = 8'd230;
a_exp0 = 10'd947; a_exp1 = 10'd63; a_exp2 = 10'd906; a_exp3 = 10'd450;
b_exp0 = 10'd974; b_exp1 = 10'd749; b_exp2 = 10'd170; b_exp3 = 10'd715;
a_sign0 = 4'd12; a_sign1 = 4'd11; a_sign2 = 4'd15; a_sign3 = 4'd16;
b_sign0 = 4'd6; b_sign1 = 4'd0; b_sign2 = 4'd7; b_sign3 = 4'd8;
@(posedge clk_i);
a_mant0 = 8'd134; a_mant1 = 8'd55; a_mant2 = 8'd78; a_mant3 = 8'd84;
b_mant0 = 8'd143; b_mant1 = 8'd43; b_mant2 = 8'd173; b_mant3 = 8'd158;
a_exp0 = 10'd7; a_exp1 = 10'd991; a_exp2 = 10'd934; a_exp3 = 10'd869;
b_exp0 = 10'd342; b_exp1 = 10'd159; b_exp2 = 10'd85; b_exp3 = 10'd922;
a_sign0 = 4'd9; a_sign1 = 4'd2; a_sign2 = 4'd10; a_sign3 = 4'd5;
b_sign0 = 4'd13; b_sign1 = 4'd1; b_sign2 = 4'd14; b_sign3 = 4'd12;
@(posedge clk_i);
a_mant0 = 8'd60; a_mant1 = 8'd60; a_mant2 = 8'd126; a_mant3 = 8'd131;
b_mant0 = 8'd27; b_mant1 = 8'd167; b_mant2 = 8'd169; b_mant3 = 8'd93;
a_exp0 = 10'd834; a_exp1 = 10'd2; a_exp2 = 10'd404; a_exp3 = 10'd554;
b_exp0 = 10'd546; b_exp1 = 10'd1010; b_exp2 = 10'd882; b_exp3 = 10'd744;
a_sign0 = 4'd16; a_sign1 = 4'd4; a_sign2 = 4'd6; a_sign3 = 4'd0;
b_sign0 = 4'd14; b_sign1 = 4'd12; b_sign2 = 4'd0; b_sign3 = 4'd12;
@(posedge clk_i);
a_mant0 = 8'd27; a_mant1 = 8'd8; a_mant2 = 8'd149; a_mant3 = 8'd226;
b_mant0 = 8'd255; b_mant1 = 8'd209; b_mant2 = 8'd118; b_mant3 = 8'd62;
a_exp0 = 10'd235; a_exp1 = 10'd129; a_exp2 = 10'd873; a_exp3 = 10'd492;
b_exp0 = 10'd389; b_exp1 = 10'd350; b_exp2 = 10'd381; b_exp3 = 10'd56;
a_sign0 = 4'd0; a_sign1 = 4'd13; a_sign2 = 4'd2; a_sign3 = 4'd15;
b_sign0 = 4'd10; b_sign1 = 4'd13; b_sign2 = 4'd11; b_sign3 = 4'd8;
@(posedge clk_i);
shared_exps0 = 8'd142;
shared_exps1 = 8'd121;
rstn = 0;
@(posedge clk_i);
rstn = 1;
a_mant0 = 8'd122; a_mant1 = 8'd136; a_mant2 = 8'd18; a_mant3 = 8'd140;
b_mant0 = 8'd203; b_mant1 = 8'd71; b_mant2 = 8'd123; b_mant3 = 8'd158;
a_exp0 = 10'd589; a_exp1 = 10'd885; a_exp2 = 10'd493; a_exp3 = 10'd339;
b_exp0 = 10'd623; b_exp1 = 10'd338; b_exp2 = 10'd317; b_exp3 = 10'd795;
a_sign0 = 4'd0; a_sign1 = 4'd0; a_sign2 = 4'd10; a_sign3 = 4'd1;
b_sign0 = 4'd13; b_sign1 = 4'd16; b_sign2 = 4'd15; b_sign3 = 4'd15;
@(posedge clk_i);
a_mant0 = 8'd53; a_mant1 = 8'd161; a_mant2 = 8'd84; a_mant3 = 8'd203;
b_mant0 = 8'd110; b_mant1 = 8'd40; b_mant2 = 8'd170; b_mant3 = 8'd85;
a_exp0 = 10'd332; a_exp1 = 10'd923; a_exp2 = 10'd127; a_exp3 = 10'd783;
b_exp0 = 10'd982; b_exp1 = 10'd587; b_exp2 = 10'd162; b_exp3 = 10'd258;
a_sign0 = 4'd10; a_sign1 = 4'd11; a_sign2 = 4'd3; a_sign3 = 4'd13;
b_sign0 = 4'd8; b_sign1 = 4'd13; b_sign2 = 4'd11; b_sign3 = 4'd5;
@(posedge clk_i);
a_mant0 = 8'd34; a_mant1 = 8'd239; a_mant2 = 8'd186; a_mant3 = 8'd247;
b_mant0 = 8'd39; b_mant1 = 8'd66; b_mant2 = 8'd213; b_mant3 = 8'd225;
a_exp0 = 10'd456; a_exp1 = 10'd18; a_exp2 = 10'd462; a_exp3 = 10'd628;
b_exp0 = 10'd310; b_exp1 = 10'd229; b_exp2 = 10'd333; b_exp3 = 10'd846;
a_sign0 = 4'd2; a_sign1 = 4'd4; a_sign2 = 4'd15; a_sign3 = 4'd7;
b_sign0 = 4'd10; b_sign1 = 4'd16; b_sign2 = 4'd6; b_sign3 = 4'd11;
@(posedge clk_i);
a_mant0 = 8'd38; a_mant1 = 8'd82; a_mant2 = 8'd105; a_mant3 = 8'd27;
b_mant0 = 8'd131; b_mant1 = 8'd239; b_mant2 = 8'd176; b_mant3 = 8'd70;
a_exp0 = 10'd482; a_exp1 = 10'd758; a_exp2 = 10'd1009; a_exp3 = 10'd772;
b_exp0 = 10'd804; b_exp1 = 10'd641; b_exp2 = 10'd340; b_exp3 = 10'd467;
a_sign0 = 4'd13; a_sign1 = 4'd4; a_sign2 = 4'd1; a_sign3 = 4'd6;
b_sign0 = 4'd2; b_sign1 = 4'd3; b_sign2 = 4'd12; b_sign3 = 4'd4;
@(posedge clk_i);
a_mant0 = 8'd240; a_mant1 = 8'd116; a_mant2 = 8'd10; a_mant3 = 8'd189;
b_mant0 = 8'd46; b_mant1 = 8'd102; b_mant2 = 8'd79; b_mant3 = 8'd6;
a_exp0 = 10'd100; a_exp1 = 10'd509; a_exp2 = 10'd743; a_exp3 = 10'd798;
b_exp0 = 10'd660; b_exp1 = 10'd323; b_exp2 = 10'd446; b_exp3 = 10'd223;
a_sign0 = 4'd14; a_sign1 = 4'd6; a_sign2 = 4'd8; a_sign3 = 4'd16;
b_sign0 = 4'd11; b_sign1 = 4'd4; b_sign2 = 4'd5; b_sign3 = 4'd12;
@(posedge clk_i);
a_mant0 = 8'd90; a_mant1 = 8'd210; a_mant2 = 8'd31; a_mant3 = 8'd85;
b_mant0 = 8'd98; b_mant1 = 8'd20; b_mant2 = 8'd201; b_mant3 = 8'd32;
a_exp0 = 10'd308; a_exp1 = 10'd463; a_exp2 = 10'd913; a_exp3 = 10'd320;
b_exp0 = 10'd752; b_exp1 = 10'd657; b_exp2 = 10'd761; b_exp3 = 10'd901;
a_sign0 = 4'd15; a_sign1 = 4'd9; a_sign2 = 4'd6; a_sign3 = 4'd2;
b_sign0 = 4'd11; b_sign1 = 4'd3; b_sign2 = 4'd9; b_sign3 = 4'd13;
@(posedge clk_i);
a_mant0 = 8'd6; a_mant1 = 8'd18; a_mant2 = 8'd157; a_mant3 = 8'd211;
b_mant0 = 8'd181; b_mant1 = 8'd120; b_mant2 = 8'd16; b_mant3 = 8'd114;
a_exp0 = 10'd939; a_exp1 = 10'd89; a_exp2 = 10'd958; a_exp3 = 10'd454;
b_exp0 = 10'd919; b_exp1 = 10'd927; b_exp2 = 10'd952; b_exp3 = 10'd567;
a_sign0 = 4'd12; a_sign1 = 4'd14; a_sign2 = 4'd2; a_sign3 = 4'd13;
b_sign0 = 4'd10; b_sign1 = 4'd0; b_sign2 = 4'd2; b_sign3 = 4'd0;
@(posedge clk_i);
shared_exps0 = 8'd141;
shared_exps1 = 8'd116;
a_mant0 = 8'd114; a_mant1 = 8'd217; a_mant2 = 8'd170; a_mant3 = 8'd107;
b_mant0 = 8'd71; b_mant1 = 8'd18; b_mant2 = 8'd86; b_mant3 = 8'd208;
a_exp0 = 10'd213; a_exp1 = 10'd851; a_exp2 = 10'd239; a_exp3 = 10'd314;
b_exp0 = 10'd55; b_exp1 = 10'd594; b_exp2 = 10'd543; b_exp3 = 10'd460;
a_sign0 = 4'd11; a_sign1 = 4'd11; a_sign2 = 4'd1; a_sign3 = 4'd0;
b_sign0 = 4'd0; b_sign1 = 4'd6; b_sign2 = 4'd13; b_sign3 = 4'd1;
@(posedge clk_i);
a_mant0 = 8'd80; a_mant1 = 8'd199; a_mant2 = 8'd120; a_mant3 = 8'd98;
b_mant0 = 8'd240; b_mant1 = 8'd232; b_mant2 = 8'd46; b_mant3 = 8'd216;
a_exp0 = 10'd237; a_exp1 = 10'd954; a_exp2 = 10'd727; a_exp3 = 10'd932;
b_exp0 = 10'd305; b_exp1 = 10'd75; b_exp2 = 10'd709; b_exp3 = 10'd592;
a_sign0 = 4'd8; a_sign1 = 4'd11; a_sign2 = 4'd15; a_sign3 = 4'd7;
b_sign0 = 4'd8; b_sign1 = 4'd3; b_sign2 = 4'd0; b_sign3 = 4'd6;
@(posedge clk_i);
a_mant0 = 8'd29; a_mant1 = 8'd247; a_mant2 = 8'd169; a_mant3 = 8'd60;
b_mant0 = 8'd155; b_mant1 = 8'd118; b_mant2 = 8'd238; b_mant3 = 8'd179;
a_exp0 = 10'd943; a_exp1 = 10'd298; a_exp2 = 10'd927; a_exp3 = 10'd907;
b_exp0 = 10'd489; b_exp1 = 10'd193; b_exp2 = 10'd524; b_exp3 = 10'd928;
a_sign0 = 4'd0; a_sign1 = 4'd6; a_sign2 = 4'd9; a_sign3 = 4'd7;
b_sign0 = 4'd4; b_sign1 = 4'd3; b_sign2 = 4'd10; b_sign3 = 4'd8;
@(posedge clk_i);
a_mant0 = 8'd182; a_mant1 = 8'd86; a_mant2 = 8'd39; a_mant3 = 8'd1;
b_mant0 = 8'd82; b_mant1 = 8'd152; b_mant2 = 8'd68; b_mant3 = 8'd93;
a_exp0 = 10'd508; a_exp1 = 10'd119; a_exp2 = 10'd485; a_exp3 = 10'd245;
b_exp0 = 10'd271; b_exp1 = 10'd746; b_exp2 = 10'd425; b_exp3 = 10'd20;
a_sign0 = 4'd7; a_sign1 = 4'd16; a_sign2 = 4'd9; a_sign3 = 4'd4;
b_sign0 = 4'd13; b_sign1 = 4'd14; b_sign2 = 4'd10; b_sign3 = 4'd0;
@(posedge clk_i);
a_mant0 = 8'd31; a_mant1 = 8'd104; a_mant2 = 8'd144; a_mant3 = 8'd179;
b_mant0 = 8'd157; b_mant1 = 8'd170; b_mant2 = 8'd22; b_mant3 = 8'd9;
a_exp0 = 10'd784; a_exp1 = 10'd458; a_exp2 = 10'd49; a_exp3 = 10'd887;
b_exp0 = 10'd1011; b_exp1 = 10'd369; b_exp2 = 10'd349; b_exp3 = 10'd946;
a_sign0 = 4'd16; a_sign1 = 4'd0; a_sign2 = 4'd1; a_sign3 = 4'd9;
b_sign0 = 4'd4; b_sign1 = 4'd4; b_sign2 = 4'd6; b_sign3 = 4'd16;
@(posedge clk_i);
a_mant0 = 8'd45; a_mant1 = 8'd250; a_mant2 = 8'd142; a_mant3 = 8'd154;
b_mant0 = 8'd184; b_mant1 = 8'd156; b_mant2 = 8'd92; b_mant3 = 8'd7;
a_exp0 = 10'd604; a_exp1 = 10'd696; a_exp2 = 10'd611; a_exp3 = 10'd519;
b_exp0 = 10'd699; b_exp1 = 10'd487; b_exp2 = 10'd763; b_exp3 = 10'd517;
a_sign0 = 4'd1; a_sign1 = 4'd9; a_sign2 = 4'd0; a_sign3 = 4'd7;
b_sign0 = 4'd6; b_sign1 = 4'd1; b_sign2 = 4'd10; b_sign3 = 4'd2;
@(posedge clk_i);
a_mant0 = 8'd167; a_mant1 = 8'd187; a_mant2 = 8'd118; a_mant3 = 8'd175;
b_mant0 = 8'd121; b_mant1 = 8'd120; b_mant2 = 8'd52; b_mant3 = 8'd240;
a_exp0 = 10'd851; a_exp1 = 10'd675; a_exp2 = 10'd822; a_exp3 = 10'd585;
b_exp0 = 10'd141; b_exp1 = 10'd998; b_exp2 = 10'd537; b_exp3 = 10'd563;
a_sign0 = 4'd10; a_sign1 = 4'd13; a_sign2 = 4'd0; a_sign3 = 4'd11;
b_sign0 = 4'd5; b_sign1 = 4'd14; b_sign2 = 4'd14; b_sign3 = 4'd3;
@(posedge clk_i);
a_mant0 = 8'd14; a_mant1 = 8'd252; a_mant2 = 8'd58; a_mant3 = 8'd91;
b_mant0 = 8'd99; b_mant1 = 8'd104; b_mant2 = 8'd13; b_mant3 = 8'd192;
a_exp0 = 10'd34; a_exp1 = 10'd425; a_exp2 = 10'd400; a_exp3 = 10'd205;
b_exp0 = 10'd298; b_exp1 = 10'd267; b_exp2 = 10'd242; b_exp3 = 10'd1008;
a_sign0 = 4'd7; a_sign1 = 4'd13; a_sign2 = 4'd7; a_sign3 = 4'd0;
b_sign0 = 4'd5; b_sign1 = 4'd14; b_sign2 = 4'd1; b_sign3 = 4'd0;
@(posedge clk_i);
shared_exps0 = 8'd149;
shared_exps1 = 8'd138;
a_mant0 = 8'd245; a_mant1 = 8'd111; a_mant2 = 8'd129; a_mant3 = 8'd212;
b_mant0 = 8'd169; b_mant1 = 8'd196; b_mant2 = 8'd28; b_mant3 = 8'd106;
a_exp0 = 10'd276; a_exp1 = 10'd192; a_exp2 = 10'd234; a_exp3 = 10'd804;
b_exp0 = 10'd428; b_exp1 = 10'd527; b_exp2 = 10'd424; b_exp3 = 10'd994;
a_sign0 = 4'd2; a_sign1 = 4'd6; a_sign2 = 4'd7; a_sign3 = 4'd6;
b_sign0 = 4'd6; b_sign1 = 4'd1; b_sign2 = 4'd13; b_sign3 = 4'd16;
@(posedge clk_i);
a_mant0 = 8'd69; a_mant1 = 8'd240; a_mant2 = 8'd139; a_mant3 = 8'd227;
b_mant0 = 8'd175; b_mant1 = 8'd30; b_mant2 = 8'd49; b_mant3 = 8'd90;
a_exp0 = 10'd684; a_exp1 = 10'd514; a_exp2 = 10'd776; a_exp3 = 10'd603;
b_exp0 = 10'd505; b_exp1 = 10'd186; b_exp2 = 10'd35; b_exp3 = 10'd676;
a_sign0 = 4'd13; a_sign1 = 4'd8; a_sign2 = 4'd10; a_sign3 = 4'd0;
b_sign0 = 4'd10; b_sign1 = 4'd12; b_sign2 = 4'd0; b_sign3 = 4'd13;
@(posedge clk_i);
a_mant0 = 8'd104; a_mant1 = 8'd41; a_mant2 = 8'd178; a_mant3 = 8'd184;
b_mant0 = 8'd227; b_mant1 = 8'd79; b_mant2 = 8'd21; b_mant3 = 8'd25;
a_exp0 = 10'd227; a_exp1 = 10'd1004; a_exp2 = 10'd1008; a_exp3 = 10'd182;
b_exp0 = 10'd660; b_exp1 = 10'd562; b_exp2 = 10'd311; b_exp3 = 10'd390;
a_sign0 = 4'd1; a_sign1 = 4'd5; a_sign2 = 4'd0; a_sign3 = 4'd0;
b_sign0 = 4'd13; b_sign1 = 4'd6; b_sign2 = 4'd6; b_sign3 = 4'd7;
@(posedge clk_i);
a_mant0 = 8'd249; a_mant1 = 8'd246; a_mant2 = 8'd148; a_mant3 = 8'd242;
b_mant0 = 8'd173; b_mant1 = 8'd73; b_mant2 = 8'd93; b_mant3 = 8'd33;
a_exp0 = 10'd101; a_exp1 = 10'd601; a_exp2 = 10'd293; a_exp3 = 10'd823;
b_exp0 = 10'd320; b_exp1 = 10'd587; b_exp2 = 10'd569; b_exp3 = 10'd928;
a_sign0 = 4'd8; a_sign1 = 4'd11; a_sign2 = 4'd0; a_sign3 = 4'd13;
b_sign0 = 4'd3; b_sign1 = 4'd16; b_sign2 = 4'd14; b_sign3 = 4'd6;
@(posedge clk_i);
a_mant0 = 8'd71; a_mant1 = 8'd141; a_mant2 = 8'd92; a_mant3 = 8'd25;
b_mant0 = 8'd139; b_mant1 = 8'd206; b_mant2 = 8'd149; b_mant3 = 8'd21;
a_exp0 = 10'd398; a_exp1 = 10'd63; a_exp2 = 10'd777; a_exp3 = 10'd345;
b_exp0 = 10'd893; b_exp1 = 10'd898; b_exp2 = 10'd716; b_exp3 = 10'd95;
a_sign0 = 4'd15; a_sign1 = 4'd3; a_sign2 = 4'd0; a_sign3 = 4'd12;
b_sign0 = 4'd16; b_sign1 = 4'd3; b_sign2 = 4'd0; b_sign3 = 4'd3;
@(posedge clk_i);
a_mant0 = 8'd14; a_mant1 = 8'd203; a_mant2 = 8'd218; a_mant3 = 8'd173;
b_mant0 = 8'd115; b_mant1 = 8'd39; b_mant2 = 8'd53; b_mant3 = 8'd34;
a_exp0 = 10'd873; a_exp1 = 10'd599; a_exp2 = 10'd712; a_exp3 = 10'd612;
b_exp0 = 10'd344; b_exp1 = 10'd593; b_exp2 = 10'd917; b_exp3 = 10'd174;
a_sign0 = 4'd10; a_sign1 = 4'd2; a_sign2 = 4'd11; a_sign3 = 4'd11;
b_sign0 = 4'd10; b_sign1 = 4'd15; b_sign2 = 4'd7; b_sign3 = 4'd13;
@(posedge clk_i);
a_mant0 = 8'd199; a_mant1 = 8'd174; a_mant2 = 8'd128; a_mant3 = 8'd197;
b_mant0 = 8'd3; b_mant1 = 8'd73; b_mant2 = 8'd133; b_mant3 = 8'd49;
a_exp0 = 10'd245; a_exp1 = 10'd10; a_exp2 = 10'd480; a_exp3 = 10'd908;
b_exp0 = 10'd638; b_exp1 = 10'd986; b_exp2 = 10'd427; b_exp3 = 10'd395;
a_sign0 = 4'd4; a_sign1 = 4'd7; a_sign2 = 4'd12; a_sign3 = 4'd10;
b_sign0 = 4'd15; b_sign1 = 4'd5; b_sign2 = 4'd8; b_sign3 = 4'd11;
@(posedge clk_i);
a_mant0 = 8'd196; a_mant1 = 8'd100; a_mant2 = 8'd212; a_mant3 = 8'd209;
b_mant0 = 8'd62; b_mant1 = 8'd53; b_mant2 = 8'd35; b_mant3 = 8'd229;
a_exp0 = 10'd443; a_exp1 = 10'd234; a_exp2 = 10'd936; a_exp3 = 10'd177;
b_exp0 = 10'd966; b_exp1 = 10'd0; b_exp2 = 10'd449; b_exp3 = 10'd593;
a_sign0 = 4'd15; a_sign1 = 4'd7; a_sign2 = 4'd2; a_sign3 = 4'd15;
b_sign0 = 4'd6; b_sign1 = 4'd6; b_sign2 = 4'd14; b_sign3 = 4'd6;
@(posedge clk_i);
shared_exps0 = 8'd118;
shared_exps1 = 8'd143;
a_mant0 = 8'd96; a_mant1 = 8'd137; a_mant2 = 8'd119; a_mant3 = 8'd112;
b_mant0 = 8'd99; b_mant1 = 8'd31; b_mant2 = 8'd177; b_mant3 = 8'd229;
a_exp0 = 10'd339; a_exp1 = 10'd540; a_exp2 = 10'd751; a_exp3 = 10'd532;
b_exp0 = 10'd543; b_exp1 = 10'd775; b_exp2 = 10'd192; b_exp3 = 10'd105;
a_sign0 = 4'd9; a_sign1 = 4'd12; a_sign2 = 4'd1; a_sign3 = 4'd9;
b_sign0 = 4'd12; b_sign1 = 4'd3; b_sign2 = 4'd13; b_sign3 = 4'd8;
@(posedge clk_i);
a_mant0 = 8'd66; a_mant1 = 8'd179; a_mant2 = 8'd109; a_mant3 = 8'd150;
b_mant0 = 8'd231; b_mant1 = 8'd99; b_mant2 = 8'd211; b_mant3 = 8'd54;
a_exp0 = 10'd545; a_exp1 = 10'd537; a_exp2 = 10'd869; a_exp3 = 10'd144;
b_exp0 = 10'd935; b_exp1 = 10'd241; b_exp2 = 10'd705; b_exp3 = 10'd667;
a_sign0 = 4'd1; a_sign1 = 4'd3; a_sign2 = 4'd13; a_sign3 = 4'd10;
b_sign0 = 4'd13; b_sign1 = 4'd12; b_sign2 = 4'd9; b_sign3 = 4'd13;
@(posedge clk_i);
a_mant0 = 8'd29; a_mant1 = 8'd67; a_mant2 = 8'd95; a_mant3 = 8'd154;
b_mant0 = 8'd116; b_mant1 = 8'd36; b_mant2 = 8'd251; b_mant3 = 8'd139;
a_exp0 = 10'd633; a_exp1 = 10'd561; a_exp2 = 10'd33; a_exp3 = 10'd575;
b_exp0 = 10'd537; b_exp1 = 10'd118; b_exp2 = 10'd852; b_exp3 = 10'd762;
a_sign0 = 4'd12; a_sign1 = 4'd15; a_sign2 = 4'd7; a_sign3 = 4'd6;
b_sign0 = 4'd11; b_sign1 = 4'd14; b_sign2 = 4'd15; b_sign3 = 4'd15;
@(posedge clk_i);
a_mant0 = 8'd231; a_mant1 = 8'd101; a_mant2 = 8'd111; a_mant3 = 8'd212;
b_mant0 = 8'd151; b_mant1 = 8'd176; b_mant2 = 8'd238; b_mant3 = 8'd231;
a_exp0 = 10'd767; a_exp1 = 10'd810; a_exp2 = 10'd982; a_exp3 = 10'd475;
b_exp0 = 10'd87; b_exp1 = 10'd42; b_exp2 = 10'd301; b_exp3 = 10'd226;
a_sign0 = 4'd4; a_sign1 = 4'd6; a_sign2 = 4'd15; a_sign3 = 4'd7;
b_sign0 = 4'd6; b_sign1 = 4'd12; b_sign2 = 4'd13; b_sign3 = 4'd4;
@(posedge clk_i);
a_mant0 = 8'd237; a_mant1 = 8'd34; a_mant2 = 8'd97; a_mant3 = 8'd189;
b_mant0 = 8'd243; b_mant1 = 8'd194; b_mant2 = 8'd81; b_mant3 = 8'd118;
a_exp0 = 10'd103; a_exp1 = 10'd413; a_exp2 = 10'd167; a_exp3 = 10'd563;
b_exp0 = 10'd864; b_exp1 = 10'd46; b_exp2 = 10'd562; b_exp3 = 10'd1009;
a_sign0 = 4'd5; a_sign1 = 4'd10; a_sign2 = 4'd6; a_sign3 = 4'd15;
b_sign0 = 4'd11; b_sign1 = 4'd9; b_sign2 = 4'd2; b_sign3 = 4'd4;
@(posedge clk_i);
a_mant0 = 8'd234; a_mant1 = 8'd93; a_mant2 = 8'd207; a_mant3 = 8'd234;
b_mant0 = 8'd80; b_mant1 = 8'd12; b_mant2 = 8'd72; b_mant3 = 8'd163;
a_exp0 = 10'd740; a_exp1 = 10'd102; a_exp2 = 10'd584; a_exp3 = 10'd212;
b_exp0 = 10'd1009; b_exp1 = 10'd982; b_exp2 = 10'd835; b_exp3 = 10'd640;
a_sign0 = 4'd8; a_sign1 = 4'd13; a_sign2 = 4'd8; a_sign3 = 4'd13;
b_sign0 = 4'd8; b_sign1 = 4'd10; b_sign2 = 4'd14; b_sign3 = 4'd1;
@(posedge clk_i);
a_mant0 = 8'd206; a_mant1 = 8'd215; a_mant2 = 8'd125; a_mant3 = 8'd116;
b_mant0 = 8'd117; b_mant1 = 8'd135; b_mant2 = 8'd47; b_mant3 = 8'd104;
a_exp0 = 10'd94; a_exp1 = 10'd758; a_exp2 = 10'd17; a_exp3 = 10'd728;
b_exp0 = 10'd985; b_exp1 = 10'd574; b_exp2 = 10'd430; b_exp3 = 10'd940;
a_sign0 = 4'd7; a_sign1 = 4'd4; a_sign2 = 4'd9; a_sign3 = 4'd6;
b_sign0 = 4'd2; b_sign1 = 4'd16; b_sign2 = 4'd6; b_sign3 = 4'd7;
@(posedge clk_i);
a_mant0 = 8'd157; a_mant1 = 8'd152; a_mant2 = 8'd245; a_mant3 = 8'd21;
b_mant0 = 8'd203; b_mant1 = 8'd183; b_mant2 = 8'd88; b_mant3 = 8'd239;
a_exp0 = 10'd868; a_exp1 = 10'd818; a_exp2 = 10'd900; a_exp3 = 10'd902;
b_exp0 = 10'd110; b_exp1 = 10'd198; b_exp2 = 10'd460; b_exp3 = 10'd203;
a_sign0 = 4'd1; a_sign1 = 4'd5; a_sign2 = 4'd12; a_sign3 = 4'd12;
b_sign0 = 4'd6; b_sign1 = 4'd16; b_sign2 = 4'd14; b_sign3 = 4'd5;
@(posedge clk_i);
shared_exps0 = 8'd121;
shared_exps1 = 8'd126;
rstn = 0;
@(posedge clk_i);
rstn = 1;
a_mant0 = 8'd138; a_mant1 = 8'd87; a_mant2 = 8'd210; a_mant3 = 8'd92;
b_mant0 = 8'd0; b_mant1 = 8'd73; b_mant2 = 8'd108; b_mant3 = 8'd102;
a_exp0 = 10'd327; a_exp1 = 10'd488; a_exp2 = 10'd478; a_exp3 = 10'd44;
b_exp0 = 10'd132; b_exp1 = 10'd112; b_exp2 = 10'd1006; b_exp3 = 10'd975;
a_sign0 = 4'd1; a_sign1 = 4'd0; a_sign2 = 4'd8; a_sign3 = 4'd11;
b_sign0 = 4'd8; b_sign1 = 4'd12; b_sign2 = 4'd0; b_sign3 = 4'd15;
@(posedge clk_i);
a_mant0 = 8'd126; a_mant1 = 8'd188; a_mant2 = 8'd104; a_mant3 = 8'd157;
b_mant0 = 8'd152; b_mant1 = 8'd182; b_mant2 = 8'd55; b_mant3 = 8'd156;
a_exp0 = 10'd339; a_exp1 = 10'd5; a_exp2 = 10'd484; a_exp3 = 10'd399;
b_exp0 = 10'd700; b_exp1 = 10'd786; b_exp2 = 10'd759; b_exp3 = 10'd909;
a_sign0 = 4'd6; a_sign1 = 4'd10; a_sign2 = 4'd12; a_sign3 = 4'd4;
b_sign0 = 4'd15; b_sign1 = 4'd12; b_sign2 = 4'd10; b_sign3 = 4'd16;
@(posedge clk_i);
a_mant0 = 8'd205; a_mant1 = 8'd32; a_mant2 = 8'd244; a_mant3 = 8'd51;
b_mant0 = 8'd55; b_mant1 = 8'd210; b_mant2 = 8'd83; b_mant3 = 8'd24;
a_exp0 = 10'd930; a_exp1 = 10'd98; a_exp2 = 10'd885; a_exp3 = 10'd595;
b_exp0 = 10'd474; b_exp1 = 10'd418; b_exp2 = 10'd422; b_exp3 = 10'd410;
a_sign0 = 4'd8; a_sign1 = 4'd1; a_sign2 = 4'd7; a_sign3 = 4'd11;
b_sign0 = 4'd8; b_sign1 = 4'd0; b_sign2 = 4'd11; b_sign3 = 4'd4;
@(posedge clk_i);
a_mant0 = 8'd214; a_mant1 = 8'd3; a_mant2 = 8'd98; a_mant3 = 8'd155;
b_mant0 = 8'd41; b_mant1 = 8'd224; b_mant2 = 8'd202; b_mant3 = 8'd105;
a_exp0 = 10'd852; a_exp1 = 10'd431; a_exp2 = 10'd355; a_exp3 = 10'd174;
b_exp0 = 10'd319; b_exp1 = 10'd1; b_exp2 = 10'd886; b_exp3 = 10'd614;
a_sign0 = 4'd8; a_sign1 = 4'd2; a_sign2 = 4'd2; a_sign3 = 4'd8;
b_sign0 = 4'd2; b_sign1 = 4'd9; b_sign2 = 4'd1; b_sign3 = 4'd5;
@(posedge clk_i);
a_mant0 = 8'd52; a_mant1 = 8'd194; a_mant2 = 8'd226; a_mant3 = 8'd80;
b_mant0 = 8'd136; b_mant1 = 8'd163; b_mant2 = 8'd84; b_mant3 = 8'd21;
a_exp0 = 10'd981; a_exp1 = 10'd655; a_exp2 = 10'd908; a_exp3 = 10'd829;
b_exp0 = 10'd86; b_exp1 = 10'd251; b_exp2 = 10'd993; b_exp3 = 10'd931;
a_sign0 = 4'd10; a_sign1 = 4'd15; a_sign2 = 4'd15; a_sign3 = 4'd7;
b_sign0 = 4'd10; b_sign1 = 4'd12; b_sign2 = 4'd2; b_sign3 = 4'd3;
@(posedge clk_i);
a_mant0 = 8'd139; a_mant1 = 8'd106; a_mant2 = 8'd164; a_mant3 = 8'd86;
b_mant0 = 8'd80; b_mant1 = 8'd53; b_mant2 = 8'd161; b_mant3 = 8'd124;
a_exp0 = 10'd946; a_exp1 = 10'd590; a_exp2 = 10'd165; a_exp3 = 10'd352;
b_exp0 = 10'd334; b_exp1 = 10'd807; b_exp2 = 10'd541; b_exp3 = 10'd915;
a_sign0 = 4'd2; a_sign1 = 4'd2; a_sign2 = 4'd13; a_sign3 = 4'd0;
b_sign0 = 4'd2; b_sign1 = 4'd0; b_sign2 = 4'd8; b_sign3 = 4'd3;
@(posedge clk_i);
a_mant0 = 8'd136; a_mant1 = 8'd114; a_mant2 = 8'd22; a_mant3 = 8'd234;
b_mant0 = 8'd227; b_mant1 = 8'd191; b_mant2 = 8'd25; b_mant3 = 8'd38;
a_exp0 = 10'd315; a_exp1 = 10'd969; a_exp2 = 10'd411; a_exp3 = 10'd72;
b_exp0 = 10'd887; b_exp1 = 10'd204; b_exp2 = 10'd99; b_exp3 = 10'd863;
a_sign0 = 4'd11; a_sign1 = 4'd5; a_sign2 = 4'd15; a_sign3 = 4'd8;
b_sign0 = 4'd1; b_sign1 = 4'd4; b_sign2 = 4'd13; b_sign3 = 4'd14;
@(posedge clk_i);
shared_exps0 = 8'd132;
shared_exps1 = 8'd122;
a_mant0 = 8'd160; a_mant1 = 8'd212; a_mant2 = 8'd131; a_mant3 = 8'd70;
b_mant0 = 8'd240; b_mant1 = 8'd255; b_mant2 = 8'd55; b_mant3 = 8'd139;
a_exp0 = 10'd60; a_exp1 = 10'd785; a_exp2 = 10'd179; a_exp3 = 10'd507;
b_exp0 = 10'd839; b_exp1 = 10'd293; b_exp2 = 10'd481; b_exp3 = 10'd216;
a_sign0 = 4'd2; a_sign1 = 4'd6; a_sign2 = 4'd8; a_sign3 = 4'd9;
b_sign0 = 4'd9; b_sign1 = 4'd2; b_sign2 = 4'd10; b_sign3 = 4'd3;
@(posedge clk_i);
a_mant0 = 8'd168; a_mant1 = 8'd37; a_mant2 = 8'd115; a_mant3 = 8'd99;
b_mant0 = 8'd141; b_mant1 = 8'd112; b_mant2 = 8'd137; b_mant3 = 8'd27;
a_exp0 = 10'd632; a_exp1 = 10'd408; a_exp2 = 10'd116; a_exp3 = 10'd982;
b_exp0 = 10'd840; b_exp1 = 10'd1018; b_exp2 = 10'd507; b_exp3 = 10'd605;
a_sign0 = 4'd9; a_sign1 = 4'd5; a_sign2 = 4'd2; a_sign3 = 4'd6;
b_sign0 = 4'd9; b_sign1 = 4'd12; b_sign2 = 4'd14; b_sign3 = 4'd12;
@(posedge clk_i);
a_mant0 = 8'd35; a_mant1 = 8'd229; a_mant2 = 8'd254; a_mant3 = 8'd126;
b_mant0 = 8'd46; b_mant1 = 8'd213; b_mant2 = 8'd145; b_mant3 = 8'd50;
a_exp0 = 10'd953; a_exp1 = 10'd764; a_exp2 = 10'd271; a_exp3 = 10'd42;
b_exp0 = 10'd121; b_exp1 = 10'd717; b_exp2 = 10'd578; b_exp3 = 10'd392;
a_sign0 = 4'd16; a_sign1 = 4'd11; a_sign2 = 4'd4; a_sign3 = 4'd3;
b_sign0 = 4'd16; b_sign1 = 4'd14; b_sign2 = 4'd6; b_sign3 = 4'd13;
@(posedge clk_i);
a_mant0 = 8'd74; a_mant1 = 8'd80; a_mant2 = 8'd70; a_mant3 = 8'd186;
b_mant0 = 8'd194; b_mant1 = 8'd236; b_mant2 = 8'd163; b_mant3 = 8'd135;
a_exp0 = 10'd56; a_exp1 = 10'd245; a_exp2 = 10'd313; a_exp3 = 10'd404;
b_exp0 = 10'd865; b_exp1 = 10'd812; b_exp2 = 10'd184; b_exp3 = 10'd47;
a_sign0 = 4'd16; a_sign1 = 4'd13; a_sign2 = 4'd9; a_sign3 = 4'd16;
b_sign0 = 4'd0; b_sign1 = 4'd6; b_sign2 = 4'd3; b_sign3 = 4'd4;
@(posedge clk_i);
a_mant0 = 8'd39; a_mant1 = 8'd39; a_mant2 = 8'd170; a_mant3 = 8'd204;
b_mant0 = 8'd216; b_mant1 = 8'd184; b_mant2 = 8'd31; b_mant3 = 8'd201;
a_exp0 = 10'd269; a_exp1 = 10'd809; a_exp2 = 10'd514; a_exp3 = 10'd157;
b_exp0 = 10'd763; b_exp1 = 10'd99; b_exp2 = 10'd213; b_exp3 = 10'd785;
a_sign0 = 4'd3; a_sign1 = 4'd4; a_sign2 = 4'd10; a_sign3 = 4'd5;
b_sign0 = 4'd4; b_sign1 = 4'd12; b_sign2 = 4'd14; b_sign3 = 4'd14;
@(posedge clk_i);
a_mant0 = 8'd233; a_mant1 = 8'd226; a_mant2 = 8'd189; a_mant3 = 8'd234;
b_mant0 = 8'd159; b_mant1 = 8'd63; b_mant2 = 8'd176; b_mant3 = 8'd117;
a_exp0 = 10'd0; a_exp1 = 10'd87; a_exp2 = 10'd413; a_exp3 = 10'd871;
b_exp0 = 10'd762; b_exp1 = 10'd85; b_exp2 = 10'd654; b_exp3 = 10'd230;
a_sign0 = 4'd16; a_sign1 = 4'd1; a_sign2 = 4'd6; a_sign3 = 4'd12;
b_sign0 = 4'd12; b_sign1 = 4'd6; b_sign2 = 4'd3; b_sign3 = 4'd3;
@(posedge clk_i);
a_mant0 = 8'd239; a_mant1 = 8'd159; a_mant2 = 8'd44; a_mant3 = 8'd92;
b_mant0 = 8'd124; b_mant1 = 8'd221; b_mant2 = 8'd245; b_mant3 = 8'd20;
a_exp0 = 10'd159; a_exp1 = 10'd398; a_exp2 = 10'd588; a_exp3 = 10'd434;
b_exp0 = 10'd419; b_exp1 = 10'd989; b_exp2 = 10'd27; b_exp3 = 10'd344;
a_sign0 = 4'd13; a_sign1 = 4'd6; a_sign2 = 4'd0; a_sign3 = 4'd9;
b_sign0 = 4'd0; b_sign1 = 4'd16; b_sign2 = 4'd1; b_sign3 = 4'd12;
@(posedge clk_i);
a_mant0 = 8'd20; a_mant1 = 8'd104; a_mant2 = 8'd175; a_mant3 = 8'd120;
b_mant0 = 8'd218; b_mant1 = 8'd121; b_mant2 = 8'd223; b_mant3 = 8'd15;
a_exp0 = 10'd895; a_exp1 = 10'd194; a_exp2 = 10'd448; a_exp3 = 10'd803;
b_exp0 = 10'd513; b_exp1 = 10'd405; b_exp2 = 10'd1002; b_exp3 = 10'd72;
a_sign0 = 4'd15; a_sign1 = 4'd7; a_sign2 = 4'd9; a_sign3 = 4'd16;
b_sign0 = 4'd16; b_sign1 = 4'd14; b_sign2 = 4'd16; b_sign3 = 4'd1;
@(posedge clk_i);
shared_exps0 = 8'd146;
shared_exps1 = 8'd154;
a_mant0 = 8'd208; a_mant1 = 8'd216; a_mant2 = 8'd127; a_mant3 = 8'd136;
b_mant0 = 8'd114; b_mant1 = 8'd230; b_mant2 = 8'd205; b_mant3 = 8'd180;
a_exp0 = 10'd410; a_exp1 = 10'd620; a_exp2 = 10'd608; a_exp3 = 10'd750;
b_exp0 = 10'd603; b_exp1 = 10'd638; b_exp2 = 10'd769; b_exp3 = 10'd597;
a_sign0 = 4'd15; a_sign1 = 4'd15; a_sign2 = 4'd3; a_sign3 = 4'd10;
b_sign0 = 4'd6; b_sign1 = 4'd9; b_sign2 = 4'd5; b_sign3 = 4'd11;
@(posedge clk_i);
a_mant0 = 8'd22; a_mant1 = 8'd47; a_mant2 = 8'd12; a_mant3 = 8'd56;
b_mant0 = 8'd40; b_mant1 = 8'd118; b_mant2 = 8'd186; b_mant3 = 8'd123;
a_exp0 = 10'd157; a_exp1 = 10'd863; a_exp2 = 10'd62; a_exp3 = 10'd1008;
b_exp0 = 10'd900; b_exp1 = 10'd763; b_exp2 = 10'd1004; b_exp3 = 10'd340;
a_sign0 = 4'd14; a_sign1 = 4'd10; a_sign2 = 4'd5; a_sign3 = 4'd1;
b_sign0 = 4'd10; b_sign1 = 4'd16; b_sign2 = 4'd12; b_sign3 = 4'd13;
@(posedge clk_i);
a_mant0 = 8'd181; a_mant1 = 8'd45; a_mant2 = 8'd114; a_mant3 = 8'd28;
b_mant0 = 8'd136; b_mant1 = 8'd148; b_mant2 = 8'd183; b_mant3 = 8'd18;
a_exp0 = 10'd21; a_exp1 = 10'd5; a_exp2 = 10'd164; a_exp3 = 10'd614;
b_exp0 = 10'd799; b_exp1 = 10'd20; b_exp2 = 10'd774; b_exp3 = 10'd393;
a_sign0 = 4'd4; a_sign1 = 4'd11; a_sign2 = 4'd0; a_sign3 = 4'd14;
b_sign0 = 4'd11; b_sign1 = 4'd1; b_sign2 = 4'd10; b_sign3 = 4'd14;
@(posedge clk_i);
a_mant0 = 8'd86; a_mant1 = 8'd189; a_mant2 = 8'd140; a_mant3 = 8'd234;
b_mant0 = 8'd216; b_mant1 = 8'd167; b_mant2 = 8'd149; b_mant3 = 8'd99;
a_exp0 = 10'd310; a_exp1 = 10'd130; a_exp2 = 10'd901; a_exp3 = 10'd87;
b_exp0 = 10'd289; b_exp1 = 10'd140; b_exp2 = 10'd572; b_exp3 = 10'd646;
a_sign0 = 4'd6; a_sign1 = 4'd6; a_sign2 = 4'd12; a_sign3 = 4'd3;
b_sign0 = 4'd13; b_sign1 = 4'd5; b_sign2 = 4'd16; b_sign3 = 4'd13;
@(posedge clk_i);
a_mant0 = 8'd213; a_mant1 = 8'd219; a_mant2 = 8'd244; a_mant3 = 8'd237;
b_mant0 = 8'd198; b_mant1 = 8'd136; b_mant2 = 8'd62; b_mant3 = 8'd24;
a_exp0 = 10'd982; a_exp1 = 10'd929; a_exp2 = 10'd373; a_exp3 = 10'd612;
b_exp0 = 10'd323; b_exp1 = 10'd451; b_exp2 = 10'd884; b_exp3 = 10'd265;
a_sign0 = 4'd13; a_sign1 = 4'd0; a_sign2 = 4'd3; a_sign3 = 4'd1;
b_sign0 = 4'd8; b_sign1 = 4'd1; b_sign2 = 4'd3; b_sign3 = 4'd9;
@(posedge clk_i);
a_mant0 = 8'd209; a_mant1 = 8'd115; a_mant2 = 8'd121; a_mant3 = 8'd10;
b_mant0 = 8'd38; b_mant1 = 8'd236; b_mant2 = 8'd11; b_mant3 = 8'd9;
a_exp0 = 10'd873; a_exp1 = 10'd470; a_exp2 = 10'd660; a_exp3 = 10'd553;
b_exp0 = 10'd251; b_exp1 = 10'd348; b_exp2 = 10'd638; b_exp3 = 10'd741;
a_sign0 = 4'd15; a_sign1 = 4'd4; a_sign2 = 4'd15; a_sign3 = 4'd2;
b_sign0 = 4'd4; b_sign1 = 4'd9; b_sign2 = 4'd2; b_sign3 = 4'd15;
@(posedge clk_i);
a_mant0 = 8'd121; a_mant1 = 8'd226; a_mant2 = 8'd175; a_mant3 = 8'd30;
b_mant0 = 8'd174; b_mant1 = 8'd159; b_mant2 = 8'd172; b_mant3 = 8'd149;
a_exp0 = 10'd912; a_exp1 = 10'd547; a_exp2 = 10'd595; a_exp3 = 10'd281;
b_exp0 = 10'd980; b_exp1 = 10'd141; b_exp2 = 10'd2; b_exp3 = 10'd205;
a_sign0 = 4'd10; a_sign1 = 4'd1; a_sign2 = 4'd11; a_sign3 = 4'd7;
b_sign0 = 4'd13; b_sign1 = 4'd0; b_sign2 = 4'd6; b_sign3 = 4'd14;
@(posedge clk_i);
a_mant0 = 8'd36; a_mant1 = 8'd125; a_mant2 = 8'd98; a_mant3 = 8'd114;
b_mant0 = 8'd93; b_mant1 = 8'd208; b_mant2 = 8'd4; b_mant3 = 8'd96;
a_exp0 = 10'd949; a_exp1 = 10'd871; a_exp2 = 10'd195; a_exp3 = 10'd115;
b_exp0 = 10'd765; b_exp1 = 10'd437; b_exp2 = 10'd55; b_exp3 = 10'd893;
a_sign0 = 4'd9; a_sign1 = 4'd12; a_sign2 = 4'd9; a_sign3 = 4'd8;
b_sign0 = 4'd14; b_sign1 = 4'd11; b_sign2 = 4'd10; b_sign3 = 4'd1;
@(posedge clk_i);
shared_exps0 = 8'd103;
shared_exps1 = 8'd114;
a_mant0 = 8'd21; a_mant1 = 8'd32; a_mant2 = 8'd146; a_mant3 = 8'd218;
b_mant0 = 8'd32; b_mant1 = 8'd100; b_mant2 = 8'd51; b_mant3 = 8'd31;
a_exp0 = 10'd720; a_exp1 = 10'd794; a_exp2 = 10'd285; a_exp3 = 10'd992;
b_exp0 = 10'd716; b_exp1 = 10'd596; b_exp2 = 10'd191; b_exp3 = 10'd779;
a_sign0 = 4'd4; a_sign1 = 4'd6; a_sign2 = 4'd0; a_sign3 = 4'd4;
b_sign0 = 4'd15; b_sign1 = 4'd14; b_sign2 = 4'd1; b_sign3 = 4'd12;
@(posedge clk_i);
a_mant0 = 8'd109; a_mant1 = 8'd210; a_mant2 = 8'd164; a_mant3 = 8'd13;
b_mant0 = 8'd102; b_mant1 = 8'd67; b_mant2 = 8'd223; b_mant3 = 8'd44;
a_exp0 = 10'd591; a_exp1 = 10'd1002; a_exp2 = 10'd117; a_exp3 = 10'd948;
b_exp0 = 10'd1022; b_exp1 = 10'd821; b_exp2 = 10'd1004; b_exp3 = 10'd757;
a_sign0 = 4'd15; a_sign1 = 4'd14; a_sign2 = 4'd8; a_sign3 = 4'd16;
b_sign0 = 4'd2; b_sign1 = 4'd8; b_sign2 = 4'd8; b_sign3 = 4'd3;
@(posedge clk_i);
a_mant0 = 8'd75; a_mant1 = 8'd59; a_mant2 = 8'd117; a_mant3 = 8'd133;
b_mant0 = 8'd29; b_mant1 = 8'd248; b_mant2 = 8'd179; b_mant3 = 8'd211;
a_exp0 = 10'd267; a_exp1 = 10'd72; a_exp2 = 10'd821; a_exp3 = 10'd788;
b_exp0 = 10'd22; b_exp1 = 10'd946; b_exp2 = 10'd227; b_exp3 = 10'd956;
a_sign0 = 4'd11; a_sign1 = 4'd1; a_sign2 = 4'd10; a_sign3 = 4'd9;
b_sign0 = 4'd7; b_sign1 = 4'd2; b_sign2 = 4'd11; b_sign3 = 4'd8;
@(posedge clk_i);
a_mant0 = 8'd200; a_mant1 = 8'd223; a_mant2 = 8'd143; a_mant3 = 8'd225;
b_mant0 = 8'd248; b_mant1 = 8'd21; b_mant2 = 8'd197; b_mant3 = 8'd225;
a_exp0 = 10'd191; a_exp1 = 10'd1001; a_exp2 = 10'd445; a_exp3 = 10'd192;
b_exp0 = 10'd236; b_exp1 = 10'd496; b_exp2 = 10'd918; b_exp3 = 10'd656;
a_sign0 = 4'd16; a_sign1 = 4'd3; a_sign2 = 4'd7; a_sign3 = 4'd2;
b_sign0 = 4'd9; b_sign1 = 4'd12; b_sign2 = 4'd1; b_sign3 = 4'd16;
@(posedge clk_i);
a_mant0 = 8'd143; a_mant1 = 8'd144; a_mant2 = 8'd174; a_mant3 = 8'd17;
b_mant0 = 8'd240; b_mant1 = 8'd154; b_mant2 = 8'd29; b_mant3 = 8'd96;
a_exp0 = 10'd894; a_exp1 = 10'd210; a_exp2 = 10'd440; a_exp3 = 10'd718;
b_exp0 = 10'd272; b_exp1 = 10'd990; b_exp2 = 10'd270; b_exp3 = 10'd148;
a_sign0 = 4'd15; a_sign1 = 4'd10; a_sign2 = 4'd9; a_sign3 = 4'd16;
b_sign0 = 4'd12; b_sign1 = 4'd6; b_sign2 = 4'd6; b_sign3 = 4'd2;
@(posedge clk_i);
a_mant0 = 8'd226; a_mant1 = 8'd98; a_mant2 = 8'd80; a_mant3 = 8'd58;
b_mant0 = 8'd120; b_mant1 = 8'd49; b_mant2 = 8'd5; b_mant3 = 8'd151;
a_exp0 = 10'd695; a_exp1 = 10'd672; a_exp2 = 10'd716; a_exp3 = 10'd535;
b_exp0 = 10'd199; b_exp1 = 10'd932; b_exp2 = 10'd28; b_exp3 = 10'd56;
a_sign0 = 4'd12; a_sign1 = 4'd2; a_sign2 = 4'd11; a_sign3 = 4'd9;
b_sign0 = 4'd3; b_sign1 = 4'd6; b_sign2 = 4'd4; b_sign3 = 4'd12;
@(posedge clk_i);
a_mant0 = 8'd37; a_mant1 = 8'd168; a_mant2 = 8'd169; a_mant3 = 8'd148;
b_mant0 = 8'd144; b_mant1 = 8'd181; b_mant2 = 8'd112; b_mant3 = 8'd34;
a_exp0 = 10'd955; a_exp1 = 10'd403; a_exp2 = 10'd177; a_exp3 = 10'd759;
b_exp0 = 10'd964; b_exp1 = 10'd533; b_exp2 = 10'd1016; b_exp3 = 10'd143;
a_sign0 = 4'd0; a_sign1 = 4'd14; a_sign2 = 4'd12; a_sign3 = 4'd15;
b_sign0 = 4'd6; b_sign1 = 4'd11; b_sign2 = 4'd11; b_sign3 = 4'd12;
@(posedge clk_i);
a_mant0 = 8'd168; a_mant1 = 8'd64; a_mant2 = 8'd246; a_mant3 = 8'd182;
b_mant0 = 8'd94; b_mant1 = 8'd33; b_mant2 = 8'd9; b_mant3 = 8'd196;
a_exp0 = 10'd68; a_exp1 = 10'd306; a_exp2 = 10'd776; a_exp3 = 10'd154;
b_exp0 = 10'd429; b_exp1 = 10'd529; b_exp2 = 10'd898; b_exp3 = 10'd815;
a_sign0 = 4'd9; a_sign1 = 4'd16; a_sign2 = 4'd3; a_sign3 = 4'd12;
b_sign0 = 4'd8; b_sign1 = 4'd0; b_sign2 = 4'd15; b_sign3 = 4'd0;
@(posedge clk_i);
shared_exps0 = 8'd154;
shared_exps1 = 8'd119;
rstn = 0;
@(posedge clk_i);
rstn = 1;
a_mant0 = 8'd24; a_mant1 = 8'd126; a_mant2 = 8'd65; a_mant3 = 8'd81;
b_mant0 = 8'd156; b_mant1 = 8'd36; b_mant2 = 8'd56; b_mant3 = 8'd205;
a_exp0 = 10'd925; a_exp1 = 10'd979; a_exp2 = 10'd879; a_exp3 = 10'd742;
b_exp0 = 10'd980; b_exp1 = 10'd394; b_exp2 = 10'd429; b_exp3 = 10'd258;
a_sign0 = 4'd14; a_sign1 = 4'd7; a_sign2 = 4'd16; a_sign3 = 4'd3;
b_sign0 = 4'd3; b_sign1 = 4'd1; b_sign2 = 4'd1; b_sign3 = 4'd11;
@(posedge clk_i);
a_mant0 = 8'd51; a_mant1 = 8'd102; a_mant2 = 8'd173; a_mant3 = 8'd199;
b_mant0 = 8'd46; b_mant1 = 8'd177; b_mant2 = 8'd107; b_mant3 = 8'd205;
a_exp0 = 10'd670; a_exp1 = 10'd32; a_exp2 = 10'd177; a_exp3 = 10'd564;
b_exp0 = 10'd345; b_exp1 = 10'd722; b_exp2 = 10'd224; b_exp3 = 10'd205;
a_sign0 = 4'd16; a_sign1 = 4'd16; a_sign2 = 4'd4; a_sign3 = 4'd9;
b_sign0 = 4'd9; b_sign1 = 4'd13; b_sign2 = 4'd14; b_sign3 = 4'd16;
@(posedge clk_i);
a_mant0 = 8'd169; a_mant1 = 8'd21; a_mant2 = 8'd87; a_mant3 = 8'd78;
b_mant0 = 8'd127; b_mant1 = 8'd99; b_mant2 = 8'd231; b_mant3 = 8'd90;
a_exp0 = 10'd727; a_exp1 = 10'd475; a_exp2 = 10'd100; a_exp3 = 10'd907;
b_exp0 = 10'd46; b_exp1 = 10'd379; b_exp2 = 10'd778; b_exp3 = 10'd544;
a_sign0 = 4'd7; a_sign1 = 4'd12; a_sign2 = 4'd1; a_sign3 = 4'd12;
b_sign0 = 4'd12; b_sign1 = 4'd4; b_sign2 = 4'd15; b_sign3 = 4'd7;
@(posedge clk_i);
a_mant0 = 8'd194; a_mant1 = 8'd63; a_mant2 = 8'd134; a_mant3 = 8'd162;
b_mant0 = 8'd127; b_mant1 = 8'd67; b_mant2 = 8'd1; b_mant3 = 8'd211;
a_exp0 = 10'd874; a_exp1 = 10'd123; a_exp2 = 10'd630; a_exp3 = 10'd921;
b_exp0 = 10'd172; b_exp1 = 10'd644; b_exp2 = 10'd627; b_exp3 = 10'd29;
a_sign0 = 4'd9; a_sign1 = 4'd16; a_sign2 = 4'd1; a_sign3 = 4'd14;
b_sign0 = 4'd4; b_sign1 = 4'd1; b_sign2 = 4'd8; b_sign3 = 4'd11;
@(posedge clk_i);
a_mant0 = 8'd209; a_mant1 = 8'd70; a_mant2 = 8'd224; a_mant3 = 8'd53;
b_mant0 = 8'd44; b_mant1 = 8'd84; b_mant2 = 8'd125; b_mant3 = 8'd77;
a_exp0 = 10'd498; a_exp1 = 10'd39; a_exp2 = 10'd438; a_exp3 = 10'd429;
b_exp0 = 10'd508; b_exp1 = 10'd639; b_exp2 = 10'd490; b_exp3 = 10'd939;
a_sign0 = 4'd7; a_sign1 = 4'd9; a_sign2 = 4'd15; a_sign3 = 4'd13;
b_sign0 = 4'd4; b_sign1 = 4'd1; b_sign2 = 4'd14; b_sign3 = 4'd12;
@(posedge clk_i);
a_mant0 = 8'd13; a_mant1 = 8'd223; a_mant2 = 8'd56; a_mant3 = 8'd155;
b_mant0 = 8'd75; b_mant1 = 8'd249; b_mant2 = 8'd50; b_mant3 = 8'd248;
a_exp0 = 10'd447; a_exp1 = 10'd278; a_exp2 = 10'd1009; a_exp3 = 10'd479;
b_exp0 = 10'd536; b_exp1 = 10'd571; b_exp2 = 10'd271; b_exp3 = 10'd50;
a_sign0 = 4'd8; a_sign1 = 4'd16; a_sign2 = 4'd7; a_sign3 = 4'd12;
b_sign0 = 4'd13; b_sign1 = 4'd2; b_sign2 = 4'd4; b_sign3 = 4'd13;
@(posedge clk_i);
a_mant0 = 8'd98; a_mant1 = 8'd28; a_mant2 = 8'd181; a_mant3 = 8'd177;
b_mant0 = 8'd160; b_mant1 = 8'd159; b_mant2 = 8'd99; b_mant3 = 8'd87;
a_exp0 = 10'd830; a_exp1 = 10'd883; a_exp2 = 10'd953; a_exp3 = 10'd949;
b_exp0 = 10'd719; b_exp1 = 10'd40; b_exp2 = 10'd844; b_exp3 = 10'd838;
a_sign0 = 4'd10; a_sign1 = 4'd11; a_sign2 = 4'd11; a_sign3 = 4'd0;
b_sign0 = 4'd13; b_sign1 = 4'd16; b_sign2 = 4'd15; b_sign3 = 4'd9;
@(posedge clk_i);
shared_exps0 = 8'd129;
shared_exps1 = 8'd125;
a_mant0 = 8'd74; a_mant1 = 8'd113; a_mant2 = 8'd93; a_mant3 = 8'd43;
b_mant0 = 8'd29; b_mant1 = 8'd87; b_mant2 = 8'd158; b_mant3 = 8'd228;
a_exp0 = 10'd255; a_exp1 = 10'd320; a_exp2 = 10'd230; a_exp3 = 10'd773;
b_exp0 = 10'd890; b_exp1 = 10'd18; b_exp2 = 10'd276; b_exp3 = 10'd68;
a_sign0 = 4'd5; a_sign1 = 4'd1; a_sign2 = 4'd8; a_sign3 = 4'd3;
b_sign0 = 4'd5; b_sign1 = 4'd9; b_sign2 = 4'd12; b_sign3 = 4'd3;
@(posedge clk_i);
a_mant0 = 8'd98; a_mant1 = 8'd108; a_mant2 = 8'd139; a_mant3 = 8'd155;
b_mant0 = 8'd199; b_mant1 = 8'd140; b_mant2 = 8'd77; b_mant3 = 8'd182;
a_exp0 = 10'd498; a_exp1 = 10'd212; a_exp2 = 10'd576; a_exp3 = 10'd494;
b_exp0 = 10'd456; b_exp1 = 10'd100; b_exp2 = 10'd431; b_exp3 = 10'd662;
a_sign0 = 4'd4; a_sign1 = 4'd12; a_sign2 = 4'd3; a_sign3 = 4'd14;
b_sign0 = 4'd14; b_sign1 = 4'd9; b_sign2 = 4'd10; b_sign3 = 4'd13;
@(posedge clk_i);
a_mant0 = 8'd75; a_mant1 = 8'd129; a_mant2 = 8'd14; a_mant3 = 8'd73;
b_mant0 = 8'd159; b_mant1 = 8'd103; b_mant2 = 8'd75; b_mant3 = 8'd85;
a_exp0 = 10'd906; a_exp1 = 10'd620; a_exp2 = 10'd405; a_exp3 = 10'd135;
b_exp0 = 10'd311; b_exp1 = 10'd145; b_exp2 = 10'd768; b_exp3 = 10'd79;
a_sign0 = 4'd16; a_sign1 = 4'd5; a_sign2 = 4'd11; a_sign3 = 4'd5;
b_sign0 = 4'd8; b_sign1 = 4'd10; b_sign2 = 4'd0; b_sign3 = 4'd8;
@(posedge clk_i);
a_mant0 = 8'd153; a_mant1 = 8'd8; a_mant2 = 8'd156; a_mant3 = 8'd49;
b_mant0 = 8'd223; b_mant1 = 8'd158; b_mant2 = 8'd62; b_mant3 = 8'd209;
a_exp0 = 10'd1004; a_exp1 = 10'd25; a_exp2 = 10'd144; a_exp3 = 10'd445;
b_exp0 = 10'd283; b_exp1 = 10'd969; b_exp2 = 10'd779; b_exp3 = 10'd548;
a_sign0 = 4'd14; a_sign1 = 4'd16; a_sign2 = 4'd10; a_sign3 = 4'd13;
b_sign0 = 4'd15; b_sign1 = 4'd16; b_sign2 = 4'd15; b_sign3 = 4'd0;
@(posedge clk_i);
a_mant0 = 8'd35; a_mant1 = 8'd223; a_mant2 = 8'd235; a_mant3 = 8'd95;
b_mant0 = 8'd1; b_mant1 = 8'd13; b_mant2 = 8'd23; b_mant3 = 8'd137;
a_exp0 = 10'd69; a_exp1 = 10'd388; a_exp2 = 10'd545; a_exp3 = 10'd13;
b_exp0 = 10'd1017; b_exp1 = 10'd963; b_exp2 = 10'd29; b_exp3 = 10'd423;
a_sign0 = 4'd6; a_sign1 = 4'd5; a_sign2 = 4'd1; a_sign3 = 4'd10;
b_sign0 = 4'd13; b_sign1 = 4'd9; b_sign2 = 4'd10; b_sign3 = 4'd4;
@(posedge clk_i);
a_mant0 = 8'd43; a_mant1 = 8'd196; a_mant2 = 8'd22; a_mant3 = 8'd188;
b_mant0 = 8'd229; b_mant1 = 8'd153; b_mant2 = 8'd22; b_mant3 = 8'd116;
a_exp0 = 10'd807; a_exp1 = 10'd676; a_exp2 = 10'd325; a_exp3 = 10'd559;
b_exp0 = 10'd933; b_exp1 = 10'd971; b_exp2 = 10'd71; b_exp3 = 10'd843;
a_sign0 = 4'd10; a_sign1 = 4'd10; a_sign2 = 4'd2; a_sign3 = 4'd1;
b_sign0 = 4'd15; b_sign1 = 4'd9; b_sign2 = 4'd10; b_sign3 = 4'd6;
@(posedge clk_i);
a_mant0 = 8'd213; a_mant1 = 8'd88; a_mant2 = 8'd181; a_mant3 = 8'd68;
b_mant0 = 8'd218; b_mant1 = 8'd225; b_mant2 = 8'd210; b_mant3 = 8'd143;
a_exp0 = 10'd150; a_exp1 = 10'd721; a_exp2 = 10'd932; a_exp3 = 10'd695;
b_exp0 = 10'd996; b_exp1 = 10'd257; b_exp2 = 10'd64; b_exp3 = 10'd138;
a_sign0 = 4'd1; a_sign1 = 4'd6; a_sign2 = 4'd3; a_sign3 = 4'd2;
b_sign0 = 4'd14; b_sign1 = 4'd5; b_sign2 = 4'd1; b_sign3 = 4'd14;
@(posedge clk_i);
a_mant0 = 8'd243; a_mant1 = 8'd142; a_mant2 = 8'd79; a_mant3 = 8'd224;
b_mant0 = 8'd114; b_mant1 = 8'd251; b_mant2 = 8'd22; b_mant3 = 8'd212;
a_exp0 = 10'd532; a_exp1 = 10'd120; a_exp2 = 10'd814; a_exp3 = 10'd1022;
b_exp0 = 10'd204; b_exp1 = 10'd795; b_exp2 = 10'd754; b_exp3 = 10'd199;
a_sign0 = 4'd16; a_sign1 = 4'd3; a_sign2 = 4'd16; a_sign3 = 4'd0;
b_sign0 = 4'd9; b_sign1 = 4'd8; b_sign2 = 4'd7; b_sign3 = 4'd6;
@(posedge clk_i);
shared_exps0 = 8'd141;
shared_exps1 = 8'd118;
a_mant0 = 8'd141; a_mant1 = 8'd170; a_mant2 = 8'd58; a_mant3 = 8'd193;
b_mant0 = 8'd95; b_mant1 = 8'd6; b_mant2 = 8'd89; b_mant3 = 8'd232;
a_exp0 = 10'd398; a_exp1 = 10'd917; a_exp2 = 10'd599; a_exp3 = 10'd900;
b_exp0 = 10'd759; b_exp1 = 10'd289; b_exp2 = 10'd288; b_exp3 = 10'd609;
a_sign0 = 4'd11; a_sign1 = 4'd11; a_sign2 = 4'd11; a_sign3 = 4'd15;
b_sign0 = 4'd8; b_sign1 = 4'd15; b_sign2 = 4'd14; b_sign3 = 4'd8;
@(posedge clk_i);
a_mant0 = 8'd253; a_mant1 = 8'd57; a_mant2 = 8'd85; a_mant3 = 8'd67;
b_mant0 = 8'd205; b_mant1 = 8'd168; b_mant2 = 8'd240; b_mant3 = 8'd117;
a_exp0 = 10'd325; a_exp1 = 10'd418; a_exp2 = 10'd272; a_exp3 = 10'd71;
b_exp0 = 10'd921; b_exp1 = 10'd856; b_exp2 = 10'd650; b_exp3 = 10'd95;
a_sign0 = 4'd13; a_sign1 = 4'd8; a_sign2 = 4'd9; a_sign3 = 4'd1;
b_sign0 = 4'd12; b_sign1 = 4'd9; b_sign2 = 4'd5; b_sign3 = 4'd4;
@(posedge clk_i);
a_mant0 = 8'd115; a_mant1 = 8'd196; a_mant2 = 8'd166; a_mant3 = 8'd151;
b_mant0 = 8'd135; b_mant1 = 8'd221; b_mant2 = 8'd6; b_mant3 = 8'd174;
a_exp0 = 10'd890; a_exp1 = 10'd975; a_exp2 = 10'd9; a_exp3 = 10'd948;
b_exp0 = 10'd850; b_exp1 = 10'd644; b_exp2 = 10'd84; b_exp3 = 10'd969;
a_sign0 = 4'd13; a_sign1 = 4'd10; a_sign2 = 4'd6; a_sign3 = 4'd11;
b_sign0 = 4'd11; b_sign1 = 4'd10; b_sign2 = 4'd16; b_sign3 = 4'd12;
@(posedge clk_i);
a_mant0 = 8'd110; a_mant1 = 8'd197; a_mant2 = 8'd68; a_mant3 = 8'd66;
b_mant0 = 8'd230; b_mant1 = 8'd104; b_mant2 = 8'd133; b_mant3 = 8'd88;
a_exp0 = 10'd583; a_exp1 = 10'd99; a_exp2 = 10'd481; a_exp3 = 10'd11;
b_exp0 = 10'd779; b_exp1 = 10'd515; b_exp2 = 10'd318; b_exp3 = 10'd253;
a_sign0 = 4'd10; a_sign1 = 4'd5; a_sign2 = 4'd16; a_sign3 = 4'd1;
b_sign0 = 4'd7; b_sign1 = 4'd3; b_sign2 = 4'd1; b_sign3 = 4'd11;
@(posedge clk_i);
a_mant0 = 8'd238; a_mant1 = 8'd159; a_mant2 = 8'd162; a_mant3 = 8'd93;
b_mant0 = 8'd64; b_mant1 = 8'd182; b_mant2 = 8'd205; b_mant3 = 8'd108;
a_exp0 = 10'd244; a_exp1 = 10'd572; a_exp2 = 10'd129; a_exp3 = 10'd996;
b_exp0 = 10'd25; b_exp1 = 10'd22; b_exp2 = 10'd946; b_exp3 = 10'd385;
a_sign0 = 4'd3; a_sign1 = 4'd0; a_sign2 = 4'd3; a_sign3 = 4'd14;
b_sign0 = 4'd14; b_sign1 = 4'd10; b_sign2 = 4'd8; b_sign3 = 4'd16;
@(posedge clk_i);
a_mant0 = 8'd178; a_mant1 = 8'd207; a_mant2 = 8'd217; a_mant3 = 8'd226;
b_mant0 = 8'd67; b_mant1 = 8'd3; b_mant2 = 8'd157; b_mant3 = 8'd169;
a_exp0 = 10'd619; a_exp1 = 10'd530; a_exp2 = 10'd832; a_exp3 = 10'd918;
b_exp0 = 10'd822; b_exp1 = 10'd679; b_exp2 = 10'd957; b_exp3 = 10'd616;
a_sign0 = 4'd14; a_sign1 = 4'd7; a_sign2 = 4'd14; a_sign3 = 4'd7;
b_sign0 = 4'd0; b_sign1 = 4'd11; b_sign2 = 4'd0; b_sign3 = 4'd4;
@(posedge clk_i);
a_mant0 = 8'd4; a_mant1 = 8'd163; a_mant2 = 8'd34; a_mant3 = 8'd26;
b_mant0 = 8'd112; b_mant1 = 8'd135; b_mant2 = 8'd155; b_mant3 = 8'd21;
a_exp0 = 10'd487; a_exp1 = 10'd40; a_exp2 = 10'd158; a_exp3 = 10'd438;
b_exp0 = 10'd826; b_exp1 = 10'd596; b_exp2 = 10'd860; b_exp3 = 10'd732;
a_sign0 = 4'd4; a_sign1 = 4'd14; a_sign2 = 4'd3; a_sign3 = 4'd13;
b_sign0 = 4'd8; b_sign1 = 4'd6; b_sign2 = 4'd2; b_sign3 = 4'd7;
@(posedge clk_i);
a_mant0 = 8'd3; a_mant1 = 8'd57; a_mant2 = 8'd27; a_mant3 = 8'd195;
b_mant0 = 8'd116; b_mant1 = 8'd206; b_mant2 = 8'd100; b_mant3 = 8'd47;
a_exp0 = 10'd411; a_exp1 = 10'd850; a_exp2 = 10'd834; a_exp3 = 10'd596;
b_exp0 = 10'd114; b_exp1 = 10'd742; b_exp2 = 10'd264; b_exp3 = 10'd266;
a_sign0 = 4'd6; a_sign1 = 4'd4; a_sign2 = 4'd13; a_sign3 = 4'd10;
b_sign0 = 4'd9; b_sign1 = 4'd4; b_sign2 = 4'd12; b_sign3 = 4'd6;
@(posedge clk_i);
shared_exps0 = 8'd109;
shared_exps1 = 8'd130;
a_mant0 = 8'd102; a_mant1 = 8'd50; a_mant2 = 8'd185; a_mant3 = 8'd237;
b_mant0 = 8'd216; b_mant1 = 8'd68; b_mant2 = 8'd184; b_mant3 = 8'd20;
a_exp0 = 10'd664; a_exp1 = 10'd24; a_exp2 = 10'd473; a_exp3 = 10'd154;
b_exp0 = 10'd768; b_exp1 = 10'd748; b_exp2 = 10'd247; b_exp3 = 10'd200;
a_sign0 = 4'd13; a_sign1 = 4'd1; a_sign2 = 4'd4; a_sign3 = 4'd2;
b_sign0 = 4'd2; b_sign1 = 4'd9; b_sign2 = 4'd3; b_sign3 = 4'd7;
@(posedge clk_i);
a_mant0 = 8'd6; a_mant1 = 8'd199; a_mant2 = 8'd152; a_mant3 = 8'd225;
b_mant0 = 8'd166; b_mant1 = 8'd250; b_mant2 = 8'd38; b_mant3 = 8'd112;
a_exp0 = 10'd633; a_exp1 = 10'd702; a_exp2 = 10'd472; a_exp3 = 10'd922;
b_exp0 = 10'd277; b_exp1 = 10'd855; b_exp2 = 10'd519; b_exp3 = 10'd917;
a_sign0 = 4'd16; a_sign1 = 4'd9; a_sign2 = 4'd6; a_sign3 = 4'd1;
b_sign0 = 4'd8; b_sign1 = 4'd10; b_sign2 = 4'd12; b_sign3 = 4'd2;
@(posedge clk_i);
a_mant0 = 8'd198; a_mant1 = 8'd163; a_mant2 = 8'd252; a_mant3 = 8'd14;
b_mant0 = 8'd189; b_mant1 = 8'd52; b_mant2 = 8'd155; b_mant3 = 8'd109;
a_exp0 = 10'd285; a_exp1 = 10'd1; a_exp2 = 10'd665; a_exp3 = 10'd55;
b_exp0 = 10'd869; b_exp1 = 10'd938; b_exp2 = 10'd189; b_exp3 = 10'd250;
a_sign0 = 4'd2; a_sign1 = 4'd11; a_sign2 = 4'd12; a_sign3 = 4'd5;
b_sign0 = 4'd1; b_sign1 = 4'd12; b_sign2 = 4'd15; b_sign3 = 4'd16;
@(posedge clk_i);
a_mant0 = 8'd156; a_mant1 = 8'd211; a_mant2 = 8'd124; a_mant3 = 8'd19;
b_mant0 = 8'd195; b_mant1 = 8'd58; b_mant2 = 8'd96; b_mant3 = 8'd130;
a_exp0 = 10'd705; a_exp1 = 10'd418; a_exp2 = 10'd649; a_exp3 = 10'd154;
b_exp0 = 10'd729; b_exp1 = 10'd72; b_exp2 = 10'd134; b_exp3 = 10'd377;
a_sign0 = 4'd0; a_sign1 = 4'd5; a_sign2 = 4'd9; a_sign3 = 4'd8;
b_sign0 = 4'd7; b_sign1 = 4'd9; b_sign2 = 4'd6; b_sign3 = 4'd4;
@(posedge clk_i);
a_mant0 = 8'd181; a_mant1 = 8'd146; a_mant2 = 8'd11; a_mant3 = 8'd166;
b_mant0 = 8'd81; b_mant1 = 8'd220; b_mant2 = 8'd152; b_mant3 = 8'd149;
a_exp0 = 10'd328; a_exp1 = 10'd737; a_exp2 = 10'd509; a_exp3 = 10'd67;
b_exp0 = 10'd501; b_exp1 = 10'd338; b_exp2 = 10'd979; b_exp3 = 10'd1012;
a_sign0 = 4'd6; a_sign1 = 4'd13; a_sign2 = 4'd8; a_sign3 = 4'd8;
b_sign0 = 4'd6; b_sign1 = 4'd2; b_sign2 = 4'd16; b_sign3 = 4'd3;
@(posedge clk_i);
a_mant0 = 8'd46; a_mant1 = 8'd231; a_mant2 = 8'd246; a_mant3 = 8'd214;
b_mant0 = 8'd179; b_mant1 = 8'd186; b_mant2 = 8'd222; b_mant3 = 8'd148;
a_exp0 = 10'd218; a_exp1 = 10'd785; a_exp2 = 10'd839; a_exp3 = 10'd761;
b_exp0 = 10'd506; b_exp1 = 10'd868; b_exp2 = 10'd592; b_exp3 = 10'd388;
a_sign0 = 4'd12; a_sign1 = 4'd2; a_sign2 = 4'd0; a_sign3 = 4'd11;
b_sign0 = 4'd1; b_sign1 = 4'd9; b_sign2 = 4'd14; b_sign3 = 4'd3;
@(posedge clk_i);
a_mant0 = 8'd103; a_mant1 = 8'd249; a_mant2 = 8'd121; a_mant3 = 8'd33;
b_mant0 = 8'd167; b_mant1 = 8'd47; b_mant2 = 8'd161; b_mant3 = 8'd71;
a_exp0 = 10'd173; a_exp1 = 10'd48; a_exp2 = 10'd993; a_exp3 = 10'd696;
b_exp0 = 10'd209; b_exp1 = 10'd85; b_exp2 = 10'd512; b_exp3 = 10'd1021;
a_sign0 = 4'd8; a_sign1 = 4'd2; a_sign2 = 4'd3; a_sign3 = 4'd2;
b_sign0 = 4'd13; b_sign1 = 4'd11; b_sign2 = 4'd10; b_sign3 = 4'd9;
@(posedge clk_i);
a_mant0 = 8'd35; a_mant1 = 8'd38; a_mant2 = 8'd30; a_mant3 = 8'd69;
b_mant0 = 8'd177; b_mant1 = 8'd156; b_mant2 = 8'd11; b_mant3 = 8'd152;
a_exp0 = 10'd1015; a_exp1 = 10'd866; a_exp2 = 10'd9; a_exp3 = 10'd721;
b_exp0 = 10'd492; b_exp1 = 10'd414; b_exp2 = 10'd945; b_exp3 = 10'd855;
a_sign0 = 4'd1; a_sign1 = 4'd13; a_sign2 = 4'd14; a_sign3 = 4'd16;
b_sign0 = 4'd7; b_sign1 = 4'd10; b_sign2 = 4'd8; b_sign3 = 4'd4;
@(posedge clk_i);
shared_exps0 = 8'd157;
shared_exps1 = 8'd140;
rstn = 0;
@(posedge clk_i);
rstn = 1;
a_mant0 = 8'd134; a_mant1 = 8'd122; a_mant2 = 8'd165; a_mant3 = 8'd80;
b_mant0 = 8'd108; b_mant1 = 8'd111; b_mant2 = 8'd24; b_mant3 = 8'd99;
a_exp0 = 10'd573; a_exp1 = 10'd140; a_exp2 = 10'd689; a_exp3 = 10'd659;
b_exp0 = 10'd508; b_exp1 = 10'd945; b_exp2 = 10'd131; b_exp3 = 10'd111;
a_sign0 = 4'd10; a_sign1 = 4'd5; a_sign2 = 4'd5; a_sign3 = 4'd13;
b_sign0 = 4'd7; b_sign1 = 4'd0; b_sign2 = 4'd1; b_sign3 = 4'd13;
@(posedge clk_i);
a_mant0 = 8'd62; a_mant1 = 8'd129; a_mant2 = 8'd102; a_mant3 = 8'd178;
b_mant0 = 8'd76; b_mant1 = 8'd88; b_mant2 = 8'd70; b_mant3 = 8'd198;
a_exp0 = 10'd182; a_exp1 = 10'd424; a_exp2 = 10'd446; a_exp3 = 10'd431;
b_exp0 = 10'd938; b_exp1 = 10'd243; b_exp2 = 10'd83; b_exp3 = 10'd532;
a_sign0 = 4'd11; a_sign1 = 4'd10; a_sign2 = 4'd4; a_sign3 = 4'd3;
b_sign0 = 4'd1; b_sign1 = 4'd15; b_sign2 = 4'd11; b_sign3 = 4'd10;
@(posedge clk_i);
a_mant0 = 8'd240; a_mant1 = 8'd123; a_mant2 = 8'd105; a_mant3 = 8'd47;
b_mant0 = 8'd143; b_mant1 = 8'd142; b_mant2 = 8'd176; b_mant3 = 8'd53;
a_exp0 = 10'd77; a_exp1 = 10'd892; a_exp2 = 10'd389; a_exp3 = 10'd1018;
b_exp0 = 10'd608; b_exp1 = 10'd751; b_exp2 = 10'd901; b_exp3 = 10'd786;
a_sign0 = 4'd13; a_sign1 = 4'd16; a_sign2 = 4'd1; a_sign3 = 4'd3;
b_sign0 = 4'd15; b_sign1 = 4'd0; b_sign2 = 4'd1; b_sign3 = 4'd6;
@(posedge clk_i);
a_mant0 = 8'd120; a_mant1 = 8'd249; a_mant2 = 8'd62; a_mant3 = 8'd31;
b_mant0 = 8'd186; b_mant1 = 8'd58; b_mant2 = 8'd232; b_mant3 = 8'd77;
a_exp0 = 10'd150; a_exp1 = 10'd596; a_exp2 = 10'd978; a_exp3 = 10'd54;
b_exp0 = 10'd108; b_exp1 = 10'd287; b_exp2 = 10'd87; b_exp3 = 10'd350;
a_sign0 = 4'd2; a_sign1 = 4'd0; a_sign2 = 4'd0; a_sign3 = 4'd15;
b_sign0 = 4'd2; b_sign1 = 4'd2; b_sign2 = 4'd2; b_sign3 = 4'd10;
@(posedge clk_i);
a_mant0 = 8'd112; a_mant1 = 8'd91; a_mant2 = 8'd1; a_mant3 = 8'd82;
b_mant0 = 8'd212; b_mant1 = 8'd113; b_mant2 = 8'd74; b_mant3 = 8'd66;
a_exp0 = 10'd869; a_exp1 = 10'd935; a_exp2 = 10'd94; a_exp3 = 10'd707;
b_exp0 = 10'd694; b_exp1 = 10'd214; b_exp2 = 10'd722; b_exp3 = 10'd637;
a_sign0 = 4'd4; a_sign1 = 4'd8; a_sign2 = 4'd1; a_sign3 = 4'd11;
b_sign0 = 4'd15; b_sign1 = 4'd12; b_sign2 = 4'd16; b_sign3 = 4'd2;
@(posedge clk_i);
a_mant0 = 8'd8; a_mant1 = 8'd47; a_mant2 = 8'd197; a_mant3 = 8'd224;
b_mant0 = 8'd245; b_mant1 = 8'd216; b_mant2 = 8'd121; b_mant3 = 8'd58;
a_exp0 = 10'd841; a_exp1 = 10'd789; a_exp2 = 10'd506; a_exp3 = 10'd447;
b_exp0 = 10'd386; b_exp1 = 10'd436; b_exp2 = 10'd934; b_exp3 = 10'd924;
a_sign0 = 4'd7; a_sign1 = 4'd3; a_sign2 = 4'd1; a_sign3 = 4'd11;
b_sign0 = 4'd14; b_sign1 = 4'd14; b_sign2 = 4'd3; b_sign3 = 4'd7;
@(posedge clk_i);
a_mant0 = 8'd25; a_mant1 = 8'd73; a_mant2 = 8'd143; a_mant3 = 8'd75;
b_mant0 = 8'd28; b_mant1 = 8'd235; b_mant2 = 8'd40; b_mant3 = 8'd244;
a_exp0 = 10'd382; a_exp1 = 10'd919; a_exp2 = 10'd792; a_exp3 = 10'd744;
b_exp0 = 10'd938; b_exp1 = 10'd408; b_exp2 = 10'd372; b_exp3 = 10'd529;
a_sign0 = 4'd16; a_sign1 = 4'd11; a_sign2 = 4'd16; a_sign3 = 4'd15;
b_sign0 = 4'd10; b_sign1 = 4'd12; b_sign2 = 4'd8; b_sign3 = 4'd10;
@(posedge clk_i);
shared_exps0 = 8'd109;
shared_exps1 = 8'd151;
a_mant0 = 8'd4; a_mant1 = 8'd113; a_mant2 = 8'd25; a_mant3 = 8'd131;
b_mant0 = 8'd8; b_mant1 = 8'd136; b_mant2 = 8'd15; b_mant3 = 8'd56;
a_exp0 = 10'd280; a_exp1 = 10'd894; a_exp2 = 10'd693; a_exp3 = 10'd482;
b_exp0 = 10'd636; b_exp1 = 10'd920; b_exp2 = 10'd206; b_exp3 = 10'd56;
a_sign0 = 4'd4; a_sign1 = 4'd11; a_sign2 = 4'd1; a_sign3 = 4'd4;
b_sign0 = 4'd4; b_sign1 = 4'd11; b_sign2 = 4'd9; b_sign3 = 4'd16;
@(posedge clk_i);
a_mant0 = 8'd73; a_mant1 = 8'd246; a_mant2 = 8'd60; a_mant3 = 8'd231;
b_mant0 = 8'd148; b_mant1 = 8'd198; b_mant2 = 8'd33; b_mant3 = 8'd214;
a_exp0 = 10'd609; a_exp1 = 10'd326; a_exp2 = 10'd500; a_exp3 = 10'd7;
b_exp0 = 10'd999; b_exp1 = 10'd163; b_exp2 = 10'd309; b_exp3 = 10'd179;
a_sign0 = 4'd15; a_sign1 = 4'd0; a_sign2 = 4'd14; a_sign3 = 4'd13;
b_sign0 = 4'd6; b_sign1 = 4'd10; b_sign2 = 4'd4; b_sign3 = 4'd13;
@(posedge clk_i);
a_mant0 = 8'd172; a_mant1 = 8'd34; a_mant2 = 8'd86; a_mant3 = 8'd146;
b_mant0 = 8'd125; b_mant1 = 8'd181; b_mant2 = 8'd44; b_mant3 = 8'd246;
a_exp0 = 10'd766; a_exp1 = 10'd145; a_exp2 = 10'd75; a_exp3 = 10'd359;
b_exp0 = 10'd606; b_exp1 = 10'd729; b_exp2 = 10'd950; b_exp3 = 10'd101;
a_sign0 = 4'd7; a_sign1 = 4'd16; a_sign2 = 4'd11; a_sign3 = 4'd4;
b_sign0 = 4'd4; b_sign1 = 4'd15; b_sign2 = 4'd1; b_sign3 = 4'd0;
@(posedge clk_i);
a_mant0 = 8'd18; a_mant1 = 8'd147; a_mant2 = 8'd141; a_mant3 = 8'd101;
b_mant0 = 8'd186; b_mant1 = 8'd119; b_mant2 = 8'd202; b_mant3 = 8'd200;
a_exp0 = 10'd53; a_exp1 = 10'd471; a_exp2 = 10'd509; a_exp3 = 10'd429;
b_exp0 = 10'd524; b_exp1 = 10'd929; b_exp2 = 10'd558; b_exp3 = 10'd946;
a_sign0 = 4'd0; a_sign1 = 4'd5; a_sign2 = 4'd9; a_sign3 = 4'd15;
b_sign0 = 4'd14; b_sign1 = 4'd15; b_sign2 = 4'd15; b_sign3 = 4'd12;
@(posedge clk_i);
a_mant0 = 8'd221; a_mant1 = 8'd108; a_mant2 = 8'd66; a_mant3 = 8'd62;
b_mant0 = 8'd241; b_mant1 = 8'd16; b_mant2 = 8'd15; b_mant3 = 8'd181;
a_exp0 = 10'd47; a_exp1 = 10'd718; a_exp2 = 10'd49; a_exp3 = 10'd46;
b_exp0 = 10'd278; b_exp1 = 10'd326; b_exp2 = 10'd317; b_exp3 = 10'd553;
a_sign0 = 4'd2; a_sign1 = 4'd5; a_sign2 = 4'd11; a_sign3 = 4'd13;
b_sign0 = 4'd13; b_sign1 = 4'd6; b_sign2 = 4'd13; b_sign3 = 4'd12;
@(posedge clk_i);
a_mant0 = 8'd0; a_mant1 = 8'd249; a_mant2 = 8'd90; a_mant3 = 8'd58;
b_mant0 = 8'd17; b_mant1 = 8'd53; b_mant2 = 8'd85; b_mant3 = 8'd45;
a_exp0 = 10'd1003; a_exp1 = 10'd962; a_exp2 = 10'd427; a_exp3 = 10'd770;
b_exp0 = 10'd852; b_exp1 = 10'd975; b_exp2 = 10'd837; b_exp3 = 10'd657;
a_sign0 = 4'd5; a_sign1 = 4'd9; a_sign2 = 4'd5; a_sign3 = 4'd5;
b_sign0 = 4'd5; b_sign1 = 4'd8; b_sign2 = 4'd7; b_sign3 = 4'd7;
@(posedge clk_i);
a_mant0 = 8'd103; a_mant1 = 8'd248; a_mant2 = 8'd221; a_mant3 = 8'd81;
b_mant0 = 8'd83; b_mant1 = 8'd161; b_mant2 = 8'd100; b_mant3 = 8'd59;
a_exp0 = 10'd106; a_exp1 = 10'd448; a_exp2 = 10'd709; a_exp3 = 10'd958;
b_exp0 = 10'd681; b_exp1 = 10'd472; b_exp2 = 10'd926; b_exp3 = 10'd36;
a_sign0 = 4'd9; a_sign1 = 4'd9; a_sign2 = 4'd13; a_sign3 = 4'd2;
b_sign0 = 4'd5; b_sign1 = 4'd16; b_sign2 = 4'd16; b_sign3 = 4'd0;
@(posedge clk_i);
a_mant0 = 8'd195; a_mant1 = 8'd131; a_mant2 = 8'd65; a_mant3 = 8'd109;
b_mant0 = 8'd59; b_mant1 = 8'd202; b_mant2 = 8'd11; b_mant3 = 8'd112;
a_exp0 = 10'd194; a_exp1 = 10'd122; a_exp2 = 10'd758; a_exp3 = 10'd912;
b_exp0 = 10'd171; b_exp1 = 10'd456; b_exp2 = 10'd40; b_exp3 = 10'd922;
a_sign0 = 4'd2; a_sign1 = 4'd6; a_sign2 = 4'd7; a_sign3 = 4'd10;
b_sign0 = 4'd16; b_sign1 = 4'd4; b_sign2 = 4'd10; b_sign3 = 4'd1;
@(posedge clk_i);
shared_exps0 = 8'd133;
shared_exps1 = 8'd144;
a_mant0 = 8'd160; a_mant1 = 8'd83; a_mant2 = 8'd44; a_mant3 = 8'd236;
b_mant0 = 8'd116; b_mant1 = 8'd212; b_mant2 = 8'd118; b_mant3 = 8'd174;
a_exp0 = 10'd197; a_exp1 = 10'd668; a_exp2 = 10'd228; a_exp3 = 10'd1004;
b_exp0 = 10'd318; b_exp1 = 10'd713; b_exp2 = 10'd216; b_exp3 = 10'd95;
a_sign0 = 4'd9; a_sign1 = 4'd5; a_sign2 = 4'd5; a_sign3 = 4'd9;
b_sign0 = 4'd13; b_sign1 = 4'd1; b_sign2 = 4'd0; b_sign3 = 4'd5;
@(posedge clk_i);
a_mant0 = 8'd99; a_mant1 = 8'd246; a_mant2 = 8'd15; a_mant3 = 8'd29;
b_mant0 = 8'd221; b_mant1 = 8'd199; b_mant2 = 8'd200; b_mant3 = 8'd140;
a_exp0 = 10'd974; a_exp1 = 10'd266; a_exp2 = 10'd87; a_exp3 = 10'd625;
b_exp0 = 10'd601; b_exp1 = 10'd85; b_exp2 = 10'd392; b_exp3 = 10'd560;
a_sign0 = 4'd14; a_sign1 = 4'd10; a_sign2 = 4'd10; a_sign3 = 4'd2;
b_sign0 = 4'd14; b_sign1 = 4'd2; b_sign2 = 4'd10; b_sign3 = 4'd8;
@(posedge clk_i);
a_mant0 = 8'd177; a_mant1 = 8'd0; a_mant2 = 8'd157; a_mant3 = 8'd89;
b_mant0 = 8'd30; b_mant1 = 8'd169; b_mant2 = 8'd46; b_mant3 = 8'd16;
a_exp0 = 10'd338; a_exp1 = 10'd406; a_exp2 = 10'd377; a_exp3 = 10'd509;
b_exp0 = 10'd147; b_exp1 = 10'd53; b_exp2 = 10'd539; b_exp3 = 10'd329;
a_sign0 = 4'd13; a_sign1 = 4'd1; a_sign2 = 4'd7; a_sign3 = 4'd1;
b_sign0 = 4'd2; b_sign1 = 4'd10; b_sign2 = 4'd13; b_sign3 = 4'd5;
@(posedge clk_i);
a_mant0 = 8'd232; a_mant1 = 8'd169; a_mant2 = 8'd153; a_mant3 = 8'd58;
b_mant0 = 8'd61; b_mant1 = 8'd197; b_mant2 = 8'd176; b_mant3 = 8'd18;
a_exp0 = 10'd590; a_exp1 = 10'd5; a_exp2 = 10'd1002; a_exp3 = 10'd155;
b_exp0 = 10'd508; b_exp1 = 10'd156; b_exp2 = 10'd454; b_exp3 = 10'd97;
a_sign0 = 4'd16; a_sign1 = 4'd13; a_sign2 = 4'd3; a_sign3 = 4'd3;
b_sign0 = 4'd14; b_sign1 = 4'd14; b_sign2 = 4'd5; b_sign3 = 4'd4;
@(posedge clk_i);
a_mant0 = 8'd146; a_mant1 = 8'd130; a_mant2 = 8'd194; a_mant3 = 8'd212;
b_mant0 = 8'd59; b_mant1 = 8'd208; b_mant2 = 8'd11; b_mant3 = 8'd211;
a_exp0 = 10'd369; a_exp1 = 10'd87; a_exp2 = 10'd136; a_exp3 = 10'd615;
b_exp0 = 10'd425; b_exp1 = 10'd534; b_exp2 = 10'd986; b_exp3 = 10'd117;
a_sign0 = 4'd2; a_sign1 = 4'd15; a_sign2 = 4'd16; a_sign3 = 4'd11;
b_sign0 = 4'd11; b_sign1 = 4'd9; b_sign2 = 4'd3; b_sign3 = 4'd6;
@(posedge clk_i);
a_mant0 = 8'd228; a_mant1 = 8'd178; a_mant2 = 8'd140; a_mant3 = 8'd194;
b_mant0 = 8'd157; b_mant1 = 8'd169; b_mant2 = 8'd92; b_mant3 = 8'd99;
a_exp0 = 10'd253; a_exp1 = 10'd421; a_exp2 = 10'd1014; a_exp3 = 10'd568;
b_exp0 = 10'd183; b_exp1 = 10'd306; b_exp2 = 10'd502; b_exp3 = 10'd156;
a_sign0 = 4'd9; a_sign1 = 4'd3; a_sign2 = 4'd9; a_sign3 = 4'd9;
b_sign0 = 4'd7; b_sign1 = 4'd13; b_sign2 = 4'd7; b_sign3 = 4'd0;
@(posedge clk_i);
a_mant0 = 8'd204; a_mant1 = 8'd206; a_mant2 = 8'd235; a_mant3 = 8'd79;
b_mant0 = 8'd135; b_mant1 = 8'd158; b_mant2 = 8'd34; b_mant3 = 8'd142;
a_exp0 = 10'd334; a_exp1 = 10'd341; a_exp2 = 10'd344; a_exp3 = 10'd765;
b_exp0 = 10'd463; b_exp1 = 10'd962; b_exp2 = 10'd959; b_exp3 = 10'd855;
a_sign0 = 4'd4; a_sign1 = 4'd16; a_sign2 = 4'd2; a_sign3 = 4'd12;
b_sign0 = 4'd13; b_sign1 = 4'd6; b_sign2 = 4'd11; b_sign3 = 4'd5;
@(posedge clk_i);
a_mant0 = 8'd164; a_mant1 = 8'd63; a_mant2 = 8'd70; a_mant3 = 8'd26;
b_mant0 = 8'd102; b_mant1 = 8'd113; b_mant2 = 8'd84; b_mant3 = 8'd142;
a_exp0 = 10'd481; a_exp1 = 10'd964; a_exp2 = 10'd501; a_exp3 = 10'd338;
b_exp0 = 10'd455; b_exp1 = 10'd97; b_exp2 = 10'd258; b_exp3 = 10'd112;
a_sign0 = 4'd5; a_sign1 = 4'd1; a_sign2 = 4'd15; a_sign3 = 4'd5;
b_sign0 = 4'd0; b_sign1 = 4'd5; b_sign2 = 4'd5; b_sign3 = 4'd1;
@(posedge clk_i);
shared_exps0 = 8'd134;
shared_exps1 = 8'd118;
a_mant0 = 8'd79; a_mant1 = 8'd228; a_mant2 = 8'd236; a_mant3 = 8'd228;
b_mant0 = 8'd252; b_mant1 = 8'd106; b_mant2 = 8'd172; b_mant3 = 8'd144;
a_exp0 = 10'd282; a_exp1 = 10'd468; a_exp2 = 10'd828; a_exp3 = 10'd631;
b_exp0 = 10'd211; b_exp1 = 10'd769; b_exp2 = 10'd885; b_exp3 = 10'd881;
a_sign0 = 4'd7; a_sign1 = 4'd5; a_sign2 = 4'd0; a_sign3 = 4'd2;
b_sign0 = 4'd6; b_sign1 = 4'd16; b_sign2 = 4'd8; b_sign3 = 4'd6;
@(posedge clk_i);
a_mant0 = 8'd241; a_mant1 = 8'd200; a_mant2 = 8'd243; a_mant3 = 8'd178;
b_mant0 = 8'd138; b_mant1 = 8'd91; b_mant2 = 8'd40; b_mant3 = 8'd215;
a_exp0 = 10'd646; a_exp1 = 10'd143; a_exp2 = 10'd794; a_exp3 = 10'd950;
b_exp0 = 10'd162; b_exp1 = 10'd38; b_exp2 = 10'd236; b_exp3 = 10'd287;
a_sign0 = 4'd4; a_sign1 = 4'd8; a_sign2 = 4'd8; a_sign3 = 4'd15;
b_sign0 = 4'd9; b_sign1 = 4'd13; b_sign2 = 4'd14; b_sign3 = 4'd10;
@(posedge clk_i);
a_mant0 = 8'd171; a_mant1 = 8'd240; a_mant2 = 8'd180; a_mant3 = 8'd155;
b_mant0 = 8'd54; b_mant1 = 8'd32; b_mant2 = 8'd234; b_mant3 = 8'd123;
a_exp0 = 10'd627; a_exp1 = 10'd52; a_exp2 = 10'd130; a_exp3 = 10'd688;
b_exp0 = 10'd37; b_exp1 = 10'd904; b_exp2 = 10'd699; b_exp3 = 10'd968;
a_sign0 = 4'd4; a_sign1 = 4'd10; a_sign2 = 4'd11; a_sign3 = 4'd8;
b_sign0 = 4'd10; b_sign1 = 4'd15; b_sign2 = 4'd5; b_sign3 = 4'd13;
@(posedge clk_i);
a_mant0 = 8'd145; a_mant1 = 8'd147; a_mant2 = 8'd64; a_mant3 = 8'd52;
b_mant0 = 8'd235; b_mant1 = 8'd24; b_mant2 = 8'd173; b_mant3 = 8'd126;
a_exp0 = 10'd693; a_exp1 = 10'd523; a_exp2 = 10'd206; a_exp3 = 10'd773;
b_exp0 = 10'd423; b_exp1 = 10'd936; b_exp2 = 10'd504; b_exp3 = 10'd854;
a_sign0 = 4'd10; a_sign1 = 4'd14; a_sign2 = 4'd9; a_sign3 = 4'd9;
b_sign0 = 4'd7; b_sign1 = 4'd15; b_sign2 = 4'd7; b_sign3 = 4'd16;
@(posedge clk_i);
a_mant0 = 8'd240; a_mant1 = 8'd198; a_mant2 = 8'd180; a_mant3 = 8'd58;
b_mant0 = 8'd135; b_mant1 = 8'd196; b_mant2 = 8'd36; b_mant3 = 8'd1;
a_exp0 = 10'd212; a_exp1 = 10'd728; a_exp2 = 10'd309; a_exp3 = 10'd69;
b_exp0 = 10'd74; b_exp1 = 10'd800; b_exp2 = 10'd346; b_exp3 = 10'd297;
a_sign0 = 4'd14; a_sign1 = 4'd0; a_sign2 = 4'd0; a_sign3 = 4'd11;
b_sign0 = 4'd13; b_sign1 = 4'd4; b_sign2 = 4'd7; b_sign3 = 4'd1;
@(posedge clk_i);
a_mant0 = 8'd150; a_mant1 = 8'd13; a_mant2 = 8'd135; a_mant3 = 8'd134;
b_mant0 = 8'd26; b_mant1 = 8'd148; b_mant2 = 8'd42; b_mant3 = 8'd167;
a_exp0 = 10'd233; a_exp1 = 10'd668; a_exp2 = 10'd623; a_exp3 = 10'd802;
b_exp0 = 10'd76; b_exp1 = 10'd135; b_exp2 = 10'd273; b_exp3 = 10'd743;
a_sign0 = 4'd13; a_sign1 = 4'd1; a_sign2 = 4'd14; a_sign3 = 4'd15;
b_sign0 = 4'd0; b_sign1 = 4'd7; b_sign2 = 4'd12; b_sign3 = 4'd6;
@(posedge clk_i);
a_mant0 = 8'd121; a_mant1 = 8'd177; a_mant2 = 8'd79; a_mant3 = 8'd124;
b_mant0 = 8'd121; b_mant1 = 8'd151; b_mant2 = 8'd150; b_mant3 = 8'd47;
a_exp0 = 10'd715; a_exp1 = 10'd124; a_exp2 = 10'd453; a_exp3 = 10'd988;
b_exp0 = 10'd904; b_exp1 = 10'd940; b_exp2 = 10'd456; b_exp3 = 10'd518;
a_sign0 = 4'd2; a_sign1 = 4'd9; a_sign2 = 4'd10; a_sign3 = 4'd11;
b_sign0 = 4'd0; b_sign1 = 4'd0; b_sign2 = 4'd16; b_sign3 = 4'd8;
@(posedge clk_i);
a_mant0 = 8'd137; a_mant1 = 8'd89; a_mant2 = 8'd88; a_mant3 = 8'd141;
b_mant0 = 8'd5; b_mant1 = 8'd180; b_mant2 = 8'd63; b_mant3 = 8'd163;
a_exp0 = 10'd502; a_exp1 = 10'd165; a_exp2 = 10'd629; a_exp3 = 10'd290;
b_exp0 = 10'd449; b_exp1 = 10'd341; b_exp2 = 10'd5; b_exp3 = 10'd83;
a_sign0 = 4'd6; a_sign1 = 4'd7; a_sign2 = 4'd0; a_sign3 = 4'd11;
b_sign0 = 4'd7; b_sign1 = 4'd15; b_sign2 = 4'd13; b_sign3 = 4'd13;
@(posedge clk_i);
shared_exps0 = 8'd112;
shared_exps1 = 8'd130;
rstn = 0;
@(posedge clk_i);
rstn = 1;
a_mant0 = 8'd61; a_mant1 = 8'd14; a_mant2 = 8'd49; a_mant3 = 8'd116;
b_mant0 = 8'd112; b_mant1 = 8'd67; b_mant2 = 8'd240; b_mant3 = 8'd75;
a_exp0 = 10'd74; a_exp1 = 10'd287; a_exp2 = 10'd305; a_exp3 = 10'd972;
b_exp0 = 10'd367; b_exp1 = 10'd886; b_exp2 = 10'd115; b_exp3 = 10'd771;
a_sign0 = 4'd10; a_sign1 = 4'd11; a_sign2 = 4'd15; a_sign3 = 4'd16;
b_sign0 = 4'd15; b_sign1 = 4'd4; b_sign2 = 4'd14; b_sign3 = 4'd0;
@(posedge clk_i);
a_mant0 = 8'd71; a_mant1 = 8'd120; a_mant2 = 8'd119; a_mant3 = 8'd226;
b_mant0 = 8'd85; b_mant1 = 8'd194; b_mant2 = 8'd202; b_mant3 = 8'd83;
a_exp0 = 10'd662; a_exp1 = 10'd103; a_exp2 = 10'd232; a_exp3 = 10'd30;
b_exp0 = 10'd764; b_exp1 = 10'd359; b_exp2 = 10'd718; b_exp3 = 10'd183;
a_sign0 = 4'd0; a_sign1 = 4'd12; a_sign2 = 4'd16; a_sign3 = 4'd12;
b_sign0 = 4'd16; b_sign1 = 4'd4; b_sign2 = 4'd12; b_sign3 = 4'd11;
@(posedge clk_i);
a_mant0 = 8'd67; a_mant1 = 8'd100; a_mant2 = 8'd160; a_mant3 = 8'd243;
b_mant0 = 8'd226; b_mant1 = 8'd120; b_mant2 = 8'd180; b_mant3 = 8'd121;
a_exp0 = 10'd499; a_exp1 = 10'd879; a_exp2 = 10'd949; a_exp3 = 10'd32;
b_exp0 = 10'd493; b_exp1 = 10'd733; b_exp2 = 10'd748; b_exp3 = 10'd999;
a_sign0 = 4'd5; a_sign1 = 4'd15; a_sign2 = 4'd4; a_sign3 = 4'd4;
b_sign0 = 4'd8; b_sign1 = 4'd9; b_sign2 = 4'd11; b_sign3 = 4'd5;
@(posedge clk_i);
a_mant0 = 8'd241; a_mant1 = 8'd164; a_mant2 = 8'd25; a_mant3 = 8'd113;
b_mant0 = 8'd133; b_mant1 = 8'd8; b_mant2 = 8'd72; b_mant3 = 8'd188;
a_exp0 = 10'd319; a_exp1 = 10'd2; a_exp2 = 10'd867; a_exp3 = 10'd318;
b_exp0 = 10'd423; b_exp1 = 10'd708; b_exp2 = 10'd664; b_exp3 = 10'd615;
a_sign0 = 4'd2; a_sign1 = 4'd0; a_sign2 = 4'd2; a_sign3 = 4'd14;
b_sign0 = 4'd4; b_sign1 = 4'd10; b_sign2 = 4'd14; b_sign3 = 4'd6;
@(posedge clk_i);
a_mant0 = 8'd119; a_mant1 = 8'd18; a_mant2 = 8'd197; a_mant3 = 8'd217;
b_mant0 = 8'd3; b_mant1 = 8'd206; b_mant2 = 8'd130; b_mant3 = 8'd49;
a_exp0 = 10'd229; a_exp1 = 10'd357; a_exp2 = 10'd280; a_exp3 = 10'd817;
b_exp0 = 10'd822; b_exp1 = 10'd343; b_exp2 = 10'd789; b_exp3 = 10'd896;
a_sign0 = 4'd11; a_sign1 = 4'd13; a_sign2 = 4'd2; a_sign3 = 4'd14;
b_sign0 = 4'd10; b_sign1 = 4'd5; b_sign2 = 4'd0; b_sign3 = 4'd12;
@(posedge clk_i);
a_mant0 = 8'd11; a_mant1 = 8'd190; a_mant2 = 8'd143; a_mant3 = 8'd12;
b_mant0 = 8'd204; b_mant1 = 8'd148; b_mant2 = 8'd179; b_mant3 = 8'd141;
a_exp0 = 10'd151; a_exp1 = 10'd443; a_exp2 = 10'd303; a_exp3 = 10'd495;
b_exp0 = 10'd193; b_exp1 = 10'd879; b_exp2 = 10'd802; b_exp3 = 10'd909;
a_sign0 = 4'd0; a_sign1 = 4'd8; a_sign2 = 4'd15; a_sign3 = 4'd4;
b_sign0 = 4'd11; b_sign1 = 4'd2; b_sign2 = 4'd3; b_sign3 = 4'd3;
@(posedge clk_i);
a_mant0 = 8'd217; a_mant1 = 8'd195; a_mant2 = 8'd101; a_mant3 = 8'd31;
b_mant0 = 8'd188; b_mant1 = 8'd87; b_mant2 = 8'd170; b_mant3 = 8'd63;
a_exp0 = 10'd224; a_exp1 = 10'd311; a_exp2 = 10'd211; a_exp3 = 10'd938;
b_exp0 = 10'd320; b_exp1 = 10'd232; b_exp2 = 10'd500; b_exp3 = 10'd120;
a_sign0 = 4'd16; a_sign1 = 4'd11; a_sign2 = 4'd5; a_sign3 = 4'd7;
b_sign0 = 4'd13; b_sign1 = 4'd4; b_sign2 = 4'd12; b_sign3 = 4'd11;
@(posedge clk_i);
shared_exps0 = 8'd109;
shared_exps1 = 8'd149;
a_mant0 = 8'd13; a_mant1 = 8'd110; a_mant2 = 8'd145; a_mant3 = 8'd202;
b_mant0 = 8'd205; b_mant1 = 8'd255; b_mant2 = 8'd56; b_mant3 = 8'd246;
a_exp0 = 10'd494; a_exp1 = 10'd557; a_exp2 = 10'd251; a_exp3 = 10'd845;
b_exp0 = 10'd143; b_exp1 = 10'd282; b_exp2 = 10'd896; b_exp3 = 10'd313;
a_sign0 = 4'd15; a_sign1 = 4'd6; a_sign2 = 4'd5; a_sign3 = 4'd7;
b_sign0 = 4'd11; b_sign1 = 4'd3; b_sign2 = 4'd5; b_sign3 = 4'd11;
@(posedge clk_i);
a_mant0 = 8'd134; a_mant1 = 8'd231; a_mant2 = 8'd91; a_mant3 = 8'd55;
b_mant0 = 8'd27; b_mant1 = 8'd255; b_mant2 = 8'd48; b_mant3 = 8'd36;
a_exp0 = 10'd1012; a_exp1 = 10'd690; a_exp2 = 10'd619; a_exp3 = 10'd227;
b_exp0 = 10'd874; b_exp1 = 10'd290; b_exp2 = 10'd867; b_exp3 = 10'd508;
a_sign0 = 4'd13; a_sign1 = 4'd3; a_sign2 = 4'd2; a_sign3 = 4'd10;
b_sign0 = 4'd9; b_sign1 = 4'd4; b_sign2 = 4'd4; b_sign3 = 4'd11;
@(posedge clk_i);
a_mant0 = 8'd104; a_mant1 = 8'd132; a_mant2 = 8'd103; a_mant3 = 8'd231;
b_mant0 = 8'd201; b_mant1 = 8'd93; b_mant2 = 8'd172; b_mant3 = 8'd69;
a_exp0 = 10'd497; a_exp1 = 10'd213; a_exp2 = 10'd998; a_exp3 = 10'd94;
b_exp0 = 10'd650; b_exp1 = 10'd1002; b_exp2 = 10'd530; b_exp3 = 10'd335;
a_sign0 = 4'd13; a_sign1 = 4'd1; a_sign2 = 4'd7; a_sign3 = 4'd8;
b_sign0 = 4'd0; b_sign1 = 4'd13; b_sign2 = 4'd9; b_sign3 = 4'd10;
@(posedge clk_i);
a_mant0 = 8'd204; a_mant1 = 8'd223; a_mant2 = 8'd250; a_mant3 = 8'd56;
b_mant0 = 8'd144; b_mant1 = 8'd95; b_mant2 = 8'd198; b_mant3 = 8'd235;
a_exp0 = 10'd311; a_exp1 = 10'd905; a_exp2 = 10'd285; a_exp3 = 10'd434;
b_exp0 = 10'd63; b_exp1 = 10'd736; b_exp2 = 10'd864; b_exp3 = 10'd370;
a_sign0 = 4'd6; a_sign1 = 4'd16; a_sign2 = 4'd7; a_sign3 = 4'd13;
b_sign0 = 4'd13; b_sign1 = 4'd0; b_sign2 = 4'd1; b_sign3 = 4'd10;
@(posedge clk_i);
a_mant0 = 8'd248; a_mant1 = 8'd136; a_mant2 = 8'd11; a_mant3 = 8'd65;
b_mant0 = 8'd119; b_mant1 = 8'd43; b_mant2 = 8'd155; b_mant3 = 8'd164;
a_exp0 = 10'd365; a_exp1 = 10'd926; a_exp2 = 10'd155; a_exp3 = 10'd88;
b_exp0 = 10'd835; b_exp1 = 10'd528; b_exp2 = 10'd687; b_exp3 = 10'd917;
a_sign0 = 4'd11; a_sign1 = 4'd7; a_sign2 = 4'd7; a_sign3 = 4'd16;
b_sign0 = 4'd10; b_sign1 = 4'd3; b_sign2 = 4'd10; b_sign3 = 4'd13;
@(posedge clk_i);
a_mant0 = 8'd220; a_mant1 = 8'd107; a_mant2 = 8'd169; a_mant3 = 8'd168;
b_mant0 = 8'd17; b_mant1 = 8'd78; b_mant2 = 8'd134; b_mant3 = 8'd125;
a_exp0 = 10'd102; a_exp1 = 10'd304; a_exp2 = 10'd608; a_exp3 = 10'd558;
b_exp0 = 10'd837; b_exp1 = 10'd740; b_exp2 = 10'd584; b_exp3 = 10'd938;
a_sign0 = 4'd6; a_sign1 = 4'd7; a_sign2 = 4'd6; a_sign3 = 4'd13;
b_sign0 = 4'd8; b_sign1 = 4'd5; b_sign2 = 4'd15; b_sign3 = 4'd5;
@(posedge clk_i);
a_mant0 = 8'd206; a_mant1 = 8'd106; a_mant2 = 8'd237; a_mant3 = 8'd219;
b_mant0 = 8'd62; b_mant1 = 8'd83; b_mant2 = 8'd49; b_mant3 = 8'd80;
a_exp0 = 10'd61; a_exp1 = 10'd426; a_exp2 = 10'd931; a_exp3 = 10'd277;
b_exp0 = 10'd567; b_exp1 = 10'd140; b_exp2 = 10'd837; b_exp3 = 10'd971;
a_sign0 = 4'd3; a_sign1 = 4'd3; a_sign2 = 4'd0; a_sign3 = 4'd10;
b_sign0 = 4'd8; b_sign1 = 4'd0; b_sign2 = 4'd8; b_sign3 = 4'd9;
@(posedge clk_i);
a_mant0 = 8'd186; a_mant1 = 8'd133; a_mant2 = 8'd61; a_mant3 = 8'd171;
b_mant0 = 8'd139; b_mant1 = 8'd69; b_mant2 = 8'd142; b_mant3 = 8'd203;
a_exp0 = 10'd395; a_exp1 = 10'd112; a_exp2 = 10'd465; a_exp3 = 10'd868;
b_exp0 = 10'd336; b_exp1 = 10'd182; b_exp2 = 10'd410; b_exp3 = 10'd220;
a_sign0 = 4'd7; a_sign1 = 4'd11; a_sign2 = 4'd13; a_sign3 = 4'd8;
b_sign0 = 4'd3; b_sign1 = 4'd8; b_sign2 = 4'd9; b_sign3 = 4'd16;
@(posedge clk_i);
shared_exps0 = 8'd122;
shared_exps1 = 8'd151;
a_mant0 = 8'd241; a_mant1 = 8'd138; a_mant2 = 8'd241; a_mant3 = 8'd106;
b_mant0 = 8'd248; b_mant1 = 8'd227; b_mant2 = 8'd67; b_mant3 = 8'd147;
a_exp0 = 10'd96; a_exp1 = 10'd139; a_exp2 = 10'd604; a_exp3 = 10'd529;
b_exp0 = 10'd301; b_exp1 = 10'd841; b_exp2 = 10'd136; b_exp3 = 10'd410;
a_sign0 = 4'd13; a_sign1 = 4'd6; a_sign2 = 4'd2; a_sign3 = 4'd4;
b_sign0 = 4'd3; b_sign1 = 4'd3; b_sign2 = 4'd14; b_sign3 = 4'd5;
@(posedge clk_i);
a_mant0 = 8'd10; a_mant1 = 8'd191; a_mant2 = 8'd82; a_mant3 = 8'd231;
b_mant0 = 8'd114; b_mant1 = 8'd165; b_mant2 = 8'd30; b_mant3 = 8'd23;
a_exp0 = 10'd384; a_exp1 = 10'd753; a_exp2 = 10'd749; a_exp3 = 10'd338;
b_exp0 = 10'd636; b_exp1 = 10'd728; b_exp2 = 10'd305; b_exp3 = 10'd232;
a_sign0 = 4'd5; a_sign1 = 4'd14; a_sign2 = 4'd11; a_sign3 = 4'd6;
b_sign0 = 4'd12; b_sign1 = 4'd11; b_sign2 = 4'd1; b_sign3 = 4'd11;
@(posedge clk_i);
a_mant0 = 8'd253; a_mant1 = 8'd207; a_mant2 = 8'd87; a_mant3 = 8'd248;
b_mant0 = 8'd17; b_mant1 = 8'd255; b_mant2 = 8'd239; b_mant3 = 8'd121;
a_exp0 = 10'd430; a_exp1 = 10'd511; a_exp2 = 10'd308; a_exp3 = 10'd786;
b_exp0 = 10'd236; b_exp1 = 10'd952; b_exp2 = 10'd888; b_exp3 = 10'd884;
a_sign0 = 4'd1; a_sign1 = 4'd5; a_sign2 = 4'd0; a_sign3 = 4'd7;
b_sign0 = 4'd3; b_sign1 = 4'd5; b_sign2 = 4'd16; b_sign3 = 4'd3;
@(posedge clk_i);
a_mant0 = 8'd93; a_mant1 = 8'd158; a_mant2 = 8'd134; a_mant3 = 8'd249;
b_mant0 = 8'd102; b_mant1 = 8'd169; b_mant2 = 8'd77; b_mant3 = 8'd157;
a_exp0 = 10'd660; a_exp1 = 10'd101; a_exp2 = 10'd129; a_exp3 = 10'd148;
b_exp0 = 10'd607; b_exp1 = 10'd160; b_exp2 = 10'd74; b_exp3 = 10'd62;
a_sign0 = 4'd8; a_sign1 = 4'd3; a_sign2 = 4'd1; a_sign3 = 4'd3;
b_sign0 = 4'd14; b_sign1 = 4'd3; b_sign2 = 4'd1; b_sign3 = 4'd13;
@(posedge clk_i);
a_mant0 = 8'd94; a_mant1 = 8'd145; a_mant2 = 8'd189; a_mant3 = 8'd135;
b_mant0 = 8'd243; b_mant1 = 8'd199; b_mant2 = 8'd35; b_mant3 = 8'd186;
a_exp0 = 10'd325; a_exp1 = 10'd482; a_exp2 = 10'd508; a_exp3 = 10'd498;
b_exp0 = 10'd326; b_exp1 = 10'd733; b_exp2 = 10'd646; b_exp3 = 10'd177;
a_sign0 = 4'd9; a_sign1 = 4'd2; a_sign2 = 4'd14; a_sign3 = 4'd9;
b_sign0 = 4'd2; b_sign1 = 4'd14; b_sign2 = 4'd5; b_sign3 = 4'd5;
@(posedge clk_i);
a_mant0 = 8'd102; a_mant1 = 8'd211; a_mant2 = 8'd223; a_mant3 = 8'd76;
b_mant0 = 8'd15; b_mant1 = 8'd125; b_mant2 = 8'd207; b_mant3 = 8'd110;
a_exp0 = 10'd608; a_exp1 = 10'd602; a_exp2 = 10'd103; a_exp3 = 10'd878;
b_exp0 = 10'd32; b_exp1 = 10'd698; b_exp2 = 10'd468; b_exp3 = 10'd1021;
a_sign0 = 4'd5; a_sign1 = 4'd14; a_sign2 = 4'd8; a_sign3 = 4'd16;
b_sign0 = 4'd1; b_sign1 = 4'd16; b_sign2 = 4'd4; b_sign3 = 4'd16;
@(posedge clk_i);
a_mant0 = 8'd59; a_mant1 = 8'd66; a_mant2 = 8'd186; a_mant3 = 8'd221;
b_mant0 = 8'd42; b_mant1 = 8'd204; b_mant2 = 8'd76; b_mant3 = 8'd171;
a_exp0 = 10'd995; a_exp1 = 10'd149; a_exp2 = 10'd963; a_exp3 = 10'd837;
b_exp0 = 10'd2; b_exp1 = 10'd175; b_exp2 = 10'd176; b_exp3 = 10'd662;
a_sign0 = 4'd1; a_sign1 = 4'd5; a_sign2 = 4'd5; a_sign3 = 4'd3;
b_sign0 = 4'd9; b_sign1 = 4'd13; b_sign2 = 4'd13; b_sign3 = 4'd4;
@(posedge clk_i);
a_mant0 = 8'd170; a_mant1 = 8'd135; a_mant2 = 8'd203; a_mant3 = 8'd117;
b_mant0 = 8'd2; b_mant1 = 8'd200; b_mant2 = 8'd25; b_mant3 = 8'd105;
a_exp0 = 10'd761; a_exp1 = 10'd378; a_exp2 = 10'd456; a_exp3 = 10'd490;
b_exp0 = 10'd515; b_exp1 = 10'd975; b_exp2 = 10'd782; b_exp3 = 10'd184;
a_sign0 = 4'd3; a_sign1 = 4'd2; a_sign2 = 4'd15; a_sign3 = 4'd3;
b_sign0 = 4'd2; b_sign1 = 4'd15; b_sign2 = 4'd2; b_sign3 = 4'd6;
@(posedge clk_i);
shared_exps0 = 8'd113;
shared_exps1 = 8'd111;
a_mant0 = 8'd113; a_mant1 = 8'd209; a_mant2 = 8'd143; a_mant3 = 8'd67;
b_mant0 = 8'd202; b_mant1 = 8'd188; b_mant2 = 8'd24; b_mant3 = 8'd235;
a_exp0 = 10'd959; a_exp1 = 10'd770; a_exp2 = 10'd935; a_exp3 = 10'd216;
b_exp0 = 10'd359; b_exp1 = 10'd266; b_exp2 = 10'd56; b_exp3 = 10'd167;
a_sign0 = 4'd11; a_sign1 = 4'd11; a_sign2 = 4'd6; a_sign3 = 4'd15;
b_sign0 = 4'd15; b_sign1 = 4'd11; b_sign2 = 4'd10; b_sign3 = 4'd10;
@(posedge clk_i);
a_mant0 = 8'd247; a_mant1 = 8'd252; a_mant2 = 8'd120; a_mant3 = 8'd170;
b_mant0 = 8'd204; b_mant1 = 8'd145; b_mant2 = 8'd199; b_mant3 = 8'd73;
a_exp0 = 10'd603; a_exp1 = 10'd381; a_exp2 = 10'd945; a_exp3 = 10'd931;
b_exp0 = 10'd1; b_exp1 = 10'd884; b_exp2 = 10'd176; b_exp3 = 10'd651;
a_sign0 = 4'd15; a_sign1 = 4'd9; a_sign2 = 4'd2; a_sign3 = 4'd13;
b_sign0 = 4'd11; b_sign1 = 4'd12; b_sign2 = 4'd8; b_sign3 = 4'd15;
@(posedge clk_i);
a_mant0 = 8'd205; a_mant1 = 8'd221; a_mant2 = 8'd218; a_mant3 = 8'd120;
b_mant0 = 8'd177; b_mant1 = 8'd74; b_mant2 = 8'd239; b_mant3 = 8'd108;
a_exp0 = 10'd150; a_exp1 = 10'd457; a_exp2 = 10'd492; a_exp3 = 10'd688;
b_exp0 = 10'd461; b_exp1 = 10'd264; b_exp2 = 10'd292; b_exp3 = 10'd69;
a_sign0 = 4'd8; a_sign1 = 4'd5; a_sign2 = 4'd0; a_sign3 = 4'd2;
b_sign0 = 4'd7; b_sign1 = 4'd8; b_sign2 = 4'd11; b_sign3 = 4'd14;
@(posedge clk_i);
a_mant0 = 8'd150; a_mant1 = 8'd33; a_mant2 = 8'd228; a_mant3 = 8'd59;
b_mant0 = 8'd253; b_mant1 = 8'd174; b_mant2 = 8'd66; b_mant3 = 8'd166;
a_exp0 = 10'd603; a_exp1 = 10'd422; a_exp2 = 10'd648; a_exp3 = 10'd455;
b_exp0 = 10'd96; b_exp1 = 10'd371; b_exp2 = 10'd828; b_exp3 = 10'd522;
a_sign0 = 4'd8; a_sign1 = 4'd15; a_sign2 = 4'd11; a_sign3 = 4'd9;
b_sign0 = 4'd1; b_sign1 = 4'd3; b_sign2 = 4'd9; b_sign3 = 4'd14;
@(posedge clk_i);
a_mant0 = 8'd255; a_mant1 = 8'd164; a_mant2 = 8'd7; a_mant3 = 8'd229;
b_mant0 = 8'd50; b_mant1 = 8'd182; b_mant2 = 8'd41; b_mant3 = 8'd66;
a_exp0 = 10'd339; a_exp1 = 10'd352; a_exp2 = 10'd26; a_exp3 = 10'd692;
b_exp0 = 10'd69; b_exp1 = 10'd756; b_exp2 = 10'd1017; b_exp3 = 10'd861;
a_sign0 = 4'd12; a_sign1 = 4'd13; a_sign2 = 4'd10; a_sign3 = 4'd11;
b_sign0 = 4'd15; b_sign1 = 4'd3; b_sign2 = 4'd4; b_sign3 = 4'd13;
@(posedge clk_i);
a_mant0 = 8'd194; a_mant1 = 8'd223; a_mant2 = 8'd70; a_mant3 = 8'd65;
b_mant0 = 8'd178; b_mant1 = 8'd129; b_mant2 = 8'd148; b_mant3 = 8'd211;
a_exp0 = 10'd368; a_exp1 = 10'd420; a_exp2 = 10'd672; a_exp3 = 10'd618;
b_exp0 = 10'd408; b_exp1 = 10'd324; b_exp2 = 10'd295; b_exp3 = 10'd895;
a_sign0 = 4'd16; a_sign1 = 4'd6; a_sign2 = 4'd6; a_sign3 = 4'd14;
b_sign0 = 4'd1; b_sign1 = 4'd16; b_sign2 = 4'd7; b_sign3 = 4'd15;
@(posedge clk_i);
a_mant0 = 8'd243; a_mant1 = 8'd105; a_mant2 = 8'd71; a_mant3 = 8'd204;
b_mant0 = 8'd184; b_mant1 = 8'd152; b_mant2 = 8'd226; b_mant3 = 8'd225;
a_exp0 = 10'd211; a_exp1 = 10'd474; a_exp2 = 10'd213; a_exp3 = 10'd567;
b_exp0 = 10'd50; b_exp1 = 10'd692; b_exp2 = 10'd229; b_exp3 = 10'd550;
a_sign0 = 4'd0; a_sign1 = 4'd13; a_sign2 = 4'd6; a_sign3 = 4'd9;
b_sign0 = 4'd10; b_sign1 = 4'd8; b_sign2 = 4'd14; b_sign3 = 4'd6;
@(posedge clk_i);
a_mant0 = 8'd210; a_mant1 = 8'd137; a_mant2 = 8'd90; a_mant3 = 8'd221;
b_mant0 = 8'd18; b_mant1 = 8'd176; b_mant2 = 8'd188; b_mant3 = 8'd7;
a_exp0 = 10'd425; a_exp1 = 10'd568; a_exp2 = 10'd794; a_exp3 = 10'd608;
b_exp0 = 10'd103; b_exp1 = 10'd499; b_exp2 = 10'd584; b_exp3 = 10'd192;
a_sign0 = 4'd6; a_sign1 = 4'd11; a_sign2 = 4'd5; a_sign3 = 4'd15;
b_sign0 = 4'd13; b_sign1 = 4'd8; b_sign2 = 4'd5; b_sign3 = 4'd9;
@(posedge clk_i);
shared_exps0 = 8'd108;
shared_exps1 = 8'd109;
rstn = 0;
@(posedge clk_i);
rstn = 1;
a_mant0 = 8'd152; a_mant1 = 8'd214; a_mant2 = 8'd195; a_mant3 = 8'd50;
b_mant0 = 8'd152; b_mant1 = 8'd62; b_mant2 = 8'd191; b_mant3 = 8'd180;
a_exp0 = 10'd212; a_exp1 = 10'd164; a_exp2 = 10'd467; a_exp3 = 10'd152;
b_exp0 = 10'd973; b_exp1 = 10'd90; b_exp2 = 10'd899; b_exp3 = 10'd398;
a_sign0 = 4'd16; a_sign1 = 4'd10; a_sign2 = 4'd3; a_sign3 = 4'd16;
b_sign0 = 4'd8; b_sign1 = 4'd8; b_sign2 = 4'd12; b_sign3 = 4'd11;
@(posedge clk_i);
a_mant0 = 8'd205; a_mant1 = 8'd155; a_mant2 = 8'd220; a_mant3 = 8'd14;
b_mant0 = 8'd185; b_mant1 = 8'd149; b_mant2 = 8'd110; b_mant3 = 8'd47;
a_exp0 = 10'd669; a_exp1 = 10'd929; a_exp2 = 10'd263; a_exp3 = 10'd418;
b_exp0 = 10'd1; b_exp1 = 10'd132; b_exp2 = 10'd107; b_exp3 = 10'd165;
a_sign0 = 4'd8; a_sign1 = 4'd3; a_sign2 = 4'd12; a_sign3 = 4'd11;
b_sign0 = 4'd10; b_sign1 = 4'd16; b_sign2 = 4'd0; b_sign3 = 4'd7;
@(posedge clk_i);
a_mant0 = 8'd164; a_mant1 = 8'd142; a_mant2 = 8'd166; a_mant3 = 8'd89;
b_mant0 = 8'd197; b_mant1 = 8'd120; b_mant2 = 8'd8; b_mant3 = 8'd233;
a_exp0 = 10'd607; a_exp1 = 10'd654; a_exp2 = 10'd134; a_exp3 = 10'd850;
b_exp0 = 10'd180; b_exp1 = 10'd160; b_exp2 = 10'd628; b_exp3 = 10'd9;
a_sign0 = 4'd2; a_sign1 = 4'd4; a_sign2 = 4'd6; a_sign3 = 4'd12;
b_sign0 = 4'd0; b_sign1 = 4'd15; b_sign2 = 4'd15; b_sign3 = 4'd16;
@(posedge clk_i);
a_mant0 = 8'd62; a_mant1 = 8'd101; a_mant2 = 8'd164; a_mant3 = 8'd173;
b_mant0 = 8'd169; b_mant1 = 8'd78; b_mant2 = 8'd244; b_mant3 = 8'd126;
a_exp0 = 10'd107; a_exp1 = 10'd1006; a_exp2 = 10'd327; a_exp3 = 10'd549;
b_exp0 = 10'd317; b_exp1 = 10'd419; b_exp2 = 10'd566; b_exp3 = 10'd984;
a_sign0 = 4'd5; a_sign1 = 4'd15; a_sign2 = 4'd3; a_sign3 = 4'd10;
b_sign0 = 4'd13; b_sign1 = 4'd11; b_sign2 = 4'd16; b_sign3 = 4'd13;
@(posedge clk_i);
a_mant0 = 8'd185; a_mant1 = 8'd53; a_mant2 = 8'd247; a_mant3 = 8'd22;
b_mant0 = 8'd77; b_mant1 = 8'd242; b_mant2 = 8'd196; b_mant3 = 8'd106;
a_exp0 = 10'd895; a_exp1 = 10'd503; a_exp2 = 10'd740; a_exp3 = 10'd450;
b_exp0 = 10'd205; b_exp1 = 10'd222; b_exp2 = 10'd834; b_exp3 = 10'd552;
a_sign0 = 4'd15; a_sign1 = 4'd13; a_sign2 = 4'd5; a_sign3 = 4'd16;
b_sign0 = 4'd2; b_sign1 = 4'd16; b_sign2 = 4'd2; b_sign3 = 4'd4;
@(posedge clk_i);
a_mant0 = 8'd226; a_mant1 = 8'd226; a_mant2 = 8'd51; a_mant3 = 8'd132;
b_mant0 = 8'd59; b_mant1 = 8'd37; b_mant2 = 8'd8; b_mant3 = 8'd236;
a_exp0 = 10'd67; a_exp1 = 10'd670; a_exp2 = 10'd676; a_exp3 = 10'd840;
b_exp0 = 10'd270; b_exp1 = 10'd988; b_exp2 = 10'd197; b_exp3 = 10'd303;
a_sign0 = 4'd11; a_sign1 = 4'd10; a_sign2 = 4'd11; a_sign3 = 4'd9;
b_sign0 = 4'd7; b_sign1 = 4'd11; b_sign2 = 4'd14; b_sign3 = 4'd5;
@(posedge clk_i);
a_mant0 = 8'd96; a_mant1 = 8'd176; a_mant2 = 8'd155; a_mant3 = 8'd159;
b_mant0 = 8'd177; b_mant1 = 8'd222; b_mant2 = 8'd130; b_mant3 = 8'd236;
a_exp0 = 10'd280; a_exp1 = 10'd987; a_exp2 = 10'd455; a_exp3 = 10'd229;
b_exp0 = 10'd73; b_exp1 = 10'd514; b_exp2 = 10'd348; b_exp3 = 10'd972;
a_sign0 = 4'd13; a_sign1 = 4'd12; a_sign2 = 4'd5; a_sign3 = 4'd6;
b_sign0 = 4'd10; b_sign1 = 4'd1; b_sign2 = 4'd15; b_sign3 = 4'd4;
@(posedge clk_i);
shared_exps0 = 8'd138;
shared_exps1 = 8'd143;
a_mant0 = 8'd68; a_mant1 = 8'd47; a_mant2 = 8'd76; a_mant3 = 8'd187;
b_mant0 = 8'd127; b_mant1 = 8'd254; b_mant2 = 8'd153; b_mant3 = 8'd237;
a_exp0 = 10'd333; a_exp1 = 10'd561; a_exp2 = 10'd591; a_exp3 = 10'd723;
b_exp0 = 10'd345; b_exp1 = 10'd204; b_exp2 = 10'd547; b_exp3 = 10'd803;
a_sign0 = 4'd1; a_sign1 = 4'd2; a_sign2 = 4'd4; a_sign3 = 4'd6;
b_sign0 = 4'd15; b_sign1 = 4'd7; b_sign2 = 4'd12; b_sign3 = 4'd12;
@(posedge clk_i);
a_mant0 = 8'd206; a_mant1 = 8'd12; a_mant2 = 8'd87; a_mant3 = 8'd137;
b_mant0 = 8'd67; b_mant1 = 8'd126; b_mant2 = 8'd90; b_mant3 = 8'd253;
a_exp0 = 10'd974; a_exp1 = 10'd300; a_exp2 = 10'd833; a_exp3 = 10'd803;
b_exp0 = 10'd769; b_exp1 = 10'd460; b_exp2 = 10'd781; b_exp3 = 10'd955;
a_sign0 = 4'd8; a_sign1 = 4'd11; a_sign2 = 4'd6; a_sign3 = 4'd12;
b_sign0 = 4'd2; b_sign1 = 4'd14; b_sign2 = 4'd15; b_sign3 = 4'd7;
@(posedge clk_i);
a_mant0 = 8'd219; a_mant1 = 8'd215; a_mant2 = 8'd76; a_mant3 = 8'd54;
b_mant0 = 8'd139; b_mant1 = 8'd142; b_mant2 = 8'd204; b_mant3 = 8'd131;
a_exp0 = 10'd791; a_exp1 = 10'd283; a_exp2 = 10'd212; a_exp3 = 10'd457;
b_exp0 = 10'd158; b_exp1 = 10'd232; b_exp2 = 10'd735; b_exp3 = 10'd920;
a_sign0 = 4'd2; a_sign1 = 4'd1; a_sign2 = 4'd7; a_sign3 = 4'd2;
b_sign0 = 4'd12; b_sign1 = 4'd5; b_sign2 = 4'd7; b_sign3 = 4'd3;
@(posedge clk_i);
a_mant0 = 8'd57; a_mant1 = 8'd166; a_mant2 = 8'd212; a_mant3 = 8'd41;
b_mant0 = 8'd177; b_mant1 = 8'd79; b_mant2 = 8'd246; b_mant3 = 8'd113;
a_exp0 = 10'd909; a_exp1 = 10'd291; a_exp2 = 10'd741; a_exp3 = 10'd671;
b_exp0 = 10'd841; b_exp1 = 10'd359; b_exp2 = 10'd743; b_exp3 = 10'd760;
a_sign0 = 4'd6; a_sign1 = 4'd16; a_sign2 = 4'd6; a_sign3 = 4'd5;
b_sign0 = 4'd4; b_sign1 = 4'd2; b_sign2 = 4'd0; b_sign3 = 4'd11;
@(posedge clk_i);
a_mant0 = 8'd142; a_mant1 = 8'd210; a_mant2 = 8'd145; a_mant3 = 8'd37;
b_mant0 = 8'd153; b_mant1 = 8'd215; b_mant2 = 8'd137; b_mant3 = 8'd192;
a_exp0 = 10'd409; a_exp1 = 10'd580; a_exp2 = 10'd544; a_exp3 = 10'd150;
b_exp0 = 10'd795; b_exp1 = 10'd92; b_exp2 = 10'd78; b_exp3 = 10'd824;
a_sign0 = 4'd10; a_sign1 = 4'd16; a_sign2 = 4'd14; a_sign3 = 4'd7;
b_sign0 = 4'd6; b_sign1 = 4'd7; b_sign2 = 4'd6; b_sign3 = 4'd14;
@(posedge clk_i);
a_mant0 = 8'd46; a_mant1 = 8'd106; a_mant2 = 8'd222; a_mant3 = 8'd105;
b_mant0 = 8'd1; b_mant1 = 8'd51; b_mant2 = 8'd183; b_mant3 = 8'd73;
a_exp0 = 10'd1017; a_exp1 = 10'd603; a_exp2 = 10'd126; a_exp3 = 10'd700;
b_exp0 = 10'd889; b_exp1 = 10'd362; b_exp2 = 10'd769; b_exp3 = 10'd560;
a_sign0 = 4'd2; a_sign1 = 4'd15; a_sign2 = 4'd8; a_sign3 = 4'd11;
b_sign0 = 4'd5; b_sign1 = 4'd9; b_sign2 = 4'd1; b_sign3 = 4'd7;
@(posedge clk_i);
a_mant0 = 8'd223; a_mant1 = 8'd165; a_mant2 = 8'd120; a_mant3 = 8'd255;
b_mant0 = 8'd253; b_mant1 = 8'd104; b_mant2 = 8'd204; b_mant3 = 8'd141;
a_exp0 = 10'd100; a_exp1 = 10'd510; a_exp2 = 10'd505; a_exp3 = 10'd618;
b_exp0 = 10'd514; b_exp1 = 10'd685; b_exp2 = 10'd1023; b_exp3 = 10'd565;
a_sign0 = 4'd11; a_sign1 = 4'd7; a_sign2 = 4'd4; a_sign3 = 4'd1;
b_sign0 = 4'd5; b_sign1 = 4'd12; b_sign2 = 4'd4; b_sign3 = 4'd0;
@(posedge clk_i);
a_mant0 = 8'd62; a_mant1 = 8'd200; a_mant2 = 8'd210; a_mant3 = 8'd121;
b_mant0 = 8'd13; b_mant1 = 8'd49; b_mant2 = 8'd4; b_mant3 = 8'd219;
a_exp0 = 10'd328; a_exp1 = 10'd959; a_exp2 = 10'd404; a_exp3 = 10'd566;
b_exp0 = 10'd998; b_exp1 = 10'd80; b_exp2 = 10'd731; b_exp3 = 10'd125;
a_sign0 = 4'd16; a_sign1 = 4'd1; a_sign2 = 4'd14; a_sign3 = 4'd8;
b_sign0 = 4'd14; b_sign1 = 4'd8; b_sign2 = 4'd15; b_sign3 = 4'd8;
@(posedge clk_i);
shared_exps0 = 8'd149;
shared_exps1 = 8'd135;
a_mant0 = 8'd166; a_mant1 = 8'd238; a_mant2 = 8'd116; a_mant3 = 8'd216;
b_mant0 = 8'd225; b_mant1 = 8'd119; b_mant2 = 8'd91; b_mant3 = 8'd83;
a_exp0 = 10'd685; a_exp1 = 10'd898; a_exp2 = 10'd989; a_exp3 = 10'd588;
b_exp0 = 10'd324; b_exp1 = 10'd869; b_exp2 = 10'd459; b_exp3 = 10'd351;
a_sign0 = 4'd12; a_sign1 = 4'd10; a_sign2 = 4'd3; a_sign3 = 4'd4;
b_sign0 = 4'd13; b_sign1 = 4'd15; b_sign2 = 4'd0; b_sign3 = 4'd1;
@(posedge clk_i);
a_mant0 = 8'd216; a_mant1 = 8'd162; a_mant2 = 8'd83; a_mant3 = 8'd90;
b_mant0 = 8'd39; b_mant1 = 8'd87; b_mant2 = 8'd138; b_mant3 = 8'd92;
a_exp0 = 10'd510; a_exp1 = 10'd964; a_exp2 = 10'd953; a_exp3 = 10'd703;
b_exp0 = 10'd805; b_exp1 = 10'd524; b_exp2 = 10'd1019; b_exp3 = 10'd356;
a_sign0 = 4'd5; a_sign1 = 4'd4; a_sign2 = 4'd3; a_sign3 = 4'd2;
b_sign0 = 4'd13; b_sign1 = 4'd2; b_sign2 = 4'd13; b_sign3 = 4'd2;
@(posedge clk_i);
a_mant0 = 8'd204; a_mant1 = 8'd110; a_mant2 = 8'd33; a_mant3 = 8'd83;
b_mant0 = 8'd196; b_mant1 = 8'd95; b_mant2 = 8'd191; b_mant3 = 8'd184;
a_exp0 = 10'd757; a_exp1 = 10'd789; a_exp2 = 10'd74; a_exp3 = 10'd587;
b_exp0 = 10'd632; b_exp1 = 10'd289; b_exp2 = 10'd1006; b_exp3 = 10'd757;
a_sign0 = 4'd8; a_sign1 = 4'd2; a_sign2 = 4'd12; a_sign3 = 4'd7;
b_sign0 = 4'd15; b_sign1 = 4'd1; b_sign2 = 4'd5; b_sign3 = 4'd14;
@(posedge clk_i);
a_mant0 = 8'd78; a_mant1 = 8'd219; a_mant2 = 8'd175; a_mant3 = 8'd255;
b_mant0 = 8'd93; b_mant1 = 8'd149; b_mant2 = 8'd185; b_mant3 = 8'd42;
a_exp0 = 10'd746; a_exp1 = 10'd307; a_exp2 = 10'd193; a_exp3 = 10'd662;
b_exp0 = 10'd116; b_exp1 = 10'd645; b_exp2 = 10'd347; b_exp3 = 10'd697;
a_sign0 = 4'd14; a_sign1 = 4'd15; a_sign2 = 4'd14; a_sign3 = 4'd13;
b_sign0 = 4'd3; b_sign1 = 4'd4; b_sign2 = 4'd8; b_sign3 = 4'd11;
@(posedge clk_i);
a_mant0 = 8'd220; a_mant1 = 8'd164; a_mant2 = 8'd114; a_mant3 = 8'd239;
b_mant0 = 8'd222; b_mant1 = 8'd18; b_mant2 = 8'd104; b_mant3 = 8'd203;
a_exp0 = 10'd50; a_exp1 = 10'd783; a_exp2 = 10'd323; a_exp3 = 10'd882;
b_exp0 = 10'd112; b_exp1 = 10'd298; b_exp2 = 10'd686; b_exp3 = 10'd440;
a_sign0 = 4'd5; a_sign1 = 4'd12; a_sign2 = 4'd11; a_sign3 = 4'd16;
b_sign0 = 4'd5; b_sign1 = 4'd13; b_sign2 = 4'd1; b_sign3 = 4'd14;
@(posedge clk_i);
a_mant0 = 8'd119; a_mant1 = 8'd64; a_mant2 = 8'd88; a_mant3 = 8'd3;
b_mant0 = 8'd199; b_mant1 = 8'd163; b_mant2 = 8'd142; b_mant3 = 8'd142;
a_exp0 = 10'd414; a_exp1 = 10'd375; a_exp2 = 10'd691; a_exp3 = 10'd547;
b_exp0 = 10'd87; b_exp1 = 10'd289; b_exp2 = 10'd255; b_exp3 = 10'd44;
a_sign0 = 4'd9; a_sign1 = 4'd11; a_sign2 = 4'd11; a_sign3 = 4'd14;
b_sign0 = 4'd5; b_sign1 = 4'd8; b_sign2 = 4'd16; b_sign3 = 4'd6;
@(posedge clk_i);
a_mant0 = 8'd15; a_mant1 = 8'd2; a_mant2 = 8'd94; a_mant3 = 8'd9;
b_mant0 = 8'd130; b_mant1 = 8'd23; b_mant2 = 8'd49; b_mant3 = 8'd169;
a_exp0 = 10'd763; a_exp1 = 10'd26; a_exp2 = 10'd300; a_exp3 = 10'd37;
b_exp0 = 10'd953; b_exp1 = 10'd229; b_exp2 = 10'd924; b_exp3 = 10'd215;
a_sign0 = 4'd7; a_sign1 = 4'd9; a_sign2 = 4'd5; a_sign3 = 4'd6;
b_sign0 = 4'd11; b_sign1 = 4'd12; b_sign2 = 4'd16; b_sign3 = 4'd2;
@(posedge clk_i);
a_mant0 = 8'd46; a_mant1 = 8'd91; a_mant2 = 8'd211; a_mant3 = 8'd112;
b_mant0 = 8'd143; b_mant1 = 8'd67; b_mant2 = 8'd94; b_mant3 = 8'd146;
a_exp0 = 10'd709; a_exp1 = 10'd110; a_exp2 = 10'd976; a_exp3 = 10'd442;
b_exp0 = 10'd240; b_exp1 = 10'd56; b_exp2 = 10'd612; b_exp3 = 10'd311;
a_sign0 = 4'd9; a_sign1 = 4'd0; a_sign2 = 4'd5; a_sign3 = 4'd0;
b_sign0 = 4'd10; b_sign1 = 4'd11; b_sign2 = 4'd0; b_sign3 = 4'd10;
@(posedge clk_i);
shared_exps0 = 8'd123;
shared_exps1 = 8'd142;
a_mant0 = 8'd169; a_mant1 = 8'd234; a_mant2 = 8'd148; a_mant3 = 8'd64;
b_mant0 = 8'd190; b_mant1 = 8'd17; b_mant2 = 8'd72; b_mant3 = 8'd51;
a_exp0 = 10'd828; a_exp1 = 10'd875; a_exp2 = 10'd372; a_exp3 = 10'd56;
b_exp0 = 10'd833; b_exp1 = 10'd277; b_exp2 = 10'd301; b_exp3 = 10'd558;
a_sign0 = 4'd4; a_sign1 = 4'd3; a_sign2 = 4'd4; a_sign3 = 4'd7;
b_sign0 = 4'd10; b_sign1 = 4'd13; b_sign2 = 4'd9; b_sign3 = 4'd14;
@(posedge clk_i);
a_mant0 = 8'd169; a_mant1 = 8'd50; a_mant2 = 8'd34; a_mant3 = 8'd75;
b_mant0 = 8'd53; b_mant1 = 8'd83; b_mant2 = 8'd213; b_mant3 = 8'd120;
a_exp0 = 10'd250; a_exp1 = 10'd380; a_exp2 = 10'd98; a_exp3 = 10'd976;
b_exp0 = 10'd445; b_exp1 = 10'd882; b_exp2 = 10'd712; b_exp3 = 10'd530;
a_sign0 = 4'd12; a_sign1 = 4'd15; a_sign2 = 4'd11; a_sign3 = 4'd15;
b_sign0 = 4'd13; b_sign1 = 4'd8; b_sign2 = 4'd11; b_sign3 = 4'd15;
@(posedge clk_i);
a_mant0 = 8'd168; a_mant1 = 8'd229; a_mant2 = 8'd230; a_mant3 = 8'd28;
b_mant0 = 8'd33; b_mant1 = 8'd4; b_mant2 = 8'd136; b_mant3 = 8'd179;
a_exp0 = 10'd919; a_exp1 = 10'd858; a_exp2 = 10'd679; a_exp3 = 10'd703;
b_exp0 = 10'd155; b_exp1 = 10'd46; b_exp2 = 10'd136; b_exp3 = 10'd824;
a_sign0 = 4'd13; a_sign1 = 4'd3; a_sign2 = 4'd10; a_sign3 = 4'd12;
b_sign0 = 4'd14; b_sign1 = 4'd7; b_sign2 = 4'd10; b_sign3 = 4'd4;
@(posedge clk_i);
a_mant0 = 8'd196; a_mant1 = 8'd11; a_mant2 = 8'd84; a_mant3 = 8'd124;
b_mant0 = 8'd165; b_mant1 = 8'd153; b_mant2 = 8'd141; b_mant3 = 8'd15;
a_exp0 = 10'd413; a_exp1 = 10'd20; a_exp2 = 10'd584; a_exp3 = 10'd498;
b_exp0 = 10'd499; b_exp1 = 10'd95; b_exp2 = 10'd15; b_exp3 = 10'd282;
a_sign0 = 4'd4; a_sign1 = 4'd8; a_sign2 = 4'd2; a_sign3 = 4'd0;
b_sign0 = 4'd5; b_sign1 = 4'd0; b_sign2 = 4'd1; b_sign3 = 4'd15;
@(posedge clk_i);
a_mant0 = 8'd93; a_mant1 = 8'd20; a_mant2 = 8'd115; a_mant3 = 8'd217;
b_mant0 = 8'd30; b_mant1 = 8'd193; b_mant2 = 8'd166; b_mant3 = 8'd143;
a_exp0 = 10'd491; a_exp1 = 10'd431; a_exp2 = 10'd440; a_exp3 = 10'd326;
b_exp0 = 10'd697; b_exp1 = 10'd824; b_exp2 = 10'd536; b_exp3 = 10'd171;
a_sign0 = 4'd8; a_sign1 = 4'd9; a_sign2 = 4'd15; a_sign3 = 4'd11;
b_sign0 = 4'd7; b_sign1 = 4'd9; b_sign2 = 4'd8; b_sign3 = 4'd4;
@(posedge clk_i);
a_mant0 = 8'd230; a_mant1 = 8'd69; a_mant2 = 8'd214; a_mant3 = 8'd89;
b_mant0 = 8'd149; b_mant1 = 8'd113; b_mant2 = 8'd98; b_mant3 = 8'd54;
a_exp0 = 10'd132; a_exp1 = 10'd869; a_exp2 = 10'd384; a_exp3 = 10'd10;
b_exp0 = 10'd487; b_exp1 = 10'd395; b_exp2 = 10'd892; b_exp3 = 10'd85;
a_sign0 = 4'd15; a_sign1 = 4'd1; a_sign2 = 4'd2; a_sign3 = 4'd2;
b_sign0 = 4'd4; b_sign1 = 4'd2; b_sign2 = 4'd8; b_sign3 = 4'd12;
@(posedge clk_i);
a_mant0 = 8'd255; a_mant1 = 8'd197; a_mant2 = 8'd74; a_mant3 = 8'd43;
b_mant0 = 8'd59; b_mant1 = 8'd142; b_mant2 = 8'd172; b_mant3 = 8'd196;
a_exp0 = 10'd598; a_exp1 = 10'd199; a_exp2 = 10'd871; a_exp3 = 10'd589;
b_exp0 = 10'd240; b_exp1 = 10'd18; b_exp2 = 10'd471; b_exp3 = 10'd759;
a_sign0 = 4'd16; a_sign1 = 4'd12; a_sign2 = 4'd8; a_sign3 = 4'd7;
b_sign0 = 4'd16; b_sign1 = 4'd4; b_sign2 = 4'd2; b_sign3 = 4'd11;
@(posedge clk_i);
a_mant0 = 8'd191; a_mant1 = 8'd41; a_mant2 = 8'd50; a_mant3 = 8'd253;
b_mant0 = 8'd235; b_mant1 = 8'd207; b_mant2 = 8'd205; b_mant3 = 8'd94;
a_exp0 = 10'd609; a_exp1 = 10'd241; a_exp2 = 10'd791; a_exp3 = 10'd237;
b_exp0 = 10'd511; b_exp1 = 10'd578; b_exp2 = 10'd244; b_exp3 = 10'd156;
a_sign0 = 4'd7; a_sign1 = 4'd15; a_sign2 = 4'd3; a_sign3 = 4'd6;
b_sign0 = 4'd3; b_sign1 = 4'd4; b_sign2 = 4'd13; b_sign3 = 4'd0;
@(posedge clk_i);
shared_exps0 = 8'd111;
shared_exps1 = 8'd75;
rstn = 0;
@(posedge clk_i);
rstn = 1;
a_mant0 = 8'd152; a_mant1 = 8'd6; a_mant2 = 8'd98; a_mant3 = 8'd162;
b_mant0 = 8'd153; b_mant1 = 8'd44; b_mant2 = 8'd85; b_mant3 = 8'd14;
a_exp0 = 10'd575; a_exp1 = 10'd906; a_exp2 = 10'd701; a_exp3 = 10'd940;
b_exp0 = 10'd485; b_exp1 = 10'd725; b_exp2 = 10'd130; b_exp3 = 10'd622;
a_sign0 = 4'd7; a_sign1 = 4'd9; a_sign2 = 4'd16; a_sign3 = 4'd14;
b_sign0 = 4'd2; b_sign1 = 4'd6; b_sign2 = 4'd1; b_sign3 = 4'd8;
@(posedge clk_i);
a_mant0 = 8'd150; a_mant1 = 8'd138; a_mant2 = 8'd3; a_mant3 = 8'd2;
b_mant0 = 8'd233; b_mant1 = 8'd197; b_mant2 = 8'd236; b_mant3 = 8'd45;
a_exp0 = 10'd312; a_exp1 = 10'd435; a_exp2 = 10'd685; a_exp3 = 10'd129;
b_exp0 = 10'd590; b_exp1 = 10'd382; b_exp2 = 10'd1015; b_exp3 = 10'd407;
a_sign0 = 4'd5; a_sign1 = 4'd13; a_sign2 = 4'd10; a_sign3 = 4'd5;
b_sign0 = 4'd4; b_sign1 = 4'd8; b_sign2 = 4'd14; b_sign3 = 4'd10;
@(posedge clk_i);
a_mant0 = 8'd50; a_mant1 = 8'd251; a_mant2 = 8'd242; a_mant3 = 8'd155;
b_mant0 = 8'd46; b_mant1 = 8'd102; b_mant2 = 8'd142; b_mant3 = 8'd83;
a_exp0 = 10'd892; a_exp1 = 10'd86; a_exp2 = 10'd250; a_exp3 = 10'd312;
b_exp0 = 10'd226; b_exp1 = 10'd768; b_exp2 = 10'd784; b_exp3 = 10'd428;
a_sign0 = 4'd14; a_sign1 = 4'd1; a_sign2 = 4'd0; a_sign3 = 4'd12;
b_sign0 = 4'd9; b_sign1 = 4'd10; b_sign2 = 4'd13; b_sign3 = 4'd4;
@(posedge clk_i);
a_mant0 = 8'd251; a_mant1 = 8'd121; a_mant2 = 8'd89; a_mant3 = 8'd25;
b_mant0 = 8'd173; b_mant1 = 8'd170; b_mant2 = 8'd107; b_mant3 = 8'd227;
a_exp0 = 10'd10; a_exp1 = 10'd902; a_exp2 = 10'd835; a_exp3 = 10'd627;
b_exp0 = 10'd525; b_exp1 = 10'd759; b_exp2 = 10'd891; b_exp3 = 10'd637;
a_sign0 = 4'd5; a_sign1 = 4'd12; a_sign2 = 4'd1; a_sign3 = 4'd1;
b_sign0 = 4'd5; b_sign1 = 4'd10; b_sign2 = 4'd15; b_sign3 = 4'd5;
@(posedge clk_i);
a_mant0 = 8'd106; a_mant1 = 8'd147; a_mant2 = 8'd67; a_mant3 = 8'd75;
b_mant0 = 8'd131; b_mant1 = 8'd37; b_mant2 = 8'd180; b_mant3 = 8'd77;
a_exp0 = 10'd400; a_exp1 = 10'd524; a_exp2 = 10'd67; a_exp3 = 10'd612;
b_exp0 = 10'd776; b_exp1 = 10'd72; b_exp2 = 10'd596; b_exp3 = 10'd792;
a_sign0 = 4'd0; a_sign1 = 4'd3; a_sign2 = 4'd13; a_sign3 = 4'd0;
b_sign0 = 4'd5; b_sign1 = 4'd11; b_sign2 = 4'd3; b_sign3 = 4'd15;
@(posedge clk_i);
a_mant0 = 8'd183; a_mant1 = 8'd120; a_mant2 = 8'd94; a_mant3 = 8'd192;
b_mant0 = 8'd17; b_mant1 = 8'd110; b_mant2 = 8'd110; b_mant3 = 8'd121;
a_exp0 = 10'd365; a_exp1 = 10'd867; a_exp2 = 10'd433; a_exp3 = 10'd120;
b_exp0 = 10'd766; b_exp1 = 10'd154; b_exp2 = 10'd1022; b_exp3 = 10'd1018;
a_sign0 = 4'd4; a_sign1 = 4'd5; a_sign2 = 4'd7; a_sign3 = 4'd9;
b_sign0 = 4'd1; b_sign1 = 4'd8; b_sign2 = 4'd3; b_sign3 = 4'd12;
@(posedge clk_i);
a_mant0 = 8'd181; a_mant1 = 8'd4; a_mant2 = 8'd235; a_mant3 = 8'd251;
b_mant0 = 8'd121; b_mant1 = 8'd169; b_mant2 = 8'd90; b_mant3 = 8'd91;
a_exp0 = 10'd285; a_exp1 = 10'd49; a_exp2 = 10'd702; a_exp3 = 10'd809;
b_exp0 = 10'd884; b_exp1 = 10'd108; b_exp2 = 10'd439; b_exp3 = 10'd180;
a_sign0 = 4'd0; a_sign1 = 4'd13; a_sign2 = 4'd10; a_sign3 = 4'd16;
b_sign0 = 4'd14; b_sign1 = 4'd16; b_sign2 = 4'd2; b_sign3 = 4'd0;
@(posedge clk_i);
shared_exps0 = 8'd134;
shared_exps1 = 8'd112;
a_mant0 = 8'd153; a_mant1 = 8'd68; a_mant2 = 8'd121; a_mant3 = 8'd65;
b_mant0 = 8'd169; b_mant1 = 8'd52; b_mant2 = 8'd52; b_mant3 = 8'd84;
a_exp0 = 10'd812; a_exp1 = 10'd227; a_exp2 = 10'd625; a_exp3 = 10'd156;
b_exp0 = 10'd641; b_exp1 = 10'd730; b_exp2 = 10'd896; b_exp3 = 10'd442;
a_sign0 = 4'd13; a_sign1 = 4'd15; a_sign2 = 4'd6; a_sign3 = 4'd13;
b_sign0 = 4'd8; b_sign1 = 4'd3; b_sign2 = 4'd0; b_sign3 = 4'd15;
@(posedge clk_i);
a_mant0 = 8'd228; a_mant1 = 8'd157; a_mant2 = 8'd122; a_mant3 = 8'd206;
b_mant0 = 8'd165; b_mant1 = 8'd252; b_mant2 = 8'd200; b_mant3 = 8'd36;
a_exp0 = 10'd211; a_exp1 = 10'd69; a_exp2 = 10'd135; a_exp3 = 10'd669;
b_exp0 = 10'd527; b_exp1 = 10'd243; b_exp2 = 10'd702; b_exp3 = 10'd880;
a_sign0 = 4'd8; a_sign1 = 4'd15; a_sign2 = 4'd11; a_sign3 = 4'd2;
b_sign0 = 4'd4; b_sign1 = 4'd11; b_sign2 = 4'd2; b_sign3 = 4'd12;
@(posedge clk_i);
a_mant0 = 8'd68; a_mant1 = 8'd135; a_mant2 = 8'd120; a_mant3 = 8'd63;
b_mant0 = 8'd200; b_mant1 = 8'd198; b_mant2 = 8'd4; b_mant3 = 8'd73;
a_exp0 = 10'd1017; a_exp1 = 10'd906; a_exp2 = 10'd996; a_exp3 = 10'd329;
b_exp0 = 10'd6; b_exp1 = 10'd657; b_exp2 = 10'd896; b_exp3 = 10'd869;
a_sign0 = 4'd8; a_sign1 = 4'd11; a_sign2 = 4'd3; a_sign3 = 4'd8;
b_sign0 = 4'd3; b_sign1 = 4'd8; b_sign2 = 4'd7; b_sign3 = 4'd5;
@(posedge clk_i);
a_mant0 = 8'd39; a_mant1 = 8'd190; a_mant2 = 8'd208; a_mant3 = 8'd115;
b_mant0 = 8'd1; b_mant1 = 8'd128; b_mant2 = 8'd84; b_mant3 = 8'd24;
a_exp0 = 10'd391; a_exp1 = 10'd825; a_exp2 = 10'd72; a_exp3 = 10'd37;
b_exp0 = 10'd958; b_exp1 = 10'd176; b_exp2 = 10'd796; b_exp3 = 10'd97;
a_sign0 = 4'd6; a_sign1 = 4'd0; a_sign2 = 4'd12; a_sign3 = 4'd2;
b_sign0 = 4'd6; b_sign1 = 4'd0; b_sign2 = 4'd6; b_sign3 = 4'd4;
@(posedge clk_i);
a_mant0 = 8'd7; a_mant1 = 8'd242; a_mant2 = 8'd88; a_mant3 = 8'd95;
b_mant0 = 8'd111; b_mant1 = 8'd157; b_mant2 = 8'd63; b_mant3 = 8'd24;
a_exp0 = 10'd734; a_exp1 = 10'd896; a_exp2 = 10'd818; a_exp3 = 10'd629;
b_exp0 = 10'd781; b_exp1 = 10'd375; b_exp2 = 10'd105; b_exp3 = 10'd426;
a_sign0 = 4'd4; a_sign1 = 4'd14; a_sign2 = 4'd15; a_sign3 = 4'd16;
b_sign0 = 4'd6; b_sign1 = 4'd16; b_sign2 = 4'd9; b_sign3 = 4'd11;
@(posedge clk_i);
a_mant0 = 8'd183; a_mant1 = 8'd94; a_mant2 = 8'd243; a_mant3 = 8'd5;
b_mant0 = 8'd29; b_mant1 = 8'd202; b_mant2 = 8'd71; b_mant3 = 8'd235;
a_exp0 = 10'd392; a_exp1 = 10'd792; a_exp2 = 10'd191; a_exp3 = 10'd236;
b_exp0 = 10'd166; b_exp1 = 10'd5; b_exp2 = 10'd783; b_exp3 = 10'd659;
a_sign0 = 4'd0; a_sign1 = 4'd16; a_sign2 = 4'd1; a_sign3 = 4'd0;
b_sign0 = 4'd1; b_sign1 = 4'd15; b_sign2 = 4'd4; b_sign3 = 4'd7;
@(posedge clk_i);
a_mant0 = 8'd56; a_mant1 = 8'd240; a_mant2 = 8'd143; a_mant3 = 8'd96;
b_mant0 = 8'd158; b_mant1 = 8'd2; b_mant2 = 8'd171; b_mant3 = 8'd22;
a_exp0 = 10'd261; a_exp1 = 10'd350; a_exp2 = 10'd599; a_exp3 = 10'd321;
b_exp0 = 10'd62; b_exp1 = 10'd206; b_exp2 = 10'd464; b_exp3 = 10'd992;
a_sign0 = 4'd2; a_sign1 = 4'd2; a_sign2 = 4'd15; a_sign3 = 4'd1;
b_sign0 = 4'd1; b_sign1 = 4'd11; b_sign2 = 4'd1; b_sign3 = 4'd16;
@(posedge clk_i);
a_mant0 = 8'd201; a_mant1 = 8'd133; a_mant2 = 8'd184; a_mant3 = 8'd99;
b_mant0 = 8'd197; b_mant1 = 8'd122; b_mant2 = 8'd170; b_mant3 = 8'd139;
a_exp0 = 10'd5; a_exp1 = 10'd180; a_exp2 = 10'd409; a_exp3 = 10'd681;
b_exp0 = 10'd27; b_exp1 = 10'd862; b_exp2 = 10'd991; b_exp3 = 10'd635;
a_sign0 = 4'd7; a_sign1 = 4'd4; a_sign2 = 4'd3; a_sign3 = 4'd5;
b_sign0 = 4'd7; b_sign1 = 4'd5; b_sign2 = 4'd1; b_sign3 = 4'd12;
@(posedge clk_i);
shared_exps0 = 8'd135;
shared_exps1 = 8'd120;
a_mant0 = 8'd136; a_mant1 = 8'd144; a_mant2 = 8'd251; a_mant3 = 8'd32;
b_mant0 = 8'd228; b_mant1 = 8'd47; b_mant2 = 8'd4; b_mant3 = 8'd179;
a_exp0 = 10'd221; a_exp1 = 10'd85; a_exp2 = 10'd906; a_exp3 = 10'd826;
b_exp0 = 10'd668; b_exp1 = 10'd118; b_exp2 = 10'd418; b_exp3 = 10'd821;
a_sign0 = 4'd6; a_sign1 = 4'd16; a_sign2 = 4'd4; a_sign3 = 4'd6;
b_sign0 = 4'd9; b_sign1 = 4'd4; b_sign2 = 4'd0; b_sign3 = 4'd13;
@(posedge clk_i);
a_mant0 = 8'd125; a_mant1 = 8'd198; a_mant2 = 8'd39; a_mant3 = 8'd219;
b_mant0 = 8'd148; b_mant1 = 8'd202; b_mant2 = 8'd9; b_mant3 = 8'd12;
a_exp0 = 10'd491; a_exp1 = 10'd424; a_exp2 = 10'd465; a_exp3 = 10'd980;
b_exp0 = 10'd283; b_exp1 = 10'd331; b_exp2 = 10'd85; b_exp3 = 10'd371;
a_sign0 = 4'd13; a_sign1 = 4'd15; a_sign2 = 4'd11; a_sign3 = 4'd4;
b_sign0 = 4'd5; b_sign1 = 4'd9; b_sign2 = 4'd0; b_sign3 = 4'd1;
@(posedge clk_i);
a_mant0 = 8'd183; a_mant1 = 8'd5; a_mant2 = 8'd253; a_mant3 = 8'd178;
b_mant0 = 8'd142; b_mant1 = 8'd89; b_mant2 = 8'd152; b_mant3 = 8'd182;
a_exp0 = 10'd430; a_exp1 = 10'd84; a_exp2 = 10'd73; a_exp3 = 10'd135;
b_exp0 = 10'd481; b_exp1 = 10'd646; b_exp2 = 10'd640; b_exp3 = 10'd32;
a_sign0 = 4'd16; a_sign1 = 4'd4; a_sign2 = 4'd16; a_sign3 = 4'd16;
b_sign0 = 4'd8; b_sign1 = 4'd9; b_sign2 = 4'd5; b_sign3 = 4'd3;
@(posedge clk_i);
a_mant0 = 8'd253; a_mant1 = 8'd54; a_mant2 = 8'd80; a_mant3 = 8'd112;
b_mant0 = 8'd72; b_mant1 = 8'd156; b_mant2 = 8'd169; b_mant3 = 8'd69;
a_exp0 = 10'd1001; a_exp1 = 10'd277; a_exp2 = 10'd858; a_exp3 = 10'd656;
b_exp0 = 10'd288; b_exp1 = 10'd100; b_exp2 = 10'd299; b_exp3 = 10'd44;
a_sign0 = 4'd2; a_sign1 = 4'd6; a_sign2 = 4'd3; a_sign3 = 4'd13;
b_sign0 = 4'd7; b_sign1 = 4'd0; b_sign2 = 4'd11; b_sign3 = 4'd1;
@(posedge clk_i);
a_mant0 = 8'd122; a_mant1 = 8'd189; a_mant2 = 8'd130; a_mant3 = 8'd234;
b_mant0 = 8'd47; b_mant1 = 8'd255; b_mant2 = 8'd86; b_mant3 = 8'd217;
a_exp0 = 10'd501; a_exp1 = 10'd720; a_exp2 = 10'd503; a_exp3 = 10'd182;
b_exp0 = 10'd696; b_exp1 = 10'd364; b_exp2 = 10'd688; b_exp3 = 10'd271;
a_sign0 = 4'd8; a_sign1 = 4'd11; a_sign2 = 4'd14; a_sign3 = 4'd2;
b_sign0 = 4'd5; b_sign1 = 4'd5; b_sign2 = 4'd5; b_sign3 = 4'd4;
@(posedge clk_i);
a_mant0 = 8'd88; a_mant1 = 8'd206; a_mant2 = 8'd77; a_mant3 = 8'd18;
b_mant0 = 8'd23; b_mant1 = 8'd231; b_mant2 = 8'd213; b_mant3 = 8'd108;
a_exp0 = 10'd877; a_exp1 = 10'd593; a_exp2 = 10'd484; a_exp3 = 10'd216;
b_exp0 = 10'd248; b_exp1 = 10'd169; b_exp2 = 10'd960; b_exp3 = 10'd814;
a_sign0 = 4'd2; a_sign1 = 4'd11; a_sign2 = 4'd10; a_sign3 = 4'd11;
b_sign0 = 4'd12; b_sign1 = 4'd1; b_sign2 = 4'd11; b_sign3 = 4'd16;
@(posedge clk_i);
a_mant0 = 8'd89; a_mant1 = 8'd244; a_mant2 = 8'd163; a_mant3 = 8'd184;
b_mant0 = 8'd21; b_mant1 = 8'd174; b_mant2 = 8'd107; b_mant3 = 8'd63;
a_exp0 = 10'd293; a_exp1 = 10'd903; a_exp2 = 10'd344; a_exp3 = 10'd452;
b_exp0 = 10'd252; b_exp1 = 10'd933; b_exp2 = 10'd747; b_exp3 = 10'd411;
a_sign0 = 4'd9; a_sign1 = 4'd3; a_sign2 = 4'd12; a_sign3 = 4'd12;
b_sign0 = 4'd5; b_sign1 = 4'd4; b_sign2 = 4'd7; b_sign3 = 4'd6;
@(posedge clk_i);
a_mant0 = 8'd21; a_mant1 = 8'd21; a_mant2 = 8'd60; a_mant3 = 8'd184;
b_mant0 = 8'd116; b_mant1 = 8'd108; b_mant2 = 8'd194; b_mant3 = 8'd115;
a_exp0 = 10'd811; a_exp1 = 10'd772; a_exp2 = 10'd867; a_exp3 = 10'd739;
b_exp0 = 10'd934; b_exp1 = 10'd873; b_exp2 = 10'd467; b_exp3 = 10'd838;
a_sign0 = 4'd15; a_sign1 = 4'd1; a_sign2 = 4'd10; a_sign3 = 4'd8;
b_sign0 = 4'd16; b_sign1 = 4'd15; b_sign2 = 4'd16; b_sign3 = 4'd0;
@(posedge clk_i);
shared_exps0 = 8'd140;
shared_exps1 = 8'd119;
a_mant0 = 8'd222; a_mant1 = 8'd33; a_mant2 = 8'd101; a_mant3 = 8'd69;
b_mant0 = 8'd88; b_mant1 = 8'd33; b_mant2 = 8'd224; b_mant3 = 8'd197;
a_exp0 = 10'd22; a_exp1 = 10'd473; a_exp2 = 10'd936; a_exp3 = 10'd456;
b_exp0 = 10'd829; b_exp1 = 10'd935; b_exp2 = 10'd603; b_exp3 = 10'd884;
a_sign0 = 4'd12; a_sign1 = 4'd6; a_sign2 = 4'd8; a_sign3 = 4'd12;
b_sign0 = 4'd3; b_sign1 = 4'd6; b_sign2 = 4'd13; b_sign3 = 4'd0;
@(posedge clk_i);
a_mant0 = 8'd116; a_mant1 = 8'd214; a_mant2 = 8'd143; a_mant3 = 8'd206;
b_mant0 = 8'd139; b_mant1 = 8'd235; b_mant2 = 8'd37; b_mant3 = 8'd203;
a_exp0 = 10'd705; a_exp1 = 10'd376; a_exp2 = 10'd754; a_exp3 = 10'd798;
b_exp0 = 10'd370; b_exp1 = 10'd249; b_exp2 = 10'd713; b_exp3 = 10'd814;
a_sign0 = 4'd11; a_sign1 = 4'd13; a_sign2 = 4'd16; a_sign3 = 4'd10;
b_sign0 = 4'd16; b_sign1 = 4'd4; b_sign2 = 4'd2; b_sign3 = 4'd8;
@(posedge clk_i);
a_mant0 = 8'd132; a_mant1 = 8'd142; a_mant2 = 8'd136; a_mant3 = 8'd238;
b_mant0 = 8'd47; b_mant1 = 8'd30; b_mant2 = 8'd226; b_mant3 = 8'd172;
a_exp0 = 10'd40; a_exp1 = 10'd359; a_exp2 = 10'd768; a_exp3 = 10'd156;
b_exp0 = 10'd84; b_exp1 = 10'd667; b_exp2 = 10'd693; b_exp3 = 10'd938;
a_sign0 = 4'd14; a_sign1 = 4'd2; a_sign2 = 4'd3; a_sign3 = 4'd14;
b_sign0 = 4'd1; b_sign1 = 4'd6; b_sign2 = 4'd10; b_sign3 = 4'd15;
@(posedge clk_i);
a_mant0 = 8'd87; a_mant1 = 8'd131; a_mant2 = 8'd52; a_mant3 = 8'd82;
b_mant0 = 8'd156; b_mant1 = 8'd32; b_mant2 = 8'd77; b_mant3 = 8'd255;
a_exp0 = 10'd528; a_exp1 = 10'd725; a_exp2 = 10'd729; a_exp3 = 10'd432;
b_exp0 = 10'd749; b_exp1 = 10'd566; b_exp2 = 10'd415; b_exp3 = 10'd46;
a_sign0 = 4'd4; a_sign1 = 4'd15; a_sign2 = 4'd12; a_sign3 = 4'd9;
b_sign0 = 4'd2; b_sign1 = 4'd1; b_sign2 = 4'd1; b_sign3 = 4'd16;
@(posedge clk_i);
a_mant0 = 8'd234; a_mant1 = 8'd196; a_mant2 = 8'd98; a_mant3 = 8'd143;
b_mant0 = 8'd76; b_mant1 = 8'd94; b_mant2 = 8'd129; b_mant3 = 8'd191;
a_exp0 = 10'd485; a_exp1 = 10'd107; a_exp2 = 10'd613; a_exp3 = 10'd12;
b_exp0 = 10'd902; b_exp1 = 10'd250; b_exp2 = 10'd439; b_exp3 = 10'd258;
a_sign0 = 4'd10; a_sign1 = 4'd8; a_sign2 = 4'd0; a_sign3 = 4'd12;
b_sign0 = 4'd11; b_sign1 = 4'd3; b_sign2 = 4'd10; b_sign3 = 4'd6;
@(posedge clk_i);
a_mant0 = 8'd14; a_mant1 = 8'd111; a_mant2 = 8'd82; a_mant3 = 8'd144;
b_mant0 = 8'd84; b_mant1 = 8'd179; b_mant2 = 8'd55; b_mant3 = 8'd66;
a_exp0 = 10'd241; a_exp1 = 10'd704; a_exp2 = 10'd803; a_exp3 = 10'd837;
b_exp0 = 10'd82; b_exp1 = 10'd6; b_exp2 = 10'd258; b_exp3 = 10'd402;
a_sign0 = 4'd1; a_sign1 = 4'd16; a_sign2 = 4'd1; a_sign3 = 4'd6;
b_sign0 = 4'd12; b_sign1 = 4'd4; b_sign2 = 4'd14; b_sign3 = 4'd11;
@(posedge clk_i);
a_mant0 = 8'd61; a_mant1 = 8'd224; a_mant2 = 8'd71; a_mant3 = 8'd196;
b_mant0 = 8'd139; b_mant1 = 8'd136; b_mant2 = 8'd107; b_mant3 = 8'd4;
a_exp0 = 10'd18; a_exp1 = 10'd980; a_exp2 = 10'd987; a_exp3 = 10'd940;
b_exp0 = 10'd324; b_exp1 = 10'd236; b_exp2 = 10'd853; b_exp3 = 10'd517;
a_sign0 = 4'd4; a_sign1 = 4'd12; a_sign2 = 4'd0; a_sign3 = 4'd12;
b_sign0 = 4'd6; b_sign1 = 4'd7; b_sign2 = 4'd6; b_sign3 = 4'd6;
@(posedge clk_i);
a_mant0 = 8'd91; a_mant1 = 8'd34; a_mant2 = 8'd96; a_mant3 = 8'd142;
b_mant0 = 8'd160; b_mant1 = 8'd244; b_mant2 = 8'd11; b_mant3 = 8'd37;
a_exp0 = 10'd91; a_exp1 = 10'd209; a_exp2 = 10'd581; a_exp3 = 10'd69;
b_exp0 = 10'd379; b_exp1 = 10'd226; b_exp2 = 10'd7; b_exp3 = 10'd797;
a_sign0 = 4'd9; a_sign1 = 4'd0; a_sign2 = 4'd8; a_sign3 = 4'd12;
b_sign0 = 4'd4; b_sign1 = 4'd7; b_sign2 = 4'd11; b_sign3 = 4'd11;
@(posedge clk_i);
shared_exps0 = 8'd136;
shared_exps1 = 8'd105;
rstn = 0;
@(posedge clk_i);
rstn = 1;
a_mant0 = 8'd229; a_mant1 = 8'd83; a_mant2 = 8'd245; a_mant3 = 8'd236;
b_mant0 = 8'd152; b_mant1 = 8'd163; b_mant2 = 8'd200; b_mant3 = 8'd122;
a_exp0 = 10'd777; a_exp1 = 10'd354; a_exp2 = 10'd30; a_exp3 = 10'd646;
b_exp0 = 10'd770; b_exp1 = 10'd779; b_exp2 = 10'd476; b_exp3 = 10'd525;
a_sign0 = 4'd6; a_sign1 = 4'd0; a_sign2 = 4'd6; a_sign3 = 4'd12;
b_sign0 = 4'd9; b_sign1 = 4'd15; b_sign2 = 4'd4; b_sign3 = 4'd15;
@(posedge clk_i);
a_mant0 = 8'd27; a_mant1 = 8'd118; a_mant2 = 8'd8; a_mant3 = 8'd122;
b_mant0 = 8'd157; b_mant1 = 8'd190; b_mant2 = 8'd126; b_mant3 = 8'd182;
a_exp0 = 10'd822; a_exp1 = 10'd204; a_exp2 = 10'd85; a_exp3 = 10'd470;
b_exp0 = 10'd123; b_exp1 = 10'd637; b_exp2 = 10'd354; b_exp3 = 10'd64;
a_sign0 = 4'd16; a_sign1 = 4'd8; a_sign2 = 4'd14; a_sign3 = 4'd15;
b_sign0 = 4'd1; b_sign1 = 4'd7; b_sign2 = 4'd2; b_sign3 = 4'd7;
@(posedge clk_i);
a_mant0 = 8'd34; a_mant1 = 8'd252; a_mant2 = 8'd82; a_mant3 = 8'd22;
b_mant0 = 8'd132; b_mant1 = 8'd205; b_mant2 = 8'd19; b_mant3 = 8'd213;
a_exp0 = 10'd346; a_exp1 = 10'd798; a_exp2 = 10'd244; a_exp3 = 10'd564;
b_exp0 = 10'd10; b_exp1 = 10'd21; b_exp2 = 10'd170; b_exp3 = 10'd915;
a_sign0 = 4'd12; a_sign1 = 4'd14; a_sign2 = 4'd14; a_sign3 = 4'd5;
b_sign0 = 4'd12; b_sign1 = 4'd7; b_sign2 = 4'd11; b_sign3 = 4'd10;
$dumpoff;
$finish;
end
endmodule
